/* Verilog module written by vlogFanout (qflow) */
/* With clock tree generation and fanout reduction */
/* and gate resizing */

module RISCV32I(
    input CLK,
    output [31:0] DMEM_ADDR,
    input [31:0] DMEM_DATA_L,
    output [31:0] DMEM_DATA_S,
    output DMEM_WEN,
    output [31:0] IMEM_ADDR,
    input [31:0] IMEM_DATA,
    input IRQ
);

wire _4972_ ;
wire _4552_ ;
wire _4132_ ;
wire _5757_ ;
wire _5337_ ;
wire _9170_ ;
wire _1677_ ;
wire _1257_ ;
wire _7903_ ;
wire _5090_ ;
wire _588_ ;
wire _168_ ;
wire _3823_ ;
wire _3403_ ;
wire _6295_ ;
wire _4608_ ;
wire _8861_ ;
wire _8441_ ;
wire _8021_ ;
wire \datapath.alu.b_4_bF$buf1  ;
wire _4781_ ;
wire _4361_ ;
wire _800_ ;
wire _5986_ ;
wire _5566_ ;
wire _5146_ ;
wire _60_ ;
wire _2783__bF$buf0 ;
wire _2783__bF$buf1 ;
wire _1486_ ;
wire _2783__bF$buf2 ;
wire _1066_ ;
wire _2783__bF$buf3 ;
wire _2783__bF$buf4 ;
wire _5586__bF$buf0 ;
wire _5586__bF$buf1 ;
wire _7712_ ;
wire _5586__bF$buf2 ;
wire _5586__bF$buf3 ;
wire _5586__bF$buf4 ;
wire _397_ ;
wire _4899__bF$buf0 ;
wire _4899__bF$buf1 ;
wire _4899__bF$buf2 ;
wire _4899__bF$buf3 ;
wire _4899__bF$buf4 ;
wire _8917_ ;
wire _4899__bF$buf5 ;
wire _4899__bF$buf6 ;
wire _4899__bF$buf7 ;
wire _4899__bF$buf8 ;
wire _4899__bF$buf9 ;
wire _3632_ ;
wire _3212_ ;
wire _4837_ ;
wire _4417_ ;
wire _8670_ ;
wire _8250_ ;
wire \datapath.immediatedecoder._06_  ;
wire _9035_ ;
wire _4590_ ;
wire _4170_ ;
wire _2903_ ;
wire _5795_ ;
wire _5375_ ;
wire _1295_ ;
wire _7941_ ;
wire _7521_ ;
wire _7101_ ;
wire _8726_ ;
wire _8306_ ;
wire _3861_ ;
wire _3441_ ;
wire _3021_ ;
wire _4646_ ;
wire _4226_ ;
wire CLK_bF$buf50 ;
wire CLK_bF$buf51 ;
wire CLK_bF$buf52 ;
wire CLK_bF$buf53 ;
wire CLK_bF$buf54 ;
wire CLK_bF$buf55 ;
wire CLK_bF$buf56 ;
wire CLK_bF$buf57 ;
wire CLK_bF$buf58 ;
wire CLK_bF$buf59 ;
wire _2712_ ;
wire _5184_ ;
wire _3917_ ;
wire _6389_ ;
wire _7750_ ;
wire _7330_ ;
wire _8955_ ;
wire _8535_ ;
wire _8115_ ;
wire _3670_ ;
wire _3250_ ;
wire _4875_ ;
wire _4455_ ;
wire _4035_ ;
wire [31:0] \datapath.memoryinterface.byte_size_store.storebyte  ;
wire _6601_ ;
wire _9073_ ;
wire _7806_ ;
wire _2941_ ;
wire _2521_ ;
wire _2101_ ;
wire _3726_ ;
wire _3306_ ;
wire _6198_ ;
wire _8764_ ;
wire _8344_ ;
wire _9129_ ;
wire _4684_ ;
wire _4264_ ;
wire _703_ ;
wire _5889_ ;
wire _5469_ ;
wire _5049_ ;
wire _6830_ ;
wire _6410_ ;
wire _1389_ ;
wire _7615_ ;
wire _2750_ ;
wire _2330_ ;
wire _3955_ ;
wire _3535_ ;
wire _3115_ ;
wire _8993_ ;
wire _8573_ ;
wire _8153_ ;
wire _19_ ;
wire _1601_ ;
wire _4493_ ;
wire _4073_ ;
wire \datapath.idinstr_20_bF$buf12  ;
wire _932_ ;
wire _512_ ;
wire _2806_ ;
wire _5698_ ;
wire _5278_ ;
wire [1:0] asel ;
wire _7418__bF$buf0 ;
wire _7418__bF$buf1 ;
wire _7418__bF$buf2 ;
wire _7418__bF$buf3 ;
wire _7418__bF$buf4 ;
wire _1198_ ;
wire _7844_ ;
wire _7424_ ;
wire _7004_ ;
wire [31:0] \datapath.registers.838[15]  ;
wire _8629_ ;
wire _8209_ ;
wire _3764_ ;
wire _3344_ ;
wire _4969_ ;
wire _4549_ ;
wire \datapath.idinstr_21_bF$buf21  ;
wire _4129_ ;
wire _5910_ ;
wire _8382_ ;
wire _1830_ ;
wire _1410_ ;
wire _9167_ ;
wire _741_ ;
wire _321_ ;
wire _2615_ ;
wire _5087_ ;
wire _7422__bF$buf0 ;
wire _7422__bF$buf1 ;
wire \datapath.idinstr_15_bF$buf26  ;
wire _7422__bF$buf2 ;
wire _7422__bF$buf3 ;
wire _7422__bF$buf4 ;
wire \datapath.idinstr_22_bF$buf30  ;
wire _7653_ ;
wire _7233_ ;
wire _8858_ ;
wire _8438_ ;
wire _8018_ ;
wire _3993_ ;
wire _3573_ ;
wire _3153_ ;
wire _4778_ ;
wire _4358_ ;
wire _8191_ ;
wire _5653__bF$buf0 ;
wire _5653__bF$buf1 ;
wire _5653__bF$buf2 ;
wire _5653__bF$buf3 ;
wire _5653__bF$buf4 ;
wire _5653__bF$buf5 ;
wire _5653__bF$buf6 ;
wire _5653__bF$buf7 ;
wire \datapath.idinstr_16_bF$buf35  ;
wire _57_ ;
wire _6924_ ;
wire _6504_ ;
wire \datapath.idinstr_20_bF$buf50  ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _7709_ ;
wire _2844_ ;
wire _2424_ ;
wire _2004_ ;
wire _3629_ ;
wire _3209_ ;
wire _7882_ ;
wire _7462_ ;
wire _7042_ ;
wire _8667_ ;
wire _8247_ ;
wire _3382_ ;
wire _4587_ ;
wire _4167_ ;
wire _606_ ;
wire _6733_ ;
wire _6313_ ;
wire _7938_ ;
wire _7518_ ;
wire _2653_ ;
wire _2233_ ;
wire _3858_ ;
wire _3438_ ;
wire _3018_ ;
wire _7691_ ;
wire _7271_ ;
wire _8896_ ;
wire _8476_ ;
wire _8056_ ;
wire _3191_ ;
wire _1924_ ;
wire _1504_ ;
wire _4396_ ;
wire _835_ ;
wire _415_ ;
wire _2709_ ;
wire _95_ ;
wire _6962_ ;
wire _6542_ ;
wire _6122_ ;
wire _7747_ ;
wire _7327_ ;
wire _2882_ ;
wire _2462_ ;
wire _2042_ ;
wire _3667_ ;
wire _3247_ ;
wire _7080_ ;
wire _5813_ ;
wire _8285_ ;
wire _1733_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _2938_ ;
wire _2518_ ;
wire _4847__bF$buf0 ;
wire _4847__bF$buf1 ;
wire _4847__bF$buf2 ;
wire _4847__bF$buf3 ;
wire _4847__bF$buf4 ;
wire _6771_ ;
wire _6351_ ;
wire _7976_ ;
wire _7556_ ;
wire _7136_ ;
wire _2691_ ;
wire _2271_ ;
wire _3896_ ;
wire _3476_ ;
wire _3056_ ;
wire _5622_ ;
wire _5202_ ;
wire _8094_ ;
wire _6827_ ;
wire _6407_ ;
wire _1962_ ;
wire _1542_ ;
wire _1122_ ;
wire _873_ ;
wire _453_ ;
wire _4851__bF$buf0 ;
wire _4851__bF$buf1 ;
wire _2747_ ;
wire _4851__bF$buf2 ;
wire _2327_ ;
wire _4851__bF$buf3 ;
wire _4851__bF$buf4 ;
wire _6580_ ;
wire _6160_ ;
wire _7785_ ;
wire _7365_ ;
wire _2080_ ;
wire _3285_ ;
wire _5851_ ;
wire _5431_ ;
wire _5011_ ;
wire _929_ ;
wire _509_ ;
wire _6636_ ;
wire _6216_ ;
wire _1771_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _2976_ ;
wire _2556_ ;
wire _2136_ ;
wire _4702_ ;
wire _7594_ ;
wire _7174_ ;
wire _2767__bF$buf0 ;
wire _2767__bF$buf1 ;
wire _2767__bF$buf2 ;
wire _2767__bF$buf3 ;
wire _2767__bF$buf4 ;
wire \datapath.idinstr_21_bF$buf18  ;
wire _5907_ ;
wire _8799_ ;
wire _8379_ ;
wire _3094_ ;
wire _1827_ ;
wire _1407_ ;
wire _4299_ ;
wire _5660_ ;
wire _5240_ ;
wire _738_ ;
wire _318_ ;
wire \datapath.idinstr_17_bF$buf3  ;
wire _6865_ ;
wire _6445_ ;
wire _6025_ ;
wire _1580_ ;
wire _1160_ ;
wire _491_ ;
wire \datapath.idinstr_22_bF$buf27  ;
wire _2785_ ;
wire _2365_ ;
wire _4931_ ;
wire _4511_ ;
wire _5716_ ;
wire _8188_ ;
wire _1636_ ;
wire _1216_ ;
wire \datapath.idinstr_21_bF$buf3  ;
wire \datapath.idinstr_20_bF$buf47  ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _6674_ ;
wire _6254_ ;
wire _7879_ ;
wire _7459_ ;
wire _7039_ ;
wire _2594_ ;
wire _2174_ ;
wire _8820_ ;
wire _8400_ ;
wire _3799_ ;
wire _3379_ ;
wire _286__bF$buf0 ;
wire _286__bF$buf1 ;
wire _286__bF$buf2 ;
wire _286__bF$buf3 ;
wire _286__bF$buf4 ;
wire _4740_ ;
wire _4320_ ;
wire _5945_ ;
wire _5525_ ;
wire _5105_ ;
wire _1865_ ;
wire _1445_ ;
wire _1025_ ;
wire _776_ ;
wire _356_ ;
wire _6483_ ;
wire _6063_ ;
wire _7688_ ;
wire _7268_ ;
wire _3188_ ;
wire _5754_ ;
wire _5334_ ;
wire _6959_ ;
wire _6539_ ;
wire _6119_ ;
wire _1674_ ;
wire _1254_ ;
wire _7900_ ;
wire _585_ ;
wire _165_ ;
wire _2879_ ;
wire _2459_ ;
wire _2039_ ;
wire _3820_ ;
wire _3400_ ;
wire _6292_ ;
wire _4605_ ;
wire _7497_ ;
wire _7077_ ;
wire _5983_ ;
wire _5563_ ;
wire _5143_ ;
wire _6768_ ;
wire _6348_ ;
wire _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _2688_ ;
wire _2268_ ;
wire _8914_ ;
wire _4834_ ;
wire _4414_ ;
wire _5619_ ;
wire _9032_ ;
wire \datapath.alu.b_2_bF$buf5  ;
wire _1959_ ;
wire _1539_ ;
wire _1119_ ;
wire _2900_ ;
wire _5792_ ;
wire _5372_ ;
wire _6997_ ;
wire _6577_ ;
wire _6157_ ;
wire _1292_ ;
wire _2497_ ;
wire _2077_ ;
wire _8723_ ;
wire _8303_ ;
wire _4643_ ;
wire _4223_ ;
wire CLK_bF$buf20 ;
wire CLK_bF$buf21 ;
wire CLK_bF$buf22 ;
wire CLK_bF$buf23 ;
wire CLK_bF$buf24 ;
wire CLK_bF$buf25 ;
wire CLK_bF$buf26 ;
wire CLK_bF$buf27 ;
wire CLK_bF$buf28 ;
wire CLK_bF$buf29 ;
wire _5848_ ;
wire _5428_ ;
wire _5008_ ;
wire _1768_ ;
wire _1348_ ;
wire _5181_ ;
wire _679_ ;
wire _259_ ;
wire [31:0] \datapath.registers.838[30]  ;
wire _3914_ ;
wire _6386_ ;
wire _8952_ ;
wire _8532_ ;
wire _8112_ ;
wire _4872_ ;
wire _4452_ ;
wire _4032_ ;
wire _5657_ ;
wire _5237_ ;
wire _9070_ ;
wire _1997_ ;
wire _1577_ ;
wire [31:0] \datapath.registers.838[6]  ;
wire _1157_ ;
wire _7803_ ;
wire _488_ ;
wire _3723_ ;
wire _3303_ ;
wire _6195_ ;
wire _4928_ ;
wire _4508_ ;
wire _8761_ ;
wire _8341_ ;
wire _9126_ ;
wire _4681_ ;
wire _4261_ ;
wire _700_ ;
wire _5886_ ;
wire _5466_ ;
wire _5046_ ;
wire _1386_ ;
wire _7612_ ;
wire _297_ ;
wire \datapath.idinstr_20_hier0_bF$buf4  ;
wire _8817_ ;
wire _3952_ ;
wire _3532_ ;
wire _3112_ ;
wire _4737_ ;
wire _4317_ ;
wire _0__1_bF$buf10 ;
wire _8990_ ;
wire _8570_ ;
wire _8150_ ;
wire _16_ ;
wire _4490_ ;
wire _4070_ ;
wire _2803_ ;
wire _5695_ ;
wire _5275_ ;
wire _1195_ ;
wire _7841_ ;
wire _7421_ ;
wire _7001_ ;
wire [31:0] \datapath.regcwb  ;
wire _8626_ ;
wire _8206_ ;
wire _3761_ ;
wire _3341_ ;
wire _4966_ ;
wire _4546_ ;
wire _4126_ ;
wire _9164_ ;
wire _2612_ ;
wire _5084_ ;
wire \datapath.idinstr_15_bF$buf23  ;
wire _3817_ ;
wire _6289_ ;
wire _7650_ ;
wire _7230_ ;
wire _8855_ ;
wire _8435_ ;
wire _8015_ ;
wire _3990_ ;
wire _3570_ ;
wire _3150_ ;
wire _4835__bF$buf0 ;
wire _4835__bF$buf1 ;
wire _4835__bF$buf2 ;
wire _4835__bF$buf3 ;
wire _4835__bF$buf4 ;
wire _4775_ ;
wire _4355_ ;
wire [31:0] \datapath.csr.mvect  ;
wire \datapath.idinstr_16_bF$buf32  ;
wire _54_ ;
wire _6921_ ;
wire _6501_ ;
wire _7706_ ;
wire _2841_ ;
wire _2421_ ;
wire _2001_ ;
wire _3626_ ;
wire _3206_ ;
wire _6098_ ;
wire _8664_ ;
wire _8244_ ;
wire _9029_ ;
wire _4584_ ;
wire _4164_ ;
wire _603_ ;
wire _5789_ ;
wire _5369_ ;
wire _6730_ ;
wire _6310_ ;
wire _1289_ ;
wire _7935_ ;
wire _7515_ ;
wire _2650_ ;
wire _2230_ ;
wire _3855_ ;
wire _3435_ ;
wire _3015_ ;
wire _8893_ ;
wire _8473_ ;
wire _8053_ ;
wire _1921_ ;
wire _1501_ ;
wire _4393_ ;
wire _832_ ;
wire _412_ ;
wire _2706_ ;
wire _5598_ ;
wire _5178_ ;
wire _92_ ;
wire _1098_ ;
wire _7744_ ;
wire _7324_ ;
wire _8949_ ;
wire _8529_ ;
wire _8109_ ;
wire _3664_ ;
wire _3244_ ;
wire _7425__bF$buf0 ;
wire _7425__bF$buf1 ;
wire _7425__bF$buf2 ;
wire _7425__bF$buf3 ;
wire _7425__bF$buf4 ;
wire _7425__bF$buf5 ;
wire _7425__bF$buf6 ;
wire _7425__bF$buf7 ;
wire _7425__bF$buf8 ;
wire _7425__bF$buf9 ;
wire _4869_ ;
wire _4449_ ;
wire _4029_ ;
wire _5810_ ;
wire _8282_ ;
wire _1730_ ;
wire _1310_ ;
wire _9067_ ;
wire _641_ ;
wire _221_ ;
wire _2935_ ;
wire _2515_ ;
wire _7973_ ;
wire _7553_ ;
wire _7133_ ;
wire _8758_ ;
wire _8338_ ;
wire _3893_ ;
wire _3473_ ;
wire _3053_ ;
wire _4678_ ;
wire _4258_ ;
wire _8091_ ;
wire _6824_ ;
wire _6404_ ;
wire _870_ ;
wire _450_ ;
wire _7609_ ;
wire _2744_ ;
wire _2324_ ;
wire _3949_ ;
wire _3529_ ;
wire _3109_ ;
wire _7782_ ;
wire _7362_ ;
wire _8987_ ;
wire _8567_ ;
wire _8147_ ;
wire _3282_ ;
wire _4487_ ;
wire _4067_ ;
wire _926_ ;
wire _506_ ;
wire _6633_ ;
wire _6213_ ;
wire _7838_ ;
wire _7418_ ;
wire _2973_ ;
wire _2553_ ;
wire _2133_ ;
wire _3758_ ;
wire _3338_ ;
wire _7591_ ;
wire _7171_ ;
wire \datapath.idinstr_21_bF$buf15  ;
wire _5904_ ;
wire _8796_ ;
wire _8376_ ;
wire _3091_ ;
wire _1824_ ;
wire _1404_ ;
wire _4296_ ;
wire _735_ ;
wire _315_ ;
wire \datapath.idinstr_17_bF$buf0  ;
wire _2609_ ;
wire _6862_ ;
wire _6442_ ;
wire _6022_ ;
wire \datapath.idinstr_22_bF$buf24  ;
wire _7647_ ;
wire _7227_ ;
wire _2782_ ;
wire _2362_ ;
wire _3987_ ;
wire _3567_ ;
wire _3147_ ;
wire _5713_ ;
wire _8185_ ;
wire \datapath.idinstr_16_bF$buf29  ;
wire _6918_ ;
wire _1633_ ;
wire _1213_ ;
wire \datapath.idinstr_21_bF$buf0  ;
wire \datapath.idinstr_20_bF$buf44  ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire _2838_ ;
wire \datapath.idinstr_15_bF$buf7  ;
wire _2418_ ;
wire _6671_ ;
wire _6251_ ;
wire \controlunit.mret  ;
wire _7876_ ;
wire _7456_ ;
wire _7036_ ;
wire _2591_ ;
wire _2171_ ;
wire IRQ ;
wire _3796_ ;
wire _3376_ ;
wire _5942_ ;
wire _5522_ ;
wire _5102_ ;
wire _6727_ ;
wire _6307_ ;
wire _1862_ ;
wire _1442_ ;
wire _1022_ ;
wire _773_ ;
wire _353_ ;
wire _2647_ ;
wire _2227_ ;
wire _6480_ ;
wire _6060_ ;
wire _7685_ ;
wire _7265_ ;
wire _3185_ ;
wire _1918_ ;
wire _5751_ ;
wire _5331_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _6956_ ;
wire _6536_ ;
wire _6116_ ;
wire _1671_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _2876_ ;
wire _2456_ ;
wire _2036_ ;
wire _4602_ ;
wire _7494_ ;
wire _7074_ ;
wire _5807_ ;
wire _8699_ ;
wire _8279_ ;
wire _1727_ ;
wire _1307_ ;
wire _4199_ ;
wire _5980_ ;
wire _5560_ ;
wire _5140_ ;
wire _638_ ;
wire _218_ ;
wire _6765_ ;
wire _6345_ ;
wire _1480_ ;
wire _1060_ ;
wire _391_ ;
wire \datapath.idinstr_24_bF$buf3  ;
wire _2685_ ;
wire _2265_ ;
wire _8911_ ;
wire _4831_ ;
wire _4411_ ;
wire _5616_ ;
wire _8088_ ;
wire \datapath.alu.b_2_bF$buf2  ;
wire _1956_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire _6994_ ;
wire _6574_ ;
wire _6154_ ;
wire _7779_ ;
wire _7359_ ;
wire _2494_ ;
wire _2074_ ;
wire _8720_ ;
wire _8300_ ;
wire _3699_ ;
wire _3279_ ;
wire _4640_ ;
wire _4220_ ;
wire _5845_ ;
wire _5425_ ;
wire _5005_ ;
wire _1765_ ;
wire _1345_ ;
wire _676_ ;
wire _256_ ;
wire _3911_ ;
wire _6383_ ;
wire _7588_ ;
wire _7168_ ;
wire _3088_ ;
wire _5510__bF$buf0 ;
wire _5510__bF$buf1 ;
wire _5510__bF$buf2 ;
wire _5510__bF$buf3 ;
wire _5510__bF$buf4 ;
wire _5510__bF$buf5 ;
wire _5510__bF$buf6 ;
wire _5510__bF$buf7 ;
wire _5654_ ;
wire _5234_ ;
wire _6859_ ;
wire _6439_ ;
wire _6019_ ;
wire _1994_ ;
wire _1574_ ;
wire _1154_ ;
wire _7800_ ;
wire _485_ ;
wire _2779_ ;
wire _2359_ ;
wire _3720_ ;
wire _3300_ ;
wire _6192_ ;
wire _4925_ ;
wire _4505_ ;
wire _7397_ ;
wire _9123_ ;
wire _5883_ ;
wire _5463_ ;
wire _5043_ ;
wire _6668_ ;
wire _6248_ ;
wire _1383_ ;
wire _294_ ;
wire _2588_ ;
wire _2168_ ;
wire \datapath.idinstr_20_hier0_bF$buf1  ;
wire _8814_ ;
wire _4734_ ;
wire _4314_ ;
wire _5939_ ;
wire _5519_ ;
wire _13_ ;
wire _1859_ ;
wire _1439_ ;
wire _1019_ ;
wire _2800_ ;
wire _5692_ ;
wire _5272_ ;
wire _6897_ ;
wire _6477_ ;
wire _6057_ ;
wire _1192_ ;
wire _2397_ ;
wire _8623_ ;
wire _8203_ ;
wire _4963_ ;
wire _4543_ ;
wire _4123_ ;
wire _5748_ ;
wire _5328_ ;
wire \datapath.alu.condtrue  ;
wire _9161_ ;
wire _1668_ ;
wire _1248_ ;
wire _5081_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire [31:0] \datapath.registers.838[20]  ;
wire \datapath.idinstr_15_bF$buf20  ;
wire _3814_ ;
wire _6286_ ;
wire _8852_ ;
wire _8432_ ;
wire _8012_ ;
wire _4772_ ;
wire _4352_ ;
wire \datapath.idinstr_21_hier0_bF$buf6  ;
wire _5977_ ;
wire _5557_ ;
wire _5137_ ;
wire _51_ ;
wire _1897_ ;
wire _1477_ ;
wire _1057_ ;
wire _7703_ ;
wire _388_ ;
wire _8908_ ;
wire _3623_ ;
wire _3203_ ;
wire _6095_ ;
wire _4828_ ;
wire _4408_ ;
wire _8661_ ;
wire _8241_ ;
wire _9026_ ;
wire _4581_ ;
wire _4161_ ;
wire _600_ ;
wire _5786_ ;
wire _5366_ ;
wire _1286_ ;
wire _7932_ ;
wire _7512_ ;
wire _197_ ;
wire _8717_ ;
wire _3852_ ;
wire _3432_ ;
wire _3012_ ;
wire _4637_ ;
wire _4217_ ;
wire _8890_ ;
wire _8470_ ;
wire _8050_ ;
wire _4390_ ;
wire _2703_ ;
wire _5595_ ;
wire _5175_ ;
wire _3908_ ;
wire _1095_ ;
wire _7741_ ;
wire _7321_ ;
wire _8946_ ;
wire _8526_ ;
wire _8106_ ;
wire _3661_ ;
wire _3241_ ;
wire _4866_ ;
wire _4446_ ;
wire _4026_ ;
wire _9064_ ;
wire _2932_ ;
wire _2512_ ;
wire _3717_ ;
wire _6189_ ;
wire _7970_ ;
wire _7550_ ;
wire _7130_ ;
wire _8755_ ;
wire _8335_ ;
wire _3890_ ;
wire _3470_ ;
wire _3050_ ;
wire _4675_ ;
wire _4255_ ;
wire _6821_ ;
wire _6401_ ;
wire _7606_ ;
wire _2741_ ;
wire _2321_ ;
wire _3946_ ;
wire _3526_ ;
wire _3106_ ;
wire _7_ ;
wire _8984_ ;
wire _8564_ ;
wire _8144_ ;
wire _4484_ ;
wire _4064_ ;
wire _923_ ;
wire _503_ ;
wire _5689_ ;
wire _5269_ ;
wire _6630_ ;
wire _6210_ ;
wire _1189_ ;
wire _7835_ ;
wire _7415_ ;
wire _2970_ ;
wire _2550_ ;
wire _2130_ ;
wire _3755_ ;
wire _3335_ ;
wire \datapath.idinstr_21_bF$buf12  ;
wire _5901_ ;
wire _8793_ ;
wire _8373_ ;
wire _1821_ ;
wire _1401_ ;
wire _9158_ ;
wire _4293_ ;
wire _732_ ;
wire _312_ ;
wire _2606_ ;
wire _5498_ ;
wire _5078_ ;
wire \datapath.idinstr_15_bF$buf17  ;
wire \datapath.idinstr_15_hier0_bF$buf5  ;
wire \datapath.idinstr_22_bF$buf21  ;
wire _7644_ ;
wire _7224_ ;
wire _8849_ ;
wire _8429_ ;
wire _8009_ ;
wire _3984_ ;
wire _3564_ ;
wire _3144_ ;
wire _4769_ ;
wire _4349_ ;
wire _5710_ ;
wire _8182_ ;
wire \datapath.idinstr_16_bF$buf26  ;
wire _48_ ;
wire _6915_ ;
wire _1630_ ;
wire _1210_ ;
wire \datapath.idinstr_20_bF$buf41  ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _2835_ ;
wire \datapath.idinstr_15_bF$buf4  ;
wire _2415_ ;
wire _7873_ ;
wire _7453_ ;
wire _7033_ ;
wire _8658_ ;
wire _8238_ ;
wire _3793_ ;
wire _3373_ ;
wire _4998_ ;
wire _4578_ ;
wire \datapath.idinstr_21_bF$buf50  ;
wire _4158_ ;
wire _6724_ ;
wire _6304_ ;
wire _770_ ;
wire _350_ ;
wire _7929_ ;
wire _7509_ ;
wire _2644_ ;
wire _2224_ ;
wire _3849_ ;
wire _3429_ ;
wire _3009_ ;
wire _7682_ ;
wire _7262_ ;
wire _8887_ ;
wire _8467_ ;
wire _8047_ ;
wire _3182_ ;
wire _1915_ ;
wire _4387_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _6953_ ;
wire _6533_ ;
wire _6113_ ;
wire _7738_ ;
wire _7318_ ;
wire _2873_ ;
wire _2453_ ;
wire _2033_ ;
wire _3658_ ;
wire _3238_ ;
wire _7491_ ;
wire _7071_ ;
wire _5804_ ;
wire _8696_ ;
wire _8276_ ;
wire [31:0] \datapath.csr._32_  ;
wire _1724_ ;
wire _1304_ ;
wire _4196_ ;
wire _635_ ;
wire _215_ ;
wire _2929_ ;
wire _2509_ ;
wire _6762_ ;
wire _6342_ ;
wire _7967_ ;
wire _7547_ ;
wire _7127_ ;
wire \datapath.idinstr_24_bF$buf0  ;
wire _2682_ ;
wire _2262_ ;
wire _3887_ ;
wire _3467_ ;
wire _3047_ ;
wire _5613_ ;
wire _8085_ ;
wire _4857__bF$buf0 ;
wire _4857__bF$buf1 ;
wire _4857__bF$buf2 ;
wire _4857__bF$buf3 ;
wire _4857__bF$buf4 ;
wire _6818_ ;
wire _1953_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire _2738_ ;
wire _2318_ ;
wire _6991_ ;
wire _6571_ ;
wire _6151_ ;
wire \controlunit.csrfile_trap_wen_bF$buf5  ;
wire _7776_ ;
wire _7356_ ;
wire _2491_ ;
wire _2071_ ;
wire \datapath.idinstr_22_bF$buf7  ;
wire _3696_ ;
wire _3276_ ;
wire _4861__bF$buf0 ;
wire _4861__bF$buf1 ;
wire _4861__bF$buf2 ;
wire _5842_ ;
wire _4861__bF$buf3 ;
wire _5422_ ;
wire _4861__bF$buf4 ;
wire _5002_ ;
wire _6627_ ;
wire _6207_ ;
wire _1762_ ;
wire _1342_ ;
wire _9099_ ;
wire _673_ ;
wire _253_ ;
wire _2967_ ;
wire _2547_ ;
wire _2127_ ;
wire _6380_ ;
wire _7585_ ;
wire _7165_ ;
wire _3085_ ;
wire _1818_ ;
wire _5651_ ;
wire _5231_ ;
wire _729_ ;
wire _309_ ;
wire _6856_ ;
wire _6436_ ;
wire _6016_ ;
wire _1991_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire \datapath.idinstr_22_bF$buf18  ;
wire _2776_ ;
wire _2356_ ;
wire _4922_ ;
wire _4502_ ;
wire _7394_ ;
wire _5707_ ;
wire _1841__bF$buf0 ;
wire _1841__bF$buf1 ;
wire _1841__bF$buf2 ;
wire _1841__bF$buf3 ;
wire _8599_ ;
wire _1841__bF$buf4 ;
wire _8179_ ;
wire _1841__bF$buf5 ;
wire _1841__bF$buf6 ;
wire _1841__bF$buf7 ;
wire _9120_ ;
wire _1627_ ;
wire _1207_ ;
wire _4099_ ;
wire _5880_ ;
wire _5460_ ;
wire _5040_ ;
wire \datapath.idinstr_20_bF$buf38  ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _6665_ ;
wire _6245_ ;
wire _1380_ ;
wire _291_ ;
wire _2585_ ;
wire _2165_ ;
wire _8811_ ;
wire _4731_ ;
wire _4311_ ;
wire \datapath.idinstr_21_bF$buf47  ;
wire _5936_ ;
wire _5516_ ;
wire _7451__bF$buf0 ;
wire _7451__bF$buf1 ;
wire _7451__bF$buf2 ;
wire _7451__bF$buf3 ;
wire _7451__bF$buf4 ;
wire _10_ ;
wire \datapath.alu.b_0_bF$buf8  ;
wire _1856_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire _6894_ ;
wire _6474_ ;
wire _6054_ ;
wire _7679_ ;
wire _7259_ ;
wire _2394_ ;
wire _8620_ ;
wire _8200_ ;
wire _3599_ ;
wire _3179_ ;
wire _4960_ ;
wire _4540_ ;
wire _4120_ ;
wire _5745_ ;
wire _5325_ ;
wire _1665_ ;
wire _1245_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _3811_ ;
wire _6283_ ;
wire \datapath.csr.mie  ;
wire _7488_ ;
wire _7068_ ;
wire \datapath.idinstr_21_hier0_bF$buf3  ;
wire _5974_ ;
wire _5554_ ;
wire _5134_ ;
wire _6759_ ;
wire _6339_ ;
wire _1894_ ;
wire _1474_ ;
wire _1054_ ;
wire _7700_ ;
wire _385_ ;
wire _2679_ ;
wire _2259_ ;
wire _8905_ ;
wire _3620_ ;
wire _3200_ ;
wire _6092_ ;
wire _4825_ ;
wire _4405_ ;
wire _7297_ ;
wire _9023_ ;
wire _5783_ ;
wire _5363_ ;
wire _6988_ ;
wire _6568_ ;
wire _6148_ ;
wire _1283_ ;
wire _194_ ;
wire _2488_ ;
wire _2068_ ;
wire _8714_ ;
wire _4634_ ;
wire _4214_ ;
wire _5839_ ;
wire _5419_ ;
wire _1759_ ;
wire _1339_ ;
wire _2700_ ;
wire _5592_ ;
wire _5172_ ;
wire _3905_ ;
wire _6797_ ;
wire _6377_ ;
wire _1092_ ;
wire _2297_ ;
wire _8943_ ;
wire _8523_ ;
wire _8103_ ;
wire _4863_ ;
wire _4443_ ;
wire _4023_ ;
wire _5648_ ;
wire _5228_ ;
wire _9061_ ;
wire _1988_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire [31:0] \datapath.registers.838[10]  ;
wire _3714_ ;
wire _6186_ ;
wire _4919_ ;
wire _8752_ ;
wire _8332_ ;
wire _9117_ ;
wire _4672_ ;
wire _4252_ ;
wire _5877_ ;
wire _5457_ ;
wire _5037_ ;
wire _1797_ ;
wire _1377_ ;
wire _7603_ ;
wire _288_ ;
wire _8808_ ;
wire _3943_ ;
wire _3523_ ;
wire _3103_ ;
wire _4_ ;
wire _4728_ ;
wire _4308_ ;
wire _8981_ ;
wire _8561_ ;
wire _8141_ ;
wire _4481_ ;
wire _4061_ ;
wire _920_ ;
wire _500_ ;
wire _5686_ ;
wire _5266_ ;
wire _1186_ ;
wire _7832_ ;
wire _7412_ ;
wire _8617_ ;
wire _3752_ ;
wire _3332_ ;
wire _4957_ ;
wire _4537_ ;
wire _4117_ ;
wire _8790_ ;
wire _8370_ ;
wire _9155_ ;
wire _4290_ ;
wire _2603_ ;
wire _5495_ ;
wire _5075_ ;
wire CLK_bF$buf140 ;
wire CLK_bF$buf141 ;
wire CLK_bF$buf142 ;
wire CLK_bF$buf143 ;
wire CLK_bF$buf144 ;
wire CLK_bF$buf145 ;
wire \datapath.idinstr_15_bF$buf14  ;
wire CLK_bF$buf146 ;
wire CLK_bF$buf147 ;
wire CLK_bF$buf148 ;
wire \datapath.csr.meta_irq  ;
wire _3808_ ;
wire CLK_bF$buf149 ;
wire \datapath.idinstr_15_hier0_bF$buf2  ;
wire _7641_ ;
wire _7221_ ;
wire _8846_ ;
wire _8426_ ;
wire _8006_ ;
wire _3981_ ;
wire _3561_ ;
wire _3141_ ;
wire _4766_ ;
wire _4346_ ;
wire \datapath.idinstr_16_bF$buf23  ;
wire _45_ ;
wire _6912_ ;
wire _2832_ ;
wire \datapath.idinstr_15_bF$buf1  ;
wire _2412_ ;
wire _4845__bF$buf0 ;
wire _4845__bF$buf1 ;
wire _4845__bF$buf2 ;
wire _4845__bF$buf3 ;
wire _4845__bF$buf4 ;
wire _3617_ ;
wire _6089_ ;
wire _7870_ ;
wire _7450_ ;
wire _7030_ ;
wire _8655_ ;
wire _8235_ ;
wire _3790_ ;
wire _3370_ ;
wire _4995_ ;
wire _4575_ ;
wire _4155_ ;
wire _6721_ ;
wire _6301_ ;
wire _7926_ ;
wire _7506_ ;
wire _2641_ ;
wire _2221_ ;
wire \datapath.idinstr_15_bF$buf52  ;
wire _3846_ ;
wire _3426_ ;
wire _3006_ ;
wire _8884_ ;
wire _8464_ ;
wire _8044_ ;
wire _1912_ ;
wire _4384_ ;
wire _823_ ;
wire _403_ ;
wire _5589_ ;
wire _5169_ ;
wire _83_ ;
wire _6950_ ;
wire _6530_ ;
wire _6110_ ;
wire _1089_ ;
wire _7735_ ;
wire _7315_ ;
wire _2870_ ;
wire _2450_ ;
wire _2030_ ;
wire _3655_ ;
wire _3235_ ;
wire _9058__bF$buf0 ;
wire _9058__bF$buf1 ;
wire _9058__bF$buf2 ;
wire _9058__bF$buf3 ;
wire _9058__bF$buf4 ;
wire _9058__bF$buf5 ;
wire _9058__bF$buf6 ;
wire _9058__bF$buf7 ;
wire _5801_ ;
wire _8693_ ;
wire _8273_ ;
wire _1721_ ;
wire _1301_ ;
wire _9058_ ;
wire _4193_ ;
wire _632_ ;
wire _212_ ;
wire _2926_ ;
wire _2506_ ;
wire _5398_ ;
wire _7964_ ;
wire _7544_ ;
wire _7124_ ;
wire \datapath.idinstr_18_bF$buf4  ;
wire [31:0] \datapath.registers.838[27]  ;
wire _8749_ ;
wire _8329_ ;
wire _3884_ ;
wire _3464_ ;
wire _3044_ ;
wire _4669_ ;
wire _4249_ ;
wire _5610_ ;
wire _8082_ ;
wire _6815_ ;
wire _1950_ ;
wire _1530_ ;
wire _1110_ ;
wire _861_ ;
wire _441_ ;
wire _2735_ ;
wire _2315_ ;
wire \controlunit.csrfile_trap_wen_bF$buf2  ;
wire _7773_ ;
wire _7353_ ;
wire \datapath.idinstr_22_bF$buf4  ;
wire _8978_ ;
wire _8558_ ;
wire _8138_ ;
wire _3693_ ;
wire _3273_ ;
wire _4898_ ;
wire _4478_ ;
wire _4058_ ;
wire _917_ ;
wire _6624_ ;
wire _6204_ ;
wire _9096_ ;
wire _670_ ;
wire _250_ ;
wire _7829_ ;
wire _7409_ ;
wire _2964_ ;
wire _2544_ ;
wire _2124_ ;
wire _3749_ ;
wire _3329_ ;
wire _7582_ ;
wire _7162_ ;
wire _8787_ ;
wire _8367_ ;
wire _3082_ ;
wire _1815_ ;
wire _4287_ ;
wire _726_ ;
wire _306_ ;
wire _6853_ ;
wire _6433_ ;
wire _6013_ ;
wire \datapath.idinstr_22_bF$buf15  ;
wire _7638_ ;
wire _7218_ ;
wire _2773_ ;
wire _2353_ ;
wire _3978_ ;
wire _3558_ ;
wire _3138_ ;
wire _7391_ ;
wire _5704_ ;
wire _8596_ ;
wire _8176_ ;
wire _6909_ ;
wire _1624_ ;
wire _1204_ ;
wire _4096_ ;
wire \datapath.idinstr_20_bF$buf35  ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _2829_ ;
wire _2409_ ;
wire _6662_ ;
wire _6242_ ;
wire _7867_ ;
wire _7447_ ;
wire _7027_ ;
wire _2582_ ;
wire _2162_ ;
wire _3787_ ;
wire _3367_ ;
wire \datapath.idinstr_21_bF$buf44  ;
wire _5933_ ;
wire _5513_ ;
wire _6718_ ;
wire \datapath.alu.b_0_bF$buf5  ;
wire _1853_ ;
wire _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _2638_ ;
wire _2218_ ;
wire _6891_ ;
wire _6471_ ;
wire _6051_ ;
wire \datapath.idinstr_15_bF$buf49  ;
wire _7676_ ;
wire _7256_ ;
wire _2391_ ;
wire _3596_ ;
wire _3176_ ;
wire _1909_ ;
wire _5742_ ;
wire _5322_ ;
wire _6947_ ;
wire _6527_ ;
wire _6107_ ;
wire _1662_ ;
wire _1242_ ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _2867_ ;
wire _2447_ ;
wire _2027_ ;
wire _9125__bF$buf0 ;
wire _9125__bF$buf1 ;
wire _9125__bF$buf2 ;
wire _9125__bF$buf3 ;
wire _9125__bF$buf4 ;
wire _6280_ ;
wire _7485_ ;
wire _7065_ ;
wire _1718_ ;
wire \datapath.idinstr_21_hier0_bF$buf0  ;
wire _5971_ ;
wire _5551_ ;
wire _5131_ ;
wire _629_ ;
wire _209_ ;
wire _6756_ ;
wire _6336_ ;
wire _1891_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _2676_ ;
wire _2256_ ;
wire _8902_ ;
wire _4822_ ;
wire _4402_ ;
wire _7294_ ;
wire _5607_ ;
wire _8499_ ;
wire _8079_ ;
wire _9020_ ;
wire _1947_ ;
wire _1527_ ;
wire [31:0] \datapath.registers.838[1]  ;
wire _1107_ ;
wire _5780_ ;
wire _5360_ ;
wire _858_ ;
wire _438_ ;
wire _6985_ ;
wire _6565_ ;
wire _6145_ ;
wire _1280_ ;
wire _191_ ;
wire _2485_ ;
wire _2065_ ;
wire _8711_ ;
wire _4631_ ;
wire _4211_ ;
wire _5836_ ;
wire _5416_ ;
wire _1756_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _3902_ ;
wire _6794_ ;
wire _6374_ ;
wire _7999_ ;
wire _7579_ ;
wire _7159_ ;
wire _2294_ ;
wire _8940_ ;
wire _8520_ ;
wire _8100_ ;
wire _3499_ ;
wire _3079_ ;
wire _4860_ ;
wire _4440_ ;
wire _4020_ ;
wire _5645_ ;
wire _5225_ ;
wire _1985_ ;
wire _1565_ ;
wire _1145_ ;
wire _896_ ;
wire _476_ ;
wire [2:0] \datapath.memexecptions  ;
wire _3711_ ;
wire _6183_ ;
wire _4916_ ;
wire _7388_ ;
wire _9114_ ;
wire _5874_ ;
wire _5454_ ;
wire _5034_ ;
wire [31:0] \datapath.alupc_4  ;
wire _6659_ ;
wire _6239_ ;
wire _1794_ ;
wire _1374_ ;
wire _7600_ ;
wire _285_ ;
wire _2999_ ;
wire _2579_ ;
wire _2159_ ;
wire _8805_ ;
wire _3940_ ;
wire _3520_ ;
wire _3100_ ;
wire [31:0] _1_ ;
wire _4725_ ;
wire _4305_ ;
wire _7197_ ;
wire _5683_ ;
wire _5263_ ;
wire _6888_ ;
wire _6468_ ;
wire _6048_ ;
wire _1183_ ;
wire _2388_ ;
wire _8614_ ;
wire _4954_ ;
wire _4534_ ;
wire _4114_ ;
wire _5739_ ;
wire _5319_ ;
wire _9152_ ;
wire _1659_ ;
wire _1239_ ;
wire _2600_ ;
wire _5492_ ;
wire _5072_ ;
wire CLK_bF$buf110 ;
wire CLK_bF$buf111 ;
wire CLK_bF$buf112 ;
wire CLK_bF$buf113 ;
wire CLK_bF$buf114 ;
wire CLK_bF$buf115 ;
wire \datapath.idinstr_15_bF$buf11  ;
wire CLK_bF$buf116 ;
wire CLK_bF$buf117 ;
wire CLK_bF$buf118 ;
wire _3805_ ;
wire CLK_bF$buf119 ;
wire _6697_ ;
wire _6277_ ;
wire _2197_ ;
wire _8843_ ;
wire _8423_ ;
wire _8003_ ;
wire _4763_ ;
wire _4343_ ;
wire _5968_ ;
wire _5548_ ;
wire _5128_ ;
wire \datapath.idinstr_16_bF$buf20  ;
wire _42_ ;
wire _1888_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _3614_ ;
wire _6086_ ;
wire _4819_ ;
wire _8652_ ;
wire _8232_ ;
wire _9017_ ;
wire _4992_ ;
wire _4572_ ;
wire _4152_ ;
wire _5777_ ;
wire _5357_ ;
wire _9190_ ;
wire _1697_ ;
wire _1277_ ;
wire _7923_ ;
wire _7503_ ;
wire _188_ ;
wire _8708_ ;
wire _3843_ ;
wire _3423_ ;
wire _3003_ ;
wire _4628_ ;
wire _4208_ ;
wire _8881_ ;
wire _8461_ ;
wire _8041_ ;
wire \datapath.idinstr_16_hier0_bF$buf4  ;
wire _4381_ ;
wire _820_ ;
wire _400_ ;
wire _5586_ ;
wire _5166_ ;
wire _80_ ;
wire _1086_ ;
wire _7732_ ;
wire _7312_ ;
wire _8937_ ;
wire _8517_ ;
wire _3652_ ;
wire _3232_ ;
wire _4857_ ;
wire _4437_ ;
wire _4017_ ;
wire _8690_ ;
wire _8270_ ;
wire _9055_ ;
wire _4190_ ;
wire _2923_ ;
wire _2503_ ;
wire _5395_ ;
wire _3708_ ;
wire _7961_ ;
wire _7541_ ;
wire _7121_ ;
wire \datapath.idinstr_18_bF$buf1  ;
wire _8746_ ;
wire _8326_ ;
wire _3881_ ;
wire _3461_ ;
wire _3041_ ;
wire _4666_ ;
wire _4246_ ;
wire _6812_ ;
wire _2732_ ;
wire _2312_ ;
wire _3937_ ;
wire _3517_ ;
wire _7770_ ;
wire _7350_ ;
wire \datapath.idinstr_22_bF$buf1  ;
wire \datapath.idinstr_16_bF$buf8  ;
wire _8975_ ;
wire _8555_ ;
wire _8135_ ;
wire _3690_ ;
wire _3270_ ;
wire _4895_ ;
wire _4475_ ;
wire _4055_ ;
wire _914_ ;
wire _6621_ ;
wire _6201_ ;
wire _9093_ ;
wire \controlunit.mret_bF$buf3  ;
wire _7826_ ;
wire _7406_ ;
wire _2961_ ;
wire _2541_ ;
wire _2121_ ;
wire _3746_ ;
wire _3326_ ;
wire \datapath.idinstr_20_bF$buf8  ;
wire _8784_ ;
wire _8364_ ;
wire _1812_ ;
wire _9149_ ;
wire _4284_ ;
wire _723_ ;
wire _303_ ;
wire _5489_ ;
wire _5069_ ;
wire _6850_ ;
wire _6430_ ;
wire _6010_ ;
wire \datapath.idinstr_22_bF$buf12  ;
wire _7635_ ;
wire _7215_ ;
wire _2770_ ;
wire _2350_ ;
wire _3975_ ;
wire _3555_ ;
wire _3135_ ;
wire _5701_ ;
wire _8593_ ;
wire _8173_ ;
wire \datapath.idinstr_16_bF$buf17  ;
wire _39_ ;
wire _6906_ ;
wire _1621_ ;
wire _1201_ ;
wire _4093_ ;
wire \datapath.idinstr_20_bF$buf32  ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _2826_ ;
wire _2406_ ;
wire \controlunit.csrfile_wen  ;
wire _5298_ ;
wire [31:0] \datapath.regcsralu  ;
wire _7864_ ;
wire _7444_ ;
wire _7024_ ;
wire [31:0] \datapath.registers.838[17]  ;
wire _8649_ ;
wire _8229_ ;
wire _3784_ ;
wire _3364_ ;
wire _4989_ ;
wire _4569_ ;
wire \datapath.idinstr_21_bF$buf41  ;
wire _4149_ ;
wire _5930_ ;
wire _5510_ ;
wire _6715_ ;
wire \datapath.alu.b_0_bF$buf2  ;
wire _1850_ ;
wire _1430_ ;
wire _1010_ ;
wire _9187_ ;
wire _761_ ;
wire _341_ ;
wire _2635_ ;
wire _2215_ ;
wire _2870__bF$buf0 ;
wire _2870__bF$buf1 ;
wire _2870__bF$buf2 ;
wire _2870__bF$buf3 ;
wire _2870__bF$buf4 ;
wire _2870__bF$buf5 ;
wire _2870__bF$buf6 ;
wire \datapath.idinstr_15_bF$buf46  ;
wire _7673_ ;
wire _7253_ ;
wire _8878_ ;
wire _8458_ ;
wire _8038_ ;
wire _3593_ ;
wire _3173_ ;
wire _1906_ ;
wire _4798_ ;
wire _4378_ ;
wire _817_ ;
wire _77_ ;
wire _6944_ ;
wire _6524_ ;
wire _6104_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _7729_ ;
wire _7309_ ;
wire _2864_ ;
wire _2444_ ;
wire _2024_ ;
wire _3649_ ;
wire _3229_ ;
wire _7482_ ;
wire _7062_ ;
wire _8687_ ;
wire _8267_ ;
wire _1715_ ;
wire _4187_ ;
wire _626_ ;
wire _206_ ;
wire _6753_ ;
wire _6333_ ;
wire _7958_ ;
wire _7538_ ;
wire _7118_ ;
wire _2673_ ;
wire _2253_ ;
wire _3878_ ;
wire _3458_ ;
wire _3038_ ;
wire _7291_ ;
wire _5604_ ;
wire _8496_ ;
wire _8076_ ;
wire _6809_ ;
wire _1944_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire _2729_ ;
wire _2309_ ;
wire _6982_ ;
wire _6562_ ;
wire _6142_ ;
wire \datapath.alu.b_3_bF$buf5  ;
wire _7767_ ;
wire _7347_ ;
wire _2482_ ;
wire _2062_ ;
wire _3687_ ;
wire _3267_ ;
wire _5833_ ;
wire _5413_ ;
wire _6618_ ;
wire _1753_ ;
wire _1333_ ;
wire _664_ ;
wire _244_ ;
wire _2958_ ;
wire _2538_ ;
wire _2118_ ;
wire _6791_ ;
wire _6371_ ;
wire _7996_ ;
wire _7576_ ;
wire _7156_ ;
wire _2291_ ;
wire _3496_ ;
wire _3076_ ;
wire _1809_ ;
wire _5642_ ;
wire _5222_ ;
wire _6847_ ;
wire _6427_ ;
wire _6007_ ;
wire _1982_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _2767_ ;
wire _2347_ ;
wire _6180_ ;
wire _4913_ ;
wire _7385_ ;
wire _9111_ ;
wire _1618_ ;
wire _5871_ ;
wire _5451_ ;
wire _5031_ ;
wire \datapath.idinstr_20_bF$buf29  ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _6656_ ;
wire _6236_ ;
wire _1791_ ;
wire _1371_ ;
wire _282_ ;
wire _2996_ ;
wire _2576_ ;
wire _2156_ ;
wire _8802_ ;
wire _4722_ ;
wire _4302_ ;
wire _7194_ ;
wire \datapath.idinstr_21_bF$buf38  ;
wire _5927_ ;
wire _5507_ ;
wire _8399_ ;
wire _1847_ ;
wire _1427_ ;
wire _1007_ ;
wire _5680_ ;
wire _5260_ ;
wire _758_ ;
wire _338_ ;
wire _6885_ ;
wire _6465_ ;
wire _6045_ ;
wire _1180_ ;
wire \datapath.idinstr_22_hier0_bF$buf4  ;
wire _2385_ ;
wire _8611_ ;
wire _4951_ ;
wire _4531_ ;
wire _4111_ ;
wire _5736_ ;
wire _5316_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _3802_ ;
wire _6694_ ;
wire _6274_ ;
wire _7899_ ;
wire _7479_ ;
wire _7059_ ;
wire _2194_ ;
wire _8840_ ;
wire _8420_ ;
wire _8000_ ;
wire _3399_ ;
wire _4760_ ;
wire _4340_ ;
wire _5965_ ;
wire _5545_ ;
wire _5125_ ;
wire _1885_ ;
wire _1465_ ;
wire _1045_ ;
wire _796_ ;
wire _376_ ;
wire _3611_ ;
wire _6083_ ;
wire _4816_ ;
wire _7288_ ;
wire _9014_ ;
wire _5774_ ;
wire _5354_ ;
wire CLK_bF$buf0 ;
wire CLK_bF$buf1 ;
wire CLK_bF$buf2 ;
wire CLK_bF$buf3 ;
wire CLK_bF$buf4 ;
wire CLK_bF$buf5 ;
wire CLK_bF$buf6 ;
wire CLK_bF$buf7 ;
wire CLK_bF$buf8 ;
wire CLK_bF$buf9 ;
wire _6979_ ;
wire _6559_ ;
wire _6139_ ;
wire _1694_ ;
wire _1274_ ;
wire _4934__bF$buf0 ;
wire _4934__bF$buf1 ;
wire _4934__bF$buf2 ;
wire _7920_ ;
wire _4934__bF$buf3 ;
wire _7500_ ;
wire _4934__bF$buf4 ;
wire _4934__bF$buf5 ;
wire _4934__bF$buf6 ;
wire _4934__bF$buf7 ;
wire _4934__bF$buf8 ;
wire _4934__bF$buf9 ;
wire _185_ ;
wire _2899_ ;
wire _2479_ ;
wire _2059_ ;
wire _8705_ ;
wire _3840_ ;
wire _3420_ ;
wire _3000_ ;
wire _4625_ ;
wire _4205_ ;
wire _7097_ ;
wire \datapath.idinstr_16_hier0_bF$buf1  ;
wire _5583_ ;
wire _5163_ ;
wire _6788_ ;
wire _6368_ ;
wire _1083_ ;
wire _2288_ ;
wire _8934_ ;
wire _8514_ ;
wire _4854_ ;
wire _4434_ ;
wire _4014_ ;
wire _5639_ ;
wire _5219_ ;
wire _9052_ ;
wire _1979_ ;
wire _1559_ ;
wire _1139_ ;
wire _2920_ ;
wire _2500_ ;
wire _5392_ ;
wire _3705_ ;
wire _6597_ ;
wire _6177_ ;
wire _2097_ ;
wire _8743_ ;
wire _8323_ ;
wire _9108_ ;
wire _4663_ ;
wire _4243_ ;
wire _5868_ ;
wire _5448_ ;
wire _5028_ ;
wire _1788_ ;
wire _1368_ ;
wire _699_ ;
wire _279_ ;
wire _3934_ ;
wire _3514_ ;
wire _4719_ ;
wire \datapath.idinstr_16_bF$buf5  ;
wire _8972_ ;
wire _8552_ ;
wire _8132_ ;
wire _4892_ ;
wire _4472_ ;
wire _4052_ ;
wire _5755__bF$buf0 ;
wire _5755__bF$buf1 ;
wire _5755__bF$buf2 ;
wire _5755__bF$buf3 ;
wire _5755__bF$buf4 ;
wire _911_ ;
wire _5677_ ;
wire _5257_ ;
wire _9090_ ;
wire \controlunit.mret_bF$buf0  ;
wire _1597_ ;
wire [31:0] \datapath.registers.838[8]  ;
wire _1177_ ;
wire _7823_ ;
wire _7403_ ;
wire _8608_ ;
wire _3743_ ;
wire _3323_ ;
wire _4948_ ;
wire \datapath.idinstr_20_bF$buf5  ;
wire _4528_ ;
wire _4108_ ;
wire _8781_ ;
wire _8361_ ;
wire _9146_ ;
wire _4281_ ;
wire _720_ ;
wire _300_ ;
wire _5486_ ;
wire _5066_ ;
wire _7632_ ;
wire _7212_ ;
wire _8837_ ;
wire _8417_ ;
wire _3972_ ;
wire _3552_ ;
wire _3132_ ;
wire _4757_ ;
wire _4337_ ;
wire _8590_ ;
wire _8170_ ;
wire \datapath.idinstr_16_bF$buf14  ;
wire _36_ ;
wire _6903_ ;
wire _4090_ ;
wire _2823_ ;
wire _2403_ ;
wire _5295_ ;
wire _3608_ ;
wire _7861_ ;
wire _7441_ ;
wire _7021_ ;
wire _8646_ ;
wire _8226_ ;
wire _3781_ ;
wire _3361_ ;
wire _4986_ ;
wire _4566_ ;
wire _4146_ ;
wire _4855__bF$buf0 ;
wire _4855__bF$buf1 ;
wire _4855__bF$buf2 ;
wire _4855__bF$buf3 ;
wire _4855__bF$buf4 ;
wire _6712_ ;
wire _9184_ ;
wire _7917_ ;
wire _2632_ ;
wire _2212_ ;
wire \datapath.idinstr_15_bF$buf43  ;
wire _3837_ ;
wire _3417_ ;
wire _7670_ ;
wire _7250_ ;
wire _8875_ ;
wire _8455_ ;
wire _8035_ ;
wire _3590_ ;
wire _3170_ ;
wire _1903_ ;
wire _4795_ ;
wire _4375_ ;
wire _814_ ;
wire _74_ ;
wire _6941_ ;
wire _6521_ ;
wire _6101_ ;
wire _7726_ ;
wire _7306_ ;
wire _2861_ ;
wire _2441_ ;
wire _2021_ ;
wire _3646_ ;
wire _3226_ ;
wire _5085__bF$buf0 ;
wire _5085__bF$buf1 ;
wire _5085__bF$buf2 ;
wire _5085__bF$buf3 ;
wire _5085__bF$buf4 ;
wire _5085__bF$buf5 ;
wire _5085__bF$buf6 ;
wire _5085__bF$buf7 ;
wire _8684_ ;
wire _8264_ ;
wire _1712_ ;
wire _9049_ ;
wire _4184_ ;
wire _623_ ;
wire _203_ ;
wire _2917_ ;
wire _5389_ ;
wire _6750_ ;
wire _6330_ ;
wire _7955_ ;
wire _7535_ ;
wire _7115_ ;
wire _2670_ ;
wire _2250_ ;
wire _3875_ ;
wire _3455_ ;
wire _3035_ ;
wire _5601_ ;
wire _8493_ ;
wire _8073_ ;
wire _6806_ ;
wire _1941_ ;
wire _1521_ ;
wire _1101_ ;
wire _852_ ;
wire _432_ ;
wire _2726_ ;
wire _2306_ ;
wire _5198_ ;
wire \datapath.alu.b_3_bF$buf2  ;
wire _7764_ ;
wire _7344_ ;
wire _8969_ ;
wire _8549_ ;
wire _8129_ ;
wire _3684_ ;
wire _3264_ ;
wire _4889_ ;
wire _4469_ ;
wire _4049_ ;
wire _5830_ ;
wire _5410_ ;
wire _908_ ;
wire _6615_ ;
wire _1750_ ;
wire _1330_ ;
wire _9087_ ;
wire _661_ ;
wire _241_ ;
wire _2955_ ;
wire _2535_ ;
wire _2115_ ;
wire _7993_ ;
wire _7573_ ;
wire _7153_ ;
wire _388__bF$buf0 ;
wire _388__bF$buf1 ;
wire _388__bF$buf2 ;
wire _388__bF$buf3 ;
wire _388__bF$buf4 ;
wire _8778_ ;
wire _8358_ ;
wire _3493_ ;
wire _3073_ ;
wire _1806_ ;
wire _4698_ ;
wire _4278_ ;
wire _717_ ;
wire _6844_ ;
wire _6424_ ;
wire _6004_ ;
wire _890_ ;
wire _470_ ;
wire _7629_ ;
wire _7209_ ;
wire _2764_ ;
wire _2344_ ;
wire _3969_ ;
wire _3549_ ;
wire _3129_ ;
wire _4910_ ;
wire _7382_ ;
wire _8587_ ;
wire _8167_ ;
wire _1615_ ;
wire _4087_ ;
wire \datapath.idinstr_20_bF$buf26  ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _6653_ ;
wire _6233_ ;
wire _7858_ ;
wire _7438_ ;
wire _7018_ ;
wire _2993_ ;
wire _2573_ ;
wire _2153_ ;
wire _3778_ ;
wire _3358_ ;
wire _7191_ ;
wire \datapath.idinstr_21_bF$buf35  ;
wire _5924_ ;
wire _5504_ ;
wire _8396_ ;
wire _6709_ ;
wire _1844_ ;
wire _1424_ ;
wire _1004_ ;
wire _755_ ;
wire _335_ ;
wire _2629_ ;
wire _2209_ ;
wire _6882_ ;
wire _6462_ ;
wire _6042_ ;
wire \datapath.idinstr_22_hier0_bF$buf1  ;
wire _7667_ ;
wire _7247_ ;
wire _2382_ ;
wire _3587_ ;
wire _3167_ ;
wire _5733_ ;
wire _5313_ ;
wire \datapath.idinstr_16_bF$buf49  ;
wire _6938_ ;
wire _6518_ ;
wire _1653_ ;
wire _1233_ ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _2858_ ;
wire _2438_ ;
wire _2018_ ;
wire _6691_ ;
wire _6271_ ;
wire _7896_ ;
wire _7476_ ;
wire _7056_ ;
wire _2191_ ;
wire _5762__bF$buf20 ;
wire _5762__bF$buf21 ;
wire _5762__bF$buf22 ;
wire _5762__bF$buf23 ;
wire _5762__bF$buf24 ;
wire _5762__bF$buf25 ;
wire _5762__bF$buf26 ;
wire _5762__bF$buf27 ;
wire _5762__bF$buf28 ;
wire _5762__bF$buf29 ;
wire _3396_ ;
wire _1709_ ;
wire _5962_ ;
wire _5542_ ;
wire _5122_ ;
wire _6747_ ;
wire _6327_ ;
wire _1882_ ;
wire _1462_ ;
wire _1042_ ;
wire _793_ ;
wire _373_ ;
wire _2667_ ;
wire _2247_ ;
wire _6080_ ;
wire _4813_ ;
wire _7285_ ;
wire _4803__bF$buf0 ;
wire _4803__bF$buf1 ;
wire _4803__bF$buf2 ;
wire _4803__bF$buf3 ;
wire _4803__bF$buf4 ;
wire _9011_ ;
wire _1938_ ;
wire _1518_ ;
wire _5771_ ;
wire _5351_ ;
wire _849_ ;
wire _429_ ;
wire _6976_ ;
wire _6556_ ;
wire _6136_ ;
wire _1691_ ;
wire _1271_ ;
wire _182_ ;
wire _2896_ ;
wire _2476_ ;
wire _2056_ ;
wire _8702_ ;
wire _4622_ ;
wire _4202_ ;
wire _7094_ ;
wire _5827_ ;
wire _5407_ ;
wire _8299_ ;
wire _1747_ ;
wire _1327_ ;
wire _5580_ ;
wire _5160_ ;
wire _658_ ;
wire _238_ ;
wire _9091__bF$buf0 ;
wire _9091__bF$buf1 ;
wire _9091__bF$buf2 ;
wire _9091__bF$buf3 ;
wire _9091__bF$buf4 ;
wire _6785_ ;
wire _6365_ ;
wire _1080_ ;
wire _2285_ ;
wire _8931_ ;
wire _8511_ ;
wire _4851_ ;
wire _4431_ ;
wire _4011_ ;
wire _5636_ ;
wire _5216_ ;
wire _3410__bF$buf0 ;
wire _3410__bF$buf1 ;
wire _3410__bF$buf2 ;
wire _3410__bF$buf3 ;
wire _1976_ ;
wire _1556_ ;
wire _1136_ ;
wire _7425__bF$buf30 ;
wire _7425__bF$buf31 ;
wire _7425__bF$buf32 ;
wire _7425__bF$buf33 ;
wire _7425__bF$buf34 ;
wire _7425__bF$buf35 ;
wire _7425__bF$buf36 ;
wire _7425__bF$buf37 ;
wire _7425__bF$buf38 ;
wire _7425__bF$buf39 ;
wire _887_ ;
wire _467_ ;
wire _3702_ ;
wire _6594_ ;
wire _6174_ ;
wire _4907_ ;
wire _7799_ ;
wire _7379_ ;
wire _2094_ ;
wire _8740_ ;
wire _8320_ ;
wire _3299_ ;
wire _9105_ ;
wire _4660_ ;
wire _4240_ ;
wire _5865_ ;
wire _5445_ ;
wire _5025_ ;
wire [31:0] \datapath.idpc  ;
wire _1785_ ;
wire _1365_ ;
wire _696_ ;
wire _276_ ;
wire _3931_ ;
wire _3511_ ;
wire _4716_ ;
wire _7188_ ;
wire \datapath.idinstr_16_bF$buf2  ;
wire _5674_ ;
wire _5254_ ;
wire _6879_ ;
wire _6459_ ;
wire _6039_ ;
wire _1594_ ;
wire _1174_ ;
wire _7820_ ;
wire _7400_ ;
wire _2799_ ;
wire _2379_ ;
wire _8605_ ;
wire _3740_ ;
wire _3320_ ;
wire _4945_ ;
wire \datapath.idinstr_20_bF$buf2  ;
wire _4525_ ;
wire _4105_ ;
wire [1:0] \datapath.regpcsel  ;
wire _9143_ ;
wire _5483_ ;
wire _5063_ ;
wire _6688_ ;
wire _6268_ ;
wire _2188_ ;
wire _8834_ ;
wire _8414_ ;
wire _4754_ ;
wire _4334_ ;
wire _5959_ ;
wire _5539_ ;
wire _5119_ ;
wire \datapath.idinstr_16_bF$buf11  ;
wire _33_ ;
wire _6900_ ;
wire _1879_ ;
wire _1459_ ;
wire _1039_ ;
wire _2820_ ;
wire _2400_ ;
wire _5292_ ;
wire _3605_ ;
wire _6497_ ;
wire _6077_ ;
wire _8643_ ;
wire _8223_ ;
wire _9008_ ;
wire _4983_ ;
wire _4563_ ;
wire _4143_ ;
wire \datapath.idinstr_19_bF$buf5  ;
wire _5768_ ;
wire _5348_ ;
wire _9181_ ;
wire _1688_ ;
wire _1268_ ;
wire _7914_ ;
wire _599_ ;
wire _179_ ;
wire [31:0] \datapath.registers.838[22]  ;
wire \datapath.idinstr_15_bF$buf40  ;
wire _3834_ ;
wire _3414_ ;
wire _4619_ ;
wire _8872_ ;
wire _8452_ ;
wire _8032_ ;
wire _1900_ ;
wire _4792_ ;
wire _4372_ ;
wire \datapath.idinstr_23_bF$buf5  ;
wire _811_ ;
wire _5997_ ;
wire _5577_ ;
wire _5157_ ;
wire _71_ ;
wire _5762__bF$buf0 ;
wire _5762__bF$buf1 ;
wire _5762__bF$buf2 ;
wire _5762__bF$buf3 ;
wire _5762__bF$buf4 ;
wire _5762__bF$buf5 ;
wire _5762__bF$buf6 ;
wire _5762__bF$buf7 ;
wire _1497_ ;
wire _5762__bF$buf8 ;
wire _1077_ ;
wire _5762__bF$buf9 ;
wire _7723_ ;
wire _7303_ ;
wire _8928_ ;
wire _8508_ ;
wire _3643_ ;
wire _3223_ ;
wire _4848_ ;
wire _4428_ ;
wire _4008_ ;
wire _8681_ ;
wire _8261_ ;
wire [31:0] \datapath.csr.csr_data  ;
wire _9046_ ;
wire _4181_ ;
wire _620_ ;
wire _200_ ;
wire _2914_ ;
wire _5386_ ;
wire _7952_ ;
wire _7532_ ;
wire _7112_ ;
wire _8737_ ;
wire _8317_ ;
wire _3872_ ;
wire _3452_ ;
wire _3032_ ;
wire _4657_ ;
wire _4237_ ;
wire _8490_ ;
wire _8070_ ;
wire _6803_ ;
wire _2723_ ;
wire _2303_ ;
wire _5195_ ;
wire _3928_ ;
wire _3508_ ;
wire _7761_ ;
wire _7341_ ;
wire _8966_ ;
wire _8546_ ;
wire _8126_ ;
wire _3681_ ;
wire _3261_ ;
wire _4886_ ;
wire _4466_ ;
wire _4046_ ;
wire _905_ ;
wire _6612_ ;
wire _9084_ ;
wire _7817_ ;
wire _2952_ ;
wire _2532_ ;
wire _2112_ ;
wire _3737_ ;
wire _3317_ ;
wire \datapath.alu.b_1_bF$buf6  ;
wire _7990_ ;
wire _7570_ ;
wire _7150_ ;
wire _8775_ ;
wire _8355_ ;
wire _3490_ ;
wire _3070_ ;
wire _1803_ ;
wire _4695_ ;
wire _4275_ ;
wire _714_ ;
wire _6841_ ;
wire _6421_ ;
wire _6001_ ;
wire [31:0] \datapath.alu.c  ;
wire _7626_ ;
wire _7206_ ;
wire _2761_ ;
wire _2341_ ;
wire _3966_ ;
wire _3546_ ;
wire _3126_ ;
wire _8584_ ;
wire _8164_ ;
wire _1612_ ;
wire _4084_ ;
wire \datapath.idinstr_20_bF$buf23  ;
wire _943_ ;
wire _523_ ;
wire _103_ ;
wire _2817_ ;
wire _5289_ ;
wire _6650_ ;
wire _6230_ ;
wire _7855_ ;
wire _7435_ ;
wire _7015_ ;
wire _2990_ ;
wire _2570_ ;
wire _2150_ ;
wire _3775_ ;
wire _3355_ ;
wire _3563__bF$buf0 ;
wire _3563__bF$buf1 ;
wire _3563__bF$buf2 ;
wire \datapath.idinstr_21_bF$buf32  ;
wire _3563__bF$buf3 ;
wire _3563__bF$buf4 ;
wire _5921_ ;
wire _5501_ ;
wire _5017__bF$buf0 ;
wire _5017__bF$buf1 ;
wire _5017__bF$buf2 ;
wire _5017__bF$buf3 ;
wire _5017__bF$buf4 ;
wire _8393_ ;
wire _5017__bF$buf5 ;
wire _5017__bF$buf6 ;
wire _5017__bF$buf7 ;
wire _6706_ ;
wire _1841_ ;
wire _1421_ ;
wire _1001_ ;
wire _9178_ ;
wire _752_ ;
wire _332_ ;
wire _2626_ ;
wire _2206_ ;
wire _5098_ ;
wire \datapath.idinstr_15_bF$buf37  ;
wire \datapath.idinstr_22_bF$buf41  ;
wire _7664_ ;
wire _7244_ ;
wire _8869_ ;
wire _8449_ ;
wire _8029_ ;
wire _3584_ ;
wire _3164_ ;
wire _4789_ ;
wire _4369_ ;
wire _5730_ ;
wire _5310_ ;
wire _808_ ;
wire \datapath.idinstr_16_bF$buf46  ;
wire _68_ ;
wire _6935_ ;
wire _6515_ ;
wire _1650_ ;
wire _1230_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _2855_ ;
wire _2435_ ;
wire _2015_ ;
wire _7893_ ;
wire _7473_ ;
wire _7053_ ;
wire _8678_ ;
wire _8258_ ;
wire _3393_ ;
wire _1706_ ;
wire _4598_ ;
wire _4178_ ;
wire _617_ ;
wire _6744_ ;
wire _6324_ ;
wire _790_ ;
wire _370_ ;
wire _7949_ ;
wire _7529_ ;
wire _7109_ ;
wire _2664_ ;
wire _2244_ ;
wire _3869_ ;
wire _3449_ ;
wire _3029_ ;
wire _4810_ ;
wire _7282_ ;
wire _8487_ ;
wire _8067_ ;
wire _1935_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _6973_ ;
wire _6553_ ;
wire _6133_ ;
wire _7758_ ;
wire _7338_ ;
wire _2893_ ;
wire _2473_ ;
wire _2053_ ;
wire _3678_ ;
wire _3258_ ;
wire _7091_ ;
wire _5824_ ;
wire _5404_ ;
wire _8296_ ;
wire _6609_ ;
wire _1744_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _2949_ ;
wire _2529_ ;
wire _2109_ ;
wire _6782_ ;
wire _6362_ ;
wire _7987_ ;
wire _7567_ ;
wire _7147_ ;
wire _2282_ ;
wire _3487_ ;
wire _3067_ ;
wire _182__bF$buf0 ;
wire _182__bF$buf1 ;
wire _182__bF$buf2 ;
wire _182__bF$buf3 ;
wire _182__bF$buf4 ;
wire _5633_ ;
wire _5213_ ;
wire _6838_ ;
wire _6418_ ;
wire _1973_ ;
wire _1553_ ;
wire _1133_ ;
wire _884_ ;
wire _464_ ;
wire _2758_ ;
wire _2338_ ;
wire _6591_ ;
wire _6171_ ;
wire _4904_ ;
wire _7796_ ;
wire _7376_ ;
wire _2091_ ;
wire \datapath.regz  ;
wire _3296_ ;
wire _9102_ ;
wire _1609_ ;
wire _5862_ ;
wire _5442_ ;
wire _5022_ ;
wire _6647_ ;
wire _6227_ ;
wire _1782_ ;
wire _1362_ ;
wire _693_ ;
wire _273_ ;
wire _2987_ ;
wire _2567_ ;
wire _2147_ ;
wire _4713_ ;
wire _7185_ ;
wire \datapath.idinstr_21_bF$buf29  ;
wire _5918_ ;
wire _1838_ ;
wire _1418_ ;
wire _5671_ ;
wire _5251_ ;
wire _749_ ;
wire _329_ ;
wire _6876_ ;
wire _6456_ ;
wire _6036_ ;
wire _1591_ ;
wire _1171_ ;
wire \datapath.idinstr_22_bF$buf38  ;
wire _2796_ ;
wire _2376_ ;
wire _8602_ ;
wire _4942_ ;
wire _4522_ ;
wire _4102_ ;
wire _5727_ ;
wire _5307_ ;
wire _8199_ ;
wire _9140_ ;
wire _1647_ ;
wire _1227_ ;
wire _5480_ ;
wire _5060_ ;
wire _978_ ;
wire _558_ ;
wire _138_ ;
wire _6685_ ;
wire _6265_ ;
wire _2185_ ;
wire _8831_ ;
wire _8411_ ;
wire _4751_ ;
wire _4331_ ;
wire _5956_ ;
wire _5536_ ;
wire _5116_ ;
wire _30_ ;
wire _1876_ ;
wire _1456_ ;
wire _1036_ ;
wire _787_ ;
wire _367_ ;
wire _3602_ ;
wire _6494_ ;
wire _6074_ ;
wire _4807_ ;
wire _7699_ ;
wire _7279_ ;
wire _8640_ ;
wire _8220_ ;
wire _2016__bF$buf0 ;
wire _2016__bF$buf1 ;
wire _2016__bF$buf2 ;
wire _2016__bF$buf3 ;
wire _3199_ ;
wire _9005_ ;
wire _4980_ ;
wire _4560_ ;
wire _4140_ ;
wire \datapath.idinstr_19_bF$buf2  ;
wire _5765_ ;
wire _5345_ ;
wire _1685_ ;
wire _1265_ ;
wire _7911_ ;
wire _596_ ;
wire _176_ ;
wire _3831_ ;
wire _3411_ ;
wire _4616_ ;
wire _7088_ ;
wire \datapath.idinstr_23_bF$buf2  ;
wire _5994_ ;
wire _5574_ ;
wire _5154_ ;
wire [31:0] \datapath.programcounter.pc_mux  ;
wire _6779_ ;
wire _6359_ ;
wire _1494_ ;
wire _1074_ ;
wire _7720_ ;
wire _7300_ ;
wire _2699_ ;
wire _2279_ ;
wire _8925_ ;
wire _8505_ ;
wire _3640_ ;
wire _3220_ ;
wire [31:0] \datapath.csr.csr_mepc  ;
wire _4845_ ;
wire _4425_ ;
wire _4005_ ;
wire _9043_ ;
wire _2911_ ;
wire _5383_ ;
wire _6588_ ;
wire _6168_ ;
wire _2088_ ;
wire _8734_ ;
wire _8314_ ;
wire _4654_ ;
wire _4234_ ;
wire _5859_ ;
wire _5439_ ;
wire _5019_ ;
wire _6800_ ;
wire _1779_ ;
wire _1359_ ;
wire _2720_ ;
wire _2300_ ;
wire _5192_ ;
wire _3925_ ;
wire _3505_ ;
wire _6397_ ;
wire _8963_ ;
wire _8543_ ;
wire _8123_ ;
wire _4883_ ;
wire _4463_ ;
wire _4043_ ;
wire _902_ ;
wire _5668_ ;
wire _5248_ ;
wire _9081_ ;
wire _1588_ ;
wire _1168_ ;
wire _7814_ ;
wire _499_ ;
wire [31:0] \datapath.registers.838[12]  ;
wire _3734_ ;
wire _3314_ ;
wire \datapath.alu.b_1_bF$buf3  ;
wire _4939_ ;
wire _4519_ ;
wire _8772_ ;
wire _8352_ ;
wire _1800_ ;
wire _9137_ ;
wire _4692_ ;
wire _4272_ ;
wire _711_ ;
wire _5897_ ;
wire _5477_ ;
wire _5057_ ;
wire _1397_ ;
wire _7623_ ;
wire _7203_ ;
wire _8828_ ;
wire _8408_ ;
wire _3963_ ;
wire _3543_ ;
wire _3123_ ;
wire _4748_ ;
wire _4328_ ;
wire _8581_ ;
wire _8161_ ;
wire _27_ ;
wire _4081_ ;
wire \datapath.idinstr_20_bF$buf20  ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire _2814_ ;
wire _5286_ ;
wire _7852_ ;
wire _7432_ ;
wire _7012_ ;
wire _8637_ ;
wire _8217_ ;
wire _3772_ ;
wire _3352_ ;
wire \datapath.idinstr_17_bF$buf14  ;
wire _4977_ ;
wire _4557_ ;
wire _4137_ ;
wire _8390_ ;
wire _6703_ ;
wire _9175_ ;
wire _7908_ ;
wire _2623_ ;
wire _2203_ ;
wire _5095_ ;
wire \datapath.idinstr_15_bF$buf34  ;
wire _3828_ ;
wire _3408_ ;
wire _7661_ ;
wire _7241_ ;
wire _8866_ ;
wire _8446_ ;
wire _8026_ ;
wire _3581_ ;
wire _3161_ ;
wire _4786_ ;
wire _4366_ ;
wire _805_ ;
wire \datapath.idinstr_16_bF$buf43  ;
wire _65_ ;
wire _6932_ ;
wire _6512_ ;
wire _7717_ ;
wire _2852_ ;
wire _2432_ ;
wire _2012_ ;
wire _3637_ ;
wire _3217_ ;
wire _7890_ ;
wire _7470_ ;
wire _7050_ ;
wire _8675_ ;
wire _8255_ ;
wire _3390_ ;
wire _1703_ ;
wire _4595_ ;
wire _4175_ ;
wire _614_ ;
wire _2908_ ;
wire _6741_ ;
wire _6321_ ;
wire _7946_ ;
wire _7526_ ;
wire _7106_ ;
wire _2661_ ;
wire _2241_ ;
wire _3866_ ;
wire _3446_ ;
wire _3026_ ;
wire _8484_ ;
wire _8064_ ;
wire _1932_ ;
wire _1512_ ;
wire _843_ ;
wire _423_ ;
wire _2717_ ;
wire _5189_ ;
wire _6970_ ;
wire _6550_ ;
wire _6130_ ;
wire _7755_ ;
wire _7335_ ;
wire _2890_ ;
wire _2470_ ;
wire _2050_ ;
wire _3675_ ;
wire _3255_ ;
wire _5821_ ;
wire _5401_ ;
wire _8293_ ;
wire _6606_ ;
wire _1741_ ;
wire _1321_ ;
wire _9078_ ;
wire _652_ ;
wire _232_ ;
wire _2946_ ;
wire _2526_ ;
wire _2106_ ;
wire _7984_ ;
wire _7564_ ;
wire _7144_ ;
wire [31:0] \datapath.registers.838[29]  ;
wire _8769_ ;
wire _8349_ ;
wire _3484_ ;
wire _3064_ ;
wire _4689_ ;
wire _4269_ ;
wire _5630_ ;
wire _5210_ ;
wire _708_ ;
wire _6835_ ;
wire _6415_ ;
wire _1970_ ;
wire _1550_ ;
wire _1130_ ;
wire _881_ ;
wire _461_ ;
wire _2755_ ;
wire _2335_ ;
wire [3:0] alusel ;
wire _4901_ ;
wire _7793_ ;
wire _7373_ ;
wire _8998_ ;
wire _8578_ ;
wire _8158_ ;
wire _3293_ ;
wire _1606_ ;
wire _4498_ ;
wire _4078_ ;
wire \datapath.idinstr_20_bF$buf17  ;
wire _937_ ;
wire _517_ ;
wire _6644_ ;
wire _6224_ ;
wire _690_ ;
wire _270_ ;
wire _7849_ ;
wire _7429_ ;
wire _7009_ ;
wire _2984_ ;
wire _2564_ ;
wire _2144_ ;
wire _3769_ ;
wire _3349_ ;
wire _4710_ ;
wire _7182_ ;
wire \datapath.idinstr_21_bF$buf26  ;
wire _5915_ ;
wire _8387_ ;
wire _1835_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _6873_ ;
wire _6453_ ;
wire _6033_ ;
wire \datapath.idinstr_22_bF$buf35  ;
wire _7658_ ;
wire _7238_ ;
wire _2793_ ;
wire _2373_ ;
wire _3998_ ;
wire _3578_ ;
wire _3158_ ;
wire _5724_ ;
wire _5304_ ;
wire _8196_ ;
wire _6929_ ;
wire _6509_ ;
wire _1644_ ;
wire _1224_ ;
wire \datapath.idinstr_20_bF$buf55  ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire _2849_ ;
wire _2429_ ;
wire _2009_ ;
wire _6682_ ;
wire _6262_ ;
wire _7887_ ;
wire _7467_ ;
wire _7047_ ;
wire _2182_ ;
wire _3387_ ;
wire _5953_ ;
wire _5533_ ;
wire _5113_ ;
wire DMEM_WEN ;
wire _6738_ ;
wire _6318_ ;
wire _1873_ ;
wire _1453_ ;
wire _1033_ ;
wire _784_ ;
wire _364_ ;
wire _2658_ ;
wire _2238_ ;
wire _6491_ ;
wire _6071_ ;
wire _4809__bF$buf0 ;
wire _4809__bF$buf1 ;
wire _4809__bF$buf2 ;
wire _4809__bF$buf3 ;
wire _4809__bF$buf4 ;
wire _4804_ ;
wire _7696_ ;
wire _7276_ ;
wire _3196_ ;
wire _9002_ ;
wire _1929_ ;
wire _1509_ ;
wire _5762_ ;
wire _5342_ ;
wire _6967_ ;
wire _6547_ ;
wire _6127_ ;
wire _1682_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _2887_ ;
wire _2467_ ;
wire _2047_ ;
wire _4813__bF$buf0 ;
wire _4813__bF$buf1 ;
wire _4813__bF$buf2 ;
wire _4813__bF$buf3 ;
wire _4813__bF$buf4 ;
wire _4613_ ;
wire _7085_ ;
wire _5818_ ;
wire _1738_ ;
wire _1318_ ;
wire _5991_ ;
wire _5571_ ;
wire _5151_ ;
wire _649_ ;
wire _229_ ;
wire _6776_ ;
wire _6356_ ;
wire _1491_ ;
wire _1071_ ;
wire _2696_ ;
wire _2276_ ;
wire _8922_ ;
wire _8502_ ;
wire _4842_ ;
wire _4422_ ;
wire _4002_ ;
wire _5627_ ;
wire _5207_ ;
wire _8099_ ;
wire _9040_ ;
wire _1967_ ;
wire _1547_ ;
wire [31:0] \datapath.registers.838[3]  ;
wire _1127_ ;
wire _5380_ ;
wire _878_ ;
wire _458_ ;
wire _6585_ ;
wire _6165_ ;
wire _2085_ ;
wire _8731_ ;
wire _8311_ ;
wire _4651_ ;
wire _4231_ ;
wire _5856_ ;
wire _5436_ ;
wire _5016_ ;
wire _1776_ ;
wire _1356_ ;
wire _687_ ;
wire _267_ ;
wire _3922_ ;
wire _3502_ ;
wire _6394_ ;
wire _4707_ ;
wire _7599_ ;
wire _7179_ ;
wire _8960_ ;
wire _8540_ ;
wire _8120_ ;
wire _3099_ ;
wire _4880_ ;
wire _4460_ ;
wire _4040_ ;
wire _5665_ ;
wire _5245_ ;
wire \datapath.idinstr_17_bF$buf8  ;
wire _1585_ ;
wire _1165_ ;
wire _7811_ ;
wire _496_ ;
wire _3731_ ;
wire _3311_ ;
wire \datapath.alu.b_1_bF$buf0  ;
wire _4936_ ;
wire _4516_ ;
wire _9134_ ;
wire \datapath.idinstr_21_bF$buf8  ;
wire _5894_ ;
wire _5474_ ;
wire _5054_ ;
wire _6679_ ;
wire _6259_ ;
wire _1394_ ;
wire _7620_ ;
wire _7200_ ;
wire _2599_ ;
wire _2179_ ;
wire _8825_ ;
wire _8405_ ;
wire _3960_ ;
wire _3540_ ;
wire _3120_ ;
wire _4745_ ;
wire _4325_ ;
wire _24_ ;
wire _2811_ ;
wire _5283_ ;
wire [31:0] IMEM_DATA ;
wire _6488_ ;
wire _6068_ ;
wire _8634_ ;
wire _8214_ ;
wire \datapath.idinstr_17_bF$buf11  ;
wire _4974_ ;
wire _4554_ ;
wire _4134_ ;
wire [7:0] \datapath.memoryinterface.byte_size_load.byteval  ;
wire _5759_ ;
wire _5339_ ;
wire _6700_ ;
wire _9172_ ;
wire _1679_ ;
wire _1259_ ;
wire _7905_ ;
wire _2620_ ;
wire _2200_ ;
wire _5092_ ;
wire \datapath.idinstr_15_bF$buf31  ;
wire _3825_ ;
wire _3405_ ;
wire _6297_ ;
wire _8863_ ;
wire _8443_ ;
wire _8023_ ;
wire \datapath.alu.b_4_bF$buf3  ;
wire _4783_ ;
wire _4363_ ;
wire _802_ ;
wire _5988_ ;
wire _5568_ ;
wire _5148_ ;
wire \datapath.idinstr_16_bF$buf40  ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire _7714_ ;
wire _399_ ;
wire _8919_ ;
wire _3634_ ;
wire _3214_ ;
wire _4839_ ;
wire _4419_ ;
wire _8672_ ;
wire _8252_ ;
wire _1700_ ;
wire _9037_ ;
wire _4592_ ;
wire _4172_ ;
wire _611_ ;
wire _2905_ ;
wire _5797_ ;
wire _5377_ ;
wire _1297_ ;
wire _7943_ ;
wire _7523_ ;
wire _7103_ ;
wire _8728_ ;
wire _8308_ ;
wire _3863_ ;
wire _3443_ ;
wire _3023_ ;
wire _4648_ ;
wire _4228_ ;
wire _8481_ ;
wire CLK_bF$buf70 ;
wire _8061_ ;
wire CLK_bF$buf71 ;
wire CLK_bF$buf72 ;
wire CLK_bF$buf73 ;
wire CLK_bF$buf74 ;
wire CLK_bF$buf75 ;
wire CLK_bF$buf76 ;
wire CLK_bF$buf77 ;
wire CLK_bF$buf78 ;
wire CLK_bF$buf79 ;
wire _840_ ;
wire _420_ ;
wire _2714_ ;
wire _5186_ ;
wire _3919_ ;
wire _7752_ ;
wire _7332_ ;
wire _8957_ ;
wire _8537_ ;
wire _8117_ ;
wire _3672_ ;
wire _3252_ ;
wire _4877_ ;
wire _4457_ ;
wire _4037_ ;
wire _8290_ ;
wire _6603_ ;
wire _9075_ ;
wire _7808_ ;
wire _2943_ ;
wire _2523_ ;
wire _2103_ ;
wire _3728_ ;
wire _3308_ ;
wire _7981_ ;
wire _7561_ ;
wire _7141_ ;
wire _8766_ ;
wire _8346_ ;
wire _3481_ ;
wire _3061_ ;
wire _4686_ ;
wire _4266_ ;
wire _705_ ;
wire _6832_ ;
wire _6412_ ;
wire _7617_ ;
wire _2752_ ;
wire _2332_ ;
wire _3957_ ;
wire _3537_ ;
wire _3117_ ;
wire _7790_ ;
wire _7370_ ;
wire _8995_ ;
wire _8575_ ;
wire _8155_ ;
wire _3290_ ;
wire _1603_ ;
wire _4495_ ;
wire _4075_ ;
wire \datapath.idinstr_20_bF$buf14  ;
wire _934_ ;
wire _514_ ;
wire _2808_ ;
wire _6641_ ;
wire _6221_ ;
wire _7846_ ;
wire _7426_ ;
wire _7006_ ;
wire _2981_ ;
wire _2561_ ;
wire _2141_ ;
wire _3766_ ;
wire _3346_ ;
wire \datapath.idinstr_21_bF$buf23  ;
wire _5342__bF$buf0 ;
wire _5342__bF$buf1 ;
wire _5342__bF$buf2 ;
wire _5342__bF$buf3 ;
wire _5342__bF$buf4 ;
wire _5912_ ;
wire _8384_ ;
wire _1832_ ;
wire _1412_ ;
wire _9169_ ;
wire _743_ ;
wire _323_ ;
wire _2617_ ;
wire _5089_ ;
wire _6870_ ;
wire _6450_ ;
wire _6030_ ;
wire \datapath.idinstr_15_bF$buf28  ;
wire \datapath.csr.mip  ;
wire \datapath.idinstr_22_bF$buf32  ;
wire _7655_ ;
wire _7235_ ;
wire _2790_ ;
wire _2370_ ;
wire _5689__bF$buf0 ;
wire _5689__bF$buf1 ;
wire _5689__bF$buf2 ;
wire _3995_ ;
wire _5689__bF$buf3 ;
wire _3575_ ;
wire _5689__bF$buf4 ;
wire _3155_ ;
wire _5721_ ;
wire _5301_ ;
wire _8193_ ;
wire \datapath.idinstr_16_bF$buf37  ;
wire _59_ ;
wire _6926_ ;
wire _6506_ ;
wire _1641_ ;
wire _1221_ ;
wire \datapath.idinstr_20_bF$buf52  ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _2846_ ;
wire _2426_ ;
wire _2006_ ;
wire _7884_ ;
wire _7464_ ;
wire _7044_ ;
wire [31:0] \datapath.registers.838[19]  ;
wire _8669_ ;
wire _8249_ ;
wire _3384_ ;
wire _4589_ ;
wire _4169_ ;
wire _5950_ ;
wire _5530_ ;
wire _5110_ ;
wire _608_ ;
wire _6735_ ;
wire _6315_ ;
wire _1870_ ;
wire _1450_ ;
wire _1030_ ;
wire _781_ ;
wire _361_ ;
wire _2655_ ;
wire _2235_ ;
wire _4801_ ;
wire _7693_ ;
wire _7273_ ;
wire _8898_ ;
wire _8478_ ;
wire _8058_ ;
wire _3193_ ;
wire _1926_ ;
wire _1506_ ;
wire _4398_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _6964_ ;
wire _6544_ ;
wire _6124_ ;
wire _590_ ;
wire _170_ ;
wire _7749_ ;
wire _7329_ ;
wire _2884_ ;
wire _2464_ ;
wire _2044_ ;
wire _3669_ ;
wire _3249_ ;
wire _4610_ ;
wire _7082_ ;
wire _5815_ ;
wire _8287_ ;
wire _1735_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire \datapath.alu.z  ;
wire _6773_ ;
wire _6353_ ;
wire _7978_ ;
wire _7558_ ;
wire _7138_ ;
wire _2693_ ;
wire _2273_ ;
wire _3898_ ;
wire _3478_ ;
wire _3058_ ;
wire _5624_ ;
wire _5204_ ;
wire _8096_ ;
wire _6829_ ;
wire _6409_ ;
wire _1964_ ;
wire _1544_ ;
wire _1124_ ;
wire _875_ ;
wire _455_ ;
wire _2749_ ;
wire _2329_ ;
wire _6582_ ;
wire _6162_ ;
wire _7787_ ;
wire _7367_ ;
wire _2082_ ;
wire _3287_ ;
wire _5853_ ;
wire _5433_ ;
wire _5013_ ;
wire _6638_ ;
wire _6218_ ;
wire _1773_ ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire _2978_ ;
wire _2558_ ;
wire _2138_ ;
wire _6391_ ;
wire _4704_ ;
wire _7596_ ;
wire _7176_ ;
wire _5909_ ;
wire _3096_ ;
wire _1829_ ;
wire _1409_ ;
wire _5662_ ;
wire _5242_ ;
wire \datapath.idinstr_17_bF$buf5  ;
wire _6867_ ;
wire _6447_ ;
wire _6027_ ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire \datapath.idinstr_22_bF$buf29  ;
wire _2787_ ;
wire _2367_ ;
wire _4933_ ;
wire _4513_ ;
wire _5718_ ;
wire _9131_ ;
wire _1638_ ;
wire _1218_ ;
wire \datapath.idinstr_21_bF$buf5  ;
wire _5891_ ;
wire _5471_ ;
wire _5051_ ;
wire \datapath.idinstr_20_bF$buf49  ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire _6676_ ;
wire _6256_ ;
wire _1391_ ;
wire _2596_ ;
wire _2176_ ;
wire _8822_ ;
wire _8402_ ;
wire _4742_ ;
wire _4322_ ;
wire _5947_ ;
wire _5527_ ;
wire _5107_ ;
wire _21_ ;
wire _1867_ ;
wire _1447_ ;
wire _1027_ ;
wire _5280_ ;
wire _778_ ;
wire _358_ ;
wire _6485_ ;
wire _6065_ ;
wire _8631_ ;
wire _8211_ ;
wire _4971_ ;
wire _4551_ ;
wire _4131_ ;
wire _5756_ ;
wire _5336_ ;
wire _1676_ ;
wire _1256_ ;
wire _7902_ ;
wire _587_ ;
wire _167_ ;
wire _3822_ ;
wire _3402_ ;
wire _6294_ ;
wire _4607_ ;
wire [31:0] \datapath._03_  ;
wire _7499_ ;
wire _7079_ ;
wire _8860_ ;
wire _8440_ ;
wire _8020_ ;
wire \datapath.alu.b_4_bF$buf0  ;
wire _4780_ ;
wire _4360_ ;
wire _5985_ ;
wire _5565_ ;
wire _5145_ ;
wire _1485_ ;
wire _1065_ ;
wire _7711_ ;
wire _396_ ;
wire _8916_ ;
wire _3631_ ;
wire _3211_ ;
wire _4836_ ;
wire _4416_ ;
wire _9034_ ;
wire \datapath.alu.b_2_bF$buf7  ;
wire _2902_ ;
wire _5794_ ;
wire _5374_ ;
wire _6999_ ;
wire _6579_ ;
wire _6159_ ;
wire _1294_ ;
wire _7940_ ;
wire _7520_ ;
wire _7100_ ;
wire _2499_ ;
wire _2079_ ;
wire _8725_ ;
wire _8305_ ;
wire _3860_ ;
wire _3440_ ;
wire _3020_ ;
wire _4645_ ;
wire _4225_ ;
wire CLK_bF$buf40 ;
wire CLK_bF$buf41 ;
wire CLK_bF$buf42 ;
wire _3557__bF$buf0 ;
wire CLK_bF$buf43 ;
wire _3557__bF$buf1 ;
wire CLK_bF$buf44 ;
wire _3557__bF$buf2 ;
wire CLK_bF$buf45 ;
wire _3557__bF$buf3 ;
wire CLK_bF$buf46 ;
wire _3557__bF$buf4 ;
wire CLK_bF$buf47 ;
wire CLK_bF$buf48 ;
wire CLK_bF$buf49 ;
wire _2711_ ;
wire _5183_ ;
wire _3916_ ;
wire _6388_ ;
wire _8954_ ;
wire _8534_ ;
wire _8114_ ;
wire _4874_ ;
wire _4454_ ;
wire _4034_ ;
wire _3561__bF$buf0 ;
wire _3561__bF$buf1 ;
wire _3561__bF$buf2 ;
wire _3561__bF$buf3 ;
wire _3561__bF$buf4 ;
wire _5659_ ;
wire _5239_ ;
wire _6600_ ;
wire _9072_ ;
wire _1999_ ;
wire _1579_ ;
wire _1159_ ;
wire _7805_ ;
wire _2940_ ;
wire _2520_ ;
wire _2100_ ;
wire _3725_ ;
wire _3305_ ;
wire _6197_ ;
wire _8763_ ;
wire _8343_ ;
wire _9128_ ;
wire _4683_ ;
wire _4263_ ;
wire _702_ ;
wire _5888_ ;
wire _5468_ ;
wire _5048_ ;
wire _1388_ ;
wire _7614_ ;
wire _299_ ;
wire \datapath.idinstr_20_hier0_bF$buf6  ;
wire _8819_ ;
wire _3954_ ;
wire _3534_ ;
wire _3114_ ;
wire _4739_ ;
wire _4319_ ;
wire _8992_ ;
wire _8572_ ;
wire _8152_ ;
wire _18_ ;
wire _1600_ ;
wire _4492_ ;
wire _4072_ ;
wire \datapath.idinstr_20_bF$buf11  ;
wire _931_ ;
wire _511_ ;
wire _2805_ ;
wire _5697_ ;
wire _5277_ ;
wire _1197_ ;
wire _7843_ ;
wire _7423_ ;
wire _7003_ ;
wire _8628_ ;
wire _8208_ ;
wire _3763_ ;
wire _3343_ ;
wire _4968_ ;
wire _4548_ ;
wire \datapath.idinstr_21_bF$buf20  ;
wire _4128_ ;
wire _8381_ ;
wire _9166_ ;
wire _740_ ;
wire _320_ ;
wire _2614_ ;
wire _5086_ ;
wire \datapath.idinstr_15_bF$buf25  ;
wire _3819_ ;
wire _7652_ ;
wire _7232_ ;
wire _8857_ ;
wire _8437_ ;
wire _8017_ ;
wire _3992_ ;
wire _3572_ ;
wire _3152_ ;
wire _4777_ ;
wire _4357_ ;
wire _8190_ ;
wire \datapath.idinstr_16_bF$buf34  ;
wire _56_ ;
wire _6923_ ;
wire _6503_ ;
wire _7708_ ;
wire _2843_ ;
wire _2423_ ;
wire _2003_ ;
wire _3628_ ;
wire _3208_ ;
wire _4969__bF$buf0 ;
wire _4969__bF$buf1 ;
wire _4969__bF$buf2 ;
wire _4969__bF$buf3 ;
wire _4969__bF$buf4 ;
wire _4969__bF$buf5 ;
wire _7881_ ;
wire _4969__bF$buf6 ;
wire _7461_ ;
wire _4969__bF$buf7 ;
wire _7041_ ;
wire _8666_ ;
wire _8246_ ;
wire _3381_ ;
wire _4586_ ;
wire _4166_ ;
wire _605_ ;
wire _6732_ ;
wire _6312_ ;
wire _7937_ ;
wire _7517_ ;
wire _2652_ ;
wire _2232_ ;
wire _3857_ ;
wire _3437_ ;
wire _3017_ ;
wire _7690_ ;
wire _7270_ ;
wire _8895_ ;
wire _8475_ ;
wire _8055_ ;
wire _3190_ ;
wire _1923_ ;
wire _1503_ ;
wire _4395_ ;
wire _834_ ;
wire _414_ ;
wire _2708_ ;
wire _94_ ;
wire _6961_ ;
wire _6541_ ;
wire _6121_ ;
wire _7746_ ;
wire _7326_ ;
wire _2881_ ;
wire _2461_ ;
wire _2041_ ;
wire _3666_ ;
wire _3246_ ;
wire _5812_ ;
wire _8284_ ;
wire _1732_ ;
wire _1312_ ;
wire _9069_ ;
wire _643_ ;
wire _223_ ;
wire _2937_ ;
wire _2517_ ;
wire _6770_ ;
wire _6350_ ;
wire _7975_ ;
wire _7555_ ;
wire _7135_ ;
wire _2690_ ;
wire _2270_ ;
wire _3895_ ;
wire _3475_ ;
wire _9092__bF$buf0 ;
wire _3055_ ;
wire _9092__bF$buf1 ;
wire _9092__bF$buf2 ;
wire _9092__bF$buf3 ;
wire _9092__bF$buf4 ;
wire _9092__bF$buf5 ;
wire _9092__bF$buf6 ;
wire _9092__bF$buf7 ;
wire _9092__bF$buf8 ;
wire [31:0] \datapath.memdataload  ;
wire _5621_ ;
wire _5201_ ;
wire _8093_ ;
wire _6826_ ;
wire _6406_ ;
wire _1961_ ;
wire _1541_ ;
wire _1121_ ;
wire _872_ ;
wire _452_ ;
wire _2746_ ;
wire _2326_ ;
wire _7784_ ;
wire _7364_ ;
wire _8989_ ;
wire _8569_ ;
wire _8149_ ;
wire _3284_ ;
wire _4489_ ;
wire _4069_ ;
wire _5850_ ;
wire _5430_ ;
wire _5010_ ;
wire _928_ ;
wire _508_ ;
wire _6635_ ;
wire _6215_ ;
wire _1770_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _2975_ ;
wire _2555_ ;
wire _2135_ ;
wire _4701_ ;
wire _7593_ ;
wire _7173_ ;
wire \datapath.idinstr_21_bF$buf17  ;
wire _5906_ ;
wire _2014__bF$buf0 ;
wire _2014__bF$buf1 ;
wire _2014__bF$buf2 ;
wire _2014__bF$buf3 ;
wire _8798_ ;
wire _8378_ ;
wire _3093_ ;
wire _1826_ ;
wire _1406_ ;
wire _4298_ ;
wire _737_ ;
wire _317_ ;
wire \datapath.idinstr_17_bF$buf2  ;
wire _6864_ ;
wire _6444_ ;
wire _6024_ ;
wire _490_ ;
wire \datapath.idinstr_22_bF$buf26  ;
wire _7649_ ;
wire _7229_ ;
wire _2784_ ;
wire _2364_ ;
wire _3989_ ;
wire _3569_ ;
wire _3149_ ;
wire _4930_ ;
wire _4510_ ;
wire _5715_ ;
wire _8187_ ;
wire _1635_ ;
wire _1215_ ;
wire \datapath.idinstr_21_bF$buf2  ;
wire \datapath.idinstr_20_bF$buf46  ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire \datapath.idinstr_15_bF$buf9  ;
wire _6673_ ;
wire _6253_ ;
wire _7878_ ;
wire _7458_ ;
wire _7038_ ;
wire _2593_ ;
wire _2173_ ;
wire _3798_ ;
wire _3378_ ;
wire _5408__bF$buf0 ;
wire _5408__bF$buf1 ;
wire _5408__bF$buf2 ;
wire _5408__bF$buf3 ;
wire _5408__bF$buf4 ;
wire _5408__bF$buf5 ;
wire _5408__bF$buf6 ;
wire _5408__bF$buf7 ;
wire _5944_ ;
wire _5524_ ;
wire _5104_ ;
wire _6729_ ;
wire _6309_ ;
wire _1864_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire [31:0] \datapath.registers.regb_data  ;
wire _2649_ ;
wire _2229_ ;
wire _6482_ ;
wire _6062_ ;
wire _7687_ ;
wire _7267_ ;
wire _3187_ ;
wire _5753_ ;
wire _5333_ ;
wire _4819__bF$buf0 ;
wire _4819__bF$buf1 ;
wire _4819__bF$buf2 ;
wire _4819__bF$buf3 ;
wire _6958_ ;
wire _4819__bF$buf4 ;
wire _6538_ ;
wire _6118_ ;
wire _1673_ ;
wire _1253_ ;
wire _584_ ;
wire _164_ ;
wire _2878_ ;
wire _2458_ ;
wire _2038_ ;
wire _6291_ ;
wire _4604_ ;
wire _7496_ ;
wire _7076_ ;
wire _5759__bF$buf0 ;
wire _5759__bF$buf1 ;
wire _5759__bF$buf2 ;
wire _5759__bF$buf3 ;
wire _5759__bF$buf4 ;
wire _5809_ ;
wire _1729_ ;
wire _1309_ ;
wire _5982_ ;
wire _5562_ ;
wire _5142_ ;
wire _4823__bF$buf0 ;
wire _4823__bF$buf1 ;
wire _4823__bF$buf2 ;
wire _4823__bF$buf3 ;
wire _4823__bF$buf4 ;
wire _6767_ ;
wire _6347_ ;
wire _1482_ ;
wire _1062_ ;
wire _393_ ;
wire \datapath.idinstr_24_bF$buf5  ;
wire _2687_ ;
wire _2267_ ;
wire _8913_ ;
wire _4833_ ;
wire _4413_ ;
wire _5618_ ;
wire _9031_ ;
wire \datapath.alu.b_2_bF$buf4  ;
wire _1958_ ;
wire _1538_ ;
wire _1118_ ;
wire _5791_ ;
wire _5371_ ;
wire _869_ ;
wire _449_ ;
wire _6996_ ;
wire _6576_ ;
wire _6156_ ;
wire _1291_ ;
wire _2496_ ;
wire _2076_ ;
wire _8722_ ;
wire _8302_ ;
wire _4642_ ;
wire _4222_ ;
wire CLK_bF$buf10 ;
wire CLK_bF$buf11 ;
wire CLK_bF$buf12 ;
wire CLK_bF$buf13 ;
wire CLK_bF$buf14 ;
wire CLK_bF$buf15 ;
wire CLK_bF$buf16 ;
wire CLK_bF$buf17 ;
wire CLK_bF$buf18 ;
wire CLK_bF$buf19 ;
wire _5847_ ;
wire _5427_ ;
wire _5007_ ;
wire _1767_ ;
wire _1347_ ;
wire _5180_ ;
wire _678_ ;
wire _258_ ;
wire _3913_ ;
wire _6385_ ;
wire _2597__bF$buf0 ;
wire _2597__bF$buf1 ;
wire _2597__bF$buf2 ;
wire _2597__bF$buf3 ;
wire _2597__bF$buf4 ;
wire _2597__bF$buf5 ;
wire _8951_ ;
wire _8531_ ;
wire _8111_ ;
wire _4871_ ;
wire _4451_ ;
wire _4031_ ;
wire _5656_ ;
wire _5236_ ;
wire _1996_ ;
wire _1576_ ;
wire _1156_ ;
wire _7802_ ;
wire _487_ ;
wire [31:0] DMEM_DATA_L ;
wire _3722_ ;
wire _3302_ ;
wire [31:0] DMEM_DATA_S ;
wire _6194_ ;
wire _4927_ ;
wire _4507_ ;
wire _7399_ ;
wire _8760_ ;
wire _8340_ ;
wire _9125_ ;
wire _4680_ ;
wire _4260_ ;
wire _5885_ ;
wire _5465_ ;
wire _5045_ ;
wire _1385_ ;
wire _7611_ ;
wire _296_ ;
wire \datapath.idinstr_20_hier0_bF$buf3  ;
wire _8816_ ;
wire _3951_ ;
wire _3531_ ;
wire _3111_ ;
wire _4736_ ;
wire _4316_ ;
wire _15_ ;
wire _2802_ ;
wire _5694_ ;
wire _5274_ ;
wire _6899_ ;
wire _6479_ ;
wire _6059_ ;
wire _1194_ ;
wire _7840_ ;
wire _7420_ ;
wire _7000_ ;
wire _2399_ ;
wire _8625_ ;
wire _8205_ ;
wire _3760_ ;
wire _3340_ ;
wire _4965_ ;
wire _4545_ ;
wire _4125_ ;
wire _9163_ ;
wire _2611_ ;
wire _5083_ ;
wire \datapath.idinstr_15_bF$buf22  ;
wire _3816_ ;
wire _6288_ ;
wire _8854_ ;
wire _8434_ ;
wire _8014_ ;
wire _4774_ ;
wire _4354_ ;
wire _5979_ ;
wire _5559_ ;
wire _5139_ ;
wire \datapath.idinstr_16_bF$buf31  ;
wire _53_ ;
wire _6920_ ;
wire _6500_ ;
wire _1899_ ;
wire _1479_ ;
wire _1059_ ;
wire _7705_ ;
wire _2840_ ;
wire _2420_ ;
wire _2000_ ;
wire _3625_ ;
wire _3205_ ;
wire _6097_ ;
wire _8663_ ;
wire _8243_ ;
wire _9028_ ;
wire _4583_ ;
wire _4163_ ;
wire _602_ ;
wire _5788_ ;
wire _5368_ ;
wire _1288_ ;
wire _7934_ ;
wire _7514_ ;
wire _199_ ;
wire [31:0] \datapath.registers.838[24]  ;
wire _8719_ ;
wire _3854_ ;
wire _3434_ ;
wire _3014_ ;
wire _4639_ ;
wire _4219_ ;
wire _8892_ ;
wire _8472_ ;
wire _8052_ ;
wire _1920_ ;
wire _1500_ ;
wire _4392_ ;
wire _831_ ;
wire _411_ ;
wire _2705_ ;
wire _5597_ ;
wire _5177_ ;
wire _91_ ;
wire _1097_ ;
wire _7743_ ;
wire _7323_ ;
wire _8948_ ;
wire _8528_ ;
wire _8108_ ;
wire _3663_ ;
wire _3243_ ;
wire _4868_ ;
wire _4448_ ;
wire _4028_ ;
wire _8281_ ;
wire _9066_ ;
wire _640_ ;
wire _220_ ;
wire _2934_ ;
wire _2514_ ;
wire _3719_ ;
wire _7972_ ;
wire _7552_ ;
wire _7132_ ;
wire _8757_ ;
wire _8337_ ;
wire _3892_ ;
wire _3472_ ;
wire _3052_ ;
wire _4677_ ;
wire _4257_ ;
wire _8090_ ;
wire _3134__bF$buf0 ;
wire _3134__bF$buf1 ;
wire _3134__bF$buf2 ;
wire _3134__bF$buf3 ;
wire _6823_ ;
wire _3134__bF$buf4 ;
wire _6403_ ;
wire _3134__bF$buf5 ;
wire CLK_hier0_bF$buf10 ;
wire CLK_hier0_bF$buf11 ;
wire _7608_ ;
wire _2743_ ;
wire _2323_ ;
wire _3948_ ;
wire _3528_ ;
wire _3108_ ;
wire _9_ ;
wire _7781_ ;
wire _7361_ ;
wire _8986_ ;
wire _8566_ ;
wire _8146_ ;
wire _3281_ ;
wire _4486_ ;
wire _4066_ ;
wire _925_ ;
wire _505_ ;
wire _6632_ ;
wire _6212_ ;
wire _7837_ ;
wire _7417_ ;
wire _2972_ ;
wire _2552_ ;
wire _2132_ ;
wire _3757_ ;
wire _3337_ ;
wire _7590_ ;
wire _7170_ ;
wire \datapath.idinstr_21_bF$buf14  ;
wire _5903_ ;
wire _8795_ ;
wire _8375_ ;
wire _3090_ ;
wire _1823_ ;
wire _1403_ ;
wire _4295_ ;
wire _734_ ;
wire _314_ ;
wire _2608_ ;
wire _6861_ ;
wire _6441_ ;
wire _6021_ ;
wire \datapath.idinstr_15_bF$buf19  ;
wire \datapath.idinstr_22_bF$buf23  ;
wire _7646_ ;
wire _7226_ ;
wire _2781_ ;
wire _2361_ ;
wire _3986_ ;
wire _3566_ ;
wire _3146_ ;
wire _5712_ ;
wire _8184_ ;
wire \datapath.idinstr_16_bF$buf28  ;
wire _6917_ ;
wire _1632_ ;
wire _1212_ ;
wire \datapath.idinstr_20_bF$buf43  ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _2837_ ;
wire \datapath.idinstr_15_bF$buf6  ;
wire _2417_ ;
wire _6670_ ;
wire _6250_ ;
wire _7875_ ;
wire _7455_ ;
wire _7035_ ;
wire _2590_ ;
wire _2170_ ;
wire _3795_ ;
wire _3375_ ;
wire _5941_ ;
wire _5521_ ;
wire _5101_ ;
wire _6726_ ;
wire _6306_ ;
wire _1861_ ;
wire _1441_ ;
wire _1021_ ;
wire _772_ ;
wire _352_ ;
wire _2646_ ;
wire _2226_ ;
wire _7684_ ;
wire _7264_ ;
wire _8889_ ;
wire _8469_ ;
wire _8049_ ;
wire _3184_ ;
wire _1917_ ;
wire _4389_ ;
wire _5750_ ;
wire _5330_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _6955_ ;
wire _6535_ ;
wire _6115_ ;
wire _1670_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _2875_ ;
wire _2455_ ;
wire _2035_ ;
wire _4601_ ;
wire _7493_ ;
wire _7073_ ;
wire _5806_ ;
wire _8698_ ;
wire _8278_ ;
wire _1726_ ;
wire _1306_ ;
wire _4198_ ;
wire _637_ ;
wire _217_ ;
wire _6764_ ;
wire _6344_ ;
wire _390_ ;
wire _7969_ ;
wire _7549_ ;
wire _7129_ ;
wire \datapath.idinstr_24_bF$buf2  ;
wire _2684_ ;
wire _2264_ ;
wire _8910_ ;
wire _3889_ ;
wire _3469_ ;
wire _3049_ ;
wire _4830_ ;
wire _4410_ ;
wire _5615_ ;
wire _8087_ ;
wire \datapath.alu.b_2_bF$buf1  ;
wire _1955_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire \datapath.tkbranch  ;
wire _6993_ ;
wire _6573_ ;
wire _6153_ ;
wire _2781__bF$buf0 ;
wire _2781__bF$buf1 ;
wire _2781__bF$buf2 ;
wire _2781__bF$buf3 ;
wire _2781__bF$buf4 ;
wire \controlunit.csrfile_trap_wen_bF$buf7  ;
wire _7778_ ;
wire _7358_ ;
wire _2493_ ;
wire _2073_ ;
wire \datapath.idinstr_22_bF$buf9  ;
wire _3698_ ;
wire _3278_ ;
wire _5844_ ;
wire _5424_ ;
wire _5004_ ;
wire _6629_ ;
wire _6209_ ;
wire _1764_ ;
wire _1344_ ;
wire _675_ ;
wire _255_ ;
wire _2969_ ;
wire _2549_ ;
wire _2129_ ;
wire _3910_ ;
wire _6382_ ;
wire _7587_ ;
wire _7167_ ;
wire _9158__bF$buf0 ;
wire _9158__bF$buf1 ;
wire _9158__bF$buf2 ;
wire _9158__bF$buf3 ;
wire _9158__bF$buf4 ;
wire _3087_ ;
wire _5653_ ;
wire _5233_ ;
wire _6858_ ;
wire _6438_ ;
wire _6018_ ;
wire _1993_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _2778_ ;
wire _2358_ ;
wire _6191_ ;
wire _4924_ ;
wire _4504_ ;
wire _7396_ ;
wire _5709_ ;
wire _9122_ ;
wire _1629_ ;
wire _1209_ ;
wire _5882_ ;
wire _5462_ ;
wire _5042_ ;
wire _6667_ ;
wire _6247_ ;
wire _1382_ ;
wire _293_ ;
wire _2587_ ;
wire _2167_ ;
wire \datapath.idinstr_20_hier0_bF$buf0  ;
wire _8813_ ;
wire _4733_ ;
wire _4313_ ;
wire \datapath.idinstr_21_bF$buf49  ;
wire _5938_ ;
wire _5518_ ;
wire _12_ ;
wire _1858_ ;
wire _1438_ ;
wire _1018_ ;
wire _5691_ ;
wire _5271_ ;
wire _769_ ;
wire _349_ ;
wire _6896_ ;
wire _6476_ ;
wire _6056_ ;
wire _1191_ ;
wire _2396_ ;
wire _8622_ ;
wire _8202_ ;
wire _4962_ ;
wire _4542_ ;
wire _4122_ ;
wire _5747_ ;
wire _5327_ ;
wire _9160_ ;
wire _1667_ ;
wire _1247_ ;
wire _5080_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _3813_ ;
wire _6285_ ;
wire _8851_ ;
wire _8431_ ;
wire _8011_ ;
wire _4771_ ;
wire _4351_ ;
wire \datapath.idinstr_21_hier0_bF$buf5  ;
wire _5976_ ;
wire _5556_ ;
wire _5136_ ;
wire _50_ ;
wire _1896_ ;
wire _1476_ ;
wire _1056_ ;
wire _7702_ ;
wire _387_ ;
wire _8907_ ;
wire _3622_ ;
wire _7420__bF$buf0 ;
wire _3202_ ;
wire _7420__bF$buf1 ;
wire _7420__bF$buf2 ;
wire _7420__bF$buf3 ;
wire _7420__bF$buf4 ;
wire _7420__bF$buf5 ;
wire _7420__bF$buf6 ;
wire _7420__bF$buf7 ;
wire _7420__bF$buf8 ;
wire _6094_ ;
wire _7420__bF$buf9 ;
wire _4827_ ;
wire _4407_ ;
wire _7299_ ;
wire _8660_ ;
wire _8240_ ;
wire _9025_ ;
wire _4580_ ;
wire _4160_ ;
wire _5785_ ;
wire _5365_ ;
wire _1285_ ;
wire _7931_ ;
wire _7511_ ;
wire _196_ ;
wire _8716_ ;
wire _3851_ ;
wire _3431_ ;
wire _3011_ ;
wire _4636_ ;
wire _4216_ ;
wire _2702_ ;
wire _5594_ ;
wire _5174_ ;
wire _3907_ ;
wire _6799_ ;
wire _6379_ ;
wire _1094_ ;
wire _7740_ ;
wire _7320_ ;
wire _2299_ ;
wire _8945_ ;
wire _8525_ ;
wire _8105_ ;
wire _3660_ ;
wire _3240_ ;
wire _4865_ ;
wire _4445_ ;
wire _4025_ ;
wire _9063_ ;
wire _2931_ ;
wire _2511_ ;
wire _3716_ ;
wire _6188_ ;
wire _8754_ ;
wire _8334_ ;
wire _9119_ ;
wire _4674_ ;
wire _4254_ ;
wire _5879_ ;
wire _5459_ ;
wire _5039_ ;
wire _6820_ ;
wire _6400_ ;
wire _1799_ ;
wire _1379_ ;
wire _7605_ ;
wire _2740_ ;
wire _2320_ ;
wire _3945_ ;
wire _3525_ ;
wire _3105_ ;
wire _6_ ;
wire _8983_ ;
wire _8563_ ;
wire _8143_ ;
wire _4483_ ;
wire _4063_ ;
wire _922_ ;
wire _502_ ;
wire _5688_ ;
wire _5268_ ;
wire _1188_ ;
wire _7834_ ;
wire _7414_ ;
wire [31:0] \datapath.registers.838[14]  ;
wire _8619_ ;
wire _3754_ ;
wire _3334_ ;
wire _4959_ ;
wire _4539_ ;
wire \datapath.idinstr_21_bF$buf11  ;
wire _4119_ ;
wire _5900_ ;
wire _8792_ ;
wire _8372_ ;
wire _1820_ ;
wire _1400_ ;
wire _9157_ ;
wire _4292_ ;
wire _731_ ;
wire _311_ ;
wire _2605_ ;
wire _5497_ ;
wire _5077_ ;
wire \datapath.idinstr_15_bF$buf16  ;
wire \datapath.idinstr_15_hier0_bF$buf4  ;
wire \datapath.idinstr_22_bF$buf20  ;
wire _7643_ ;
wire _7223_ ;
wire _8848_ ;
wire _8428_ ;
wire _8008_ ;
wire _3983_ ;
wire _3563_ ;
wire _3143_ ;
wire _4768_ ;
wire _4348_ ;
wire _8181_ ;
wire \datapath.idinstr_16_bF$buf25  ;
wire _47_ ;
wire _6914_ ;
wire \datapath.idinstr_20_bF$buf40  ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _2834_ ;
wire \datapath.idinstr_15_bF$buf3  ;
wire _2414_ ;
wire _3619_ ;
wire _7872_ ;
wire _7452_ ;
wire _7032_ ;
wire _8657_ ;
wire _8237_ ;
wire _3792_ ;
wire _3372_ ;
wire _4997_ ;
wire _4577_ ;
wire _4157_ ;
wire _6723_ ;
wire _6303_ ;
wire _7928_ ;
wire _7508_ ;
wire _2643_ ;
wire _2223_ ;
wire \datapath.idinstr_15_bF$buf54  ;
wire _3848_ ;
wire _3428_ ;
wire _3008_ ;
wire _7681_ ;
wire _7261_ ;
wire _8886_ ;
wire _8466_ ;
wire _8046_ ;
wire _3181_ ;
wire _1914_ ;
wire _4386_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _6952_ ;
wire _6532_ ;
wire _6112_ ;
wire _7737_ ;
wire _7317_ ;
wire _2872_ ;
wire _2452_ ;
wire _2032_ ;
wire _3657_ ;
wire _3237_ ;
wire _7490_ ;
wire _7070_ ;
wire _5803_ ;
wire _8695_ ;
wire _8275_ ;
wire _1723_ ;
wire _1303_ ;
wire _4195_ ;
wire _634_ ;
wire _214_ ;
wire _2928_ ;
wire _2508_ ;
wire _6761_ ;
wire _6341_ ;
wire _7966_ ;
wire _7546_ ;
wire _7126_ ;
wire _2681_ ;
wire _2261_ ;
wire \datapath.idinstr_18_bF$buf6  ;
wire _3886_ ;
wire _3466_ ;
wire _3046_ ;
wire _5612_ ;
wire _8084_ ;
wire _6817_ ;
wire _1952_ ;
wire _1532_ ;
wire _1112_ ;
wire _863_ ;
wire _443_ ;
wire _2737_ ;
wire _2317_ ;
wire _6990_ ;
wire _6570_ ;
wire _6150_ ;
wire \controlunit.csrfile_trap_wen_bF$buf4  ;
wire _7775_ ;
wire _7355_ ;
wire _2490_ ;
wire _2070_ ;
wire \datapath.idinstr_22_bF$buf6  ;
wire _3695_ ;
wire _3275_ ;
wire _5841_ ;
wire _5421_ ;
wire _5001_ ;
wire _919_ ;
wire _6626_ ;
wire _6206_ ;
wire _1761_ ;
wire _1341_ ;
wire _9098_ ;
wire _672_ ;
wire _252_ ;
wire _2966_ ;
wire _2546_ ;
wire _2126_ ;
wire _7584_ ;
wire _7164_ ;
wire _8789_ ;
wire _8369_ ;
wire _3084_ ;
wire _1817_ ;
wire _4289_ ;
wire _5650_ ;
wire _5230_ ;
wire _728_ ;
wire _308_ ;
wire [1:0] \controlunit.pc_sel  ;
wire _6855_ ;
wire _6435_ ;
wire _6015_ ;
wire _1990_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire \datapath.idinstr_22_bF$buf17  ;
wire _2775_ ;
wire _2355_ ;
wire _2118__bF$buf0 ;
wire _2118__bF$buf1 ;
wire _2118__bF$buf2 ;
wire _2118__bF$buf3 ;
wire _4921_ ;
wire _4501_ ;
wire _7393_ ;
wire _5706_ ;
wire _8598_ ;
wire _8178_ ;
wire _1626_ ;
wire _1206_ ;
wire _4098_ ;
wire \datapath.idinstr_20_bF$buf37  ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire _6664_ ;
wire _6244_ ;
wire _290_ ;
wire _7869_ ;
wire _7449_ ;
wire _7029_ ;
wire _2584_ ;
wire _2164_ ;
wire _8810_ ;
wire _3789_ ;
wire _3369_ ;
wire _4730_ ;
wire _4310_ ;
wire \datapath.idinstr_21_bF$buf46  ;
wire _5935_ ;
wire _5515_ ;
wire \datapath.alu.b_0_bF$buf7  ;
wire _1855_ ;
wire _1435_ ;
wire _1015_ ;
wire _766_ ;
wire _346_ ;
wire _6893_ ;
wire _6473_ ;
wire _6053_ ;
wire _7678_ ;
wire _7258_ ;
wire _2393_ ;
wire _3598_ ;
wire _3178_ ;
wire _5744_ ;
wire _5324_ ;
wire [29:0] \datapath.csr._26_  ;
wire _6949_ ;
wire _6529_ ;
wire _6109_ ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire _2869_ ;
wire _2449_ ;
wire _2029_ ;
wire _3810_ ;
wire _6282_ ;
wire _7487_ ;
wire _7067_ ;
wire _4829__bF$buf0 ;
wire _4829__bF$buf1 ;
wire _4829__bF$buf2 ;
wire _4829__bF$buf3 ;
wire _4829__bF$buf4 ;
wire \datapath.idinstr_21_hier0_bF$buf2  ;
wire _5973_ ;
wire _5553_ ;
wire _5133_ ;
wire _6758_ ;
wire _6338_ ;
wire _1893_ ;
wire _1473_ ;
wire _1053_ ;
wire _384_ ;
wire _2678_ ;
wire _2258_ ;
wire _8904_ ;
wire _6091_ ;
wire _4824_ ;
wire _4404_ ;
wire _7296_ ;
wire _5609_ ;
wire _4833__bF$buf0 ;
wire _4833__bF$buf1 ;
wire _4833__bF$buf2 ;
wire _4833__bF$buf3 ;
wire _4833__bF$buf4 ;
wire _9022_ ;
wire _1949_ ;
wire _1529_ ;
wire _1109_ ;
wire _5782_ ;
wire _5362_ ;
wire [1:0] \controlunit.wb_sel  ;
wire _6987_ ;
wire _6567_ ;
wire _6147_ ;
wire _1282_ ;
wire _193_ ;
wire _2487_ ;
wire _2067_ ;
wire _8713_ ;
wire _4633_ ;
wire _4213_ ;
wire _5838_ ;
wire _5418_ ;
wire _1758_ ;
wire _1338_ ;
wire _5591_ ;
wire _5171_ ;
wire _669_ ;
wire _249_ ;
wire _3904_ ;
wire _6796_ ;
wire _6376_ ;
wire _1091_ ;
wire _2296_ ;
wire _8942_ ;
wire _8522_ ;
wire _8102_ ;
wire [31:0] \datapath.alupc  ;
wire _7419__bF$buf0 ;
wire _7419__bF$buf1 ;
wire _4862_ ;
wire _7419__bF$buf2 ;
wire _4442_ ;
wire _7419__bF$buf3 ;
wire _4022_ ;
wire _7419__bF$buf4 ;
wire _7419__bF$buf5 ;
wire _7419__bF$buf6 ;
wire _7419__bF$buf7 ;
wire _7419__bF$buf8 ;
wire _7419__bF$buf9 ;
wire _5647_ ;
wire _5227_ ;
wire _9060_ ;
wire _1987_ ;
wire _1567_ ;
wire [31:0] \datapath.registers.838[5]  ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _3713_ ;
wire _6185_ ;
wire _4918_ ;
wire _8751_ ;
wire _8331_ ;
wire _7423__bF$buf0 ;
wire _7423__bF$buf1 ;
wire _7423__bF$buf2 ;
wire _7423__bF$buf3 ;
wire _7423__bF$buf4 ;
wire _7423__bF$buf5 ;
wire _7423__bF$buf6 ;
wire _7423__bF$buf7 ;
wire _9116_ ;
wire _4671_ ;
wire _4251_ ;
wire _5876_ ;
wire _5456_ ;
wire _5036_ ;
wire _1796_ ;
wire _1376_ ;
wire _7602_ ;
wire _287_ ;
wire _8807_ ;
wire _3942_ ;
wire _3522_ ;
wire _3102_ ;
wire [3:0] _3_ ;
wire _4727_ ;
wire _4307_ ;
wire _7199_ ;
wire _8980_ ;
wire _8560_ ;
wire _8140_ ;
wire _4480_ ;
wire _4060_ ;
wire _5685_ ;
wire _5265_ ;
wire _1185_ ;
wire _7831_ ;
wire _7411_ ;
wire _8616_ ;
wire _3751_ ;
wire _3331_ ;
wire _4956_ ;
wire _4536_ ;
wire _4116_ ;
wire _9154_ ;
wire _2602_ ;
wire _5494_ ;
wire _5074_ ;
wire CLK_bF$buf130 ;
wire CLK_bF$buf131 ;
wire CLK_bF$buf132 ;
wire CLK_bF$buf133 ;
wire CLK_bF$buf134 ;
wire CLK_bF$buf135 ;
wire \datapath.idinstr_15_bF$buf13  ;
wire CLK_bF$buf136 ;
wire CLK_bF$buf137 ;
wire CLK_bF$buf138 ;
wire _3807_ ;
wire CLK_bF$buf139 ;
wire \datapath.idinstr_15_hier0_bF$buf1  ;
wire _6699_ ;
wire _6279_ ;
wire _7640_ ;
wire _7220_ ;
wire _2199_ ;
wire _8845_ ;
wire _8425_ ;
wire _8005_ ;
wire _3980_ ;
wire _3560_ ;
wire _3140_ ;
wire _4765_ ;
wire _4345_ ;
wire \datapath.idinstr_16_bF$buf22  ;
wire _44_ ;
wire _6911_ ;
wire _2831_ ;
wire \datapath.idinstr_15_bF$buf0  ;
wire _2411_ ;
wire _3616_ ;
wire _6088_ ;
wire _4900__bF$buf0 ;
wire _4900__bF$buf1 ;
wire _4900__bF$buf2 ;
wire _4900__bF$buf3 ;
wire _4900__bF$buf4 ;
wire _8654_ ;
wire _8234_ ;
wire _9019_ ;
wire _4994_ ;
wire _4574_ ;
wire _4154_ ;
wire _5779_ ;
wire _5359_ ;
wire _6720_ ;
wire _6300_ ;
wire _1699_ ;
wire _1279_ ;
wire _7925_ ;
wire _7505_ ;
wire _2640_ ;
wire _2220_ ;
wire \datapath.idinstr_15_bF$buf51  ;
wire _3845_ ;
wire _3425_ ;
wire _3005_ ;
wire _8883_ ;
wire _8463_ ;
wire _8043_ ;
wire \datapath.idinstr_16_hier0_bF$buf6  ;
wire _1911_ ;
wire _4383_ ;
wire _822_ ;
wire _402_ ;
wire _5588_ ;
wire _5168_ ;
wire _82_ ;
wire _1088_ ;
wire _7734_ ;
wire _7314_ ;
wire _8939_ ;
wire _8519_ ;
wire _3654_ ;
wire _3234_ ;
wire _4859_ ;
wire _4439_ ;
wire _4019_ ;
wire _5800_ ;
wire _8692_ ;
wire _8272_ ;
wire _1720_ ;
wire _1300_ ;
wire _9057_ ;
wire _4192_ ;
wire _631_ ;
wire _211_ ;
wire _2925_ ;
wire _2505_ ;
wire _5397_ ;
wire _7963_ ;
wire _7543_ ;
wire _7123_ ;
wire \datapath.idinstr_18_bF$buf3  ;
wire _8748_ ;
wire _8328_ ;
wire _3883_ ;
wire _3463_ ;
wire _3043_ ;
wire _0__1_bF$buf0 ;
wire _0__1_bF$buf1 ;
wire _0__1_bF$buf2 ;
wire _0__1_bF$buf3 ;
wire _0__1_bF$buf4 ;
wire _0__1_bF$buf5 ;
wire _0__1_bF$buf6 ;
wire _0__1_bF$buf7 ;
wire _4668_ ;
wire _0__1_bF$buf8 ;
wire _4248_ ;
wire _0__1_bF$buf9 ;
wire _8081_ ;
wire _189__bF$buf0 ;
wire _189__bF$buf1 ;
wire _189__bF$buf2 ;
wire _189__bF$buf3 ;
wire _189__bF$buf4 ;
wire _6814_ ;
wire _860_ ;
wire _440_ ;
wire _2734_ ;
wire _2314_ ;
wire _3939_ ;
wire _3519_ ;
wire \controlunit.csrfile_trap_wen_bF$buf1  ;
wire _7772_ ;
wire _7352_ ;
wire \datapath.idinstr_22_bF$buf3  ;
wire _8977_ ;
wire _8557_ ;
wire _8137_ ;
wire _3692_ ;
wire _3272_ ;
wire _4897_ ;
wire _4477_ ;
wire _4057_ ;
wire _916_ ;
wire _6623_ ;
wire _6203_ ;
wire _287__bF$buf0 ;
wire _287__bF$buf1 ;
wire _287__bF$buf2 ;
wire _287__bF$buf3 ;
wire _9095_ ;
wire _287__bF$buf4 ;
wire _7828_ ;
wire _7408_ ;
wire _2963_ ;
wire _2543_ ;
wire _2123_ ;
wire _3748_ ;
wire _3328_ ;
wire _7581_ ;
wire _7161_ ;
wire _8786_ ;
wire _8366_ ;
wire _3081_ ;
wire _1814_ ;
wire _4286_ ;
wire _725_ ;
wire _305_ ;
wire _6852_ ;
wire _6432_ ;
wire _6012_ ;
wire \datapath.idinstr_22_bF$buf14  ;
wire _7637_ ;
wire _7217_ ;
wire _2772_ ;
wire _2352_ ;
wire _3977_ ;
wire _3557_ ;
wire _3137_ ;
wire _7390_ ;
wire _5703_ ;
wire _8595_ ;
wire _8175_ ;
wire \datapath.idinstr_16_bF$buf19  ;
wire _6908_ ;
wire _1623_ ;
wire _1203_ ;
wire _4095_ ;
wire \datapath.idinstr_20_bF$buf34  ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _2828_ ;
wire _2408_ ;
wire _6661_ ;
wire _6241_ ;
wire _7866_ ;
wire _7446_ ;
wire _7026_ ;
wire _2581_ ;
wire _2161_ ;
wire _3786_ ;
wire _3366_ ;
wire \datapath.idinstr_21_bF$buf43  ;
wire _5932_ ;
wire _5512_ ;
wire _6717_ ;
wire \datapath.alu.b_0_bF$buf4  ;
wire _1852_ ;
wire _1432_ ;
wire _1012_ ;
wire _9189_ ;
wire _763_ ;
wire _343_ ;
wire _2637_ ;
wire _2217_ ;
wire _6890_ ;
wire _6470_ ;
wire _6050_ ;
wire \datapath.idinstr_15_bF$buf48  ;
wire _7675_ ;
wire _7255_ ;
wire _2390_ ;
wire _3595_ ;
wire _3175_ ;
wire _1908_ ;
wire _5741_ ;
wire _5321_ ;
wire _819_ ;
wire _79_ ;
wire _6946_ ;
wire _6526_ ;
wire _6106_ ;
wire _1661_ ;
wire _1241_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _2866_ ;
wire _2446_ ;
wire _2026_ ;
wire _7484_ ;
wire _7064_ ;
wire _2027__bF$buf0 ;
wire _2027__bF$buf1 ;
wire _2027__bF$buf2 ;
wire _2027__bF$buf3 ;
wire _8689_ ;
wire _8269_ ;
wire _1717_ ;
wire _4189_ ;
wire _5970_ ;
wire _5550_ ;
wire _5130_ ;
wire _628_ ;
wire _208_ ;
wire _6755_ ;
wire _6335_ ;
wire _1890_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _2675_ ;
wire _2255_ ;
wire _8901_ ;
wire _4821_ ;
wire _4401_ ;
wire _7293_ ;
wire _5606_ ;
wire _8498_ ;
wire _8078_ ;
wire _1946_ ;
wire _1526_ ;
wire _1106_ ;
wire _857_ ;
wire _437_ ;
wire _6984_ ;
wire _6564_ ;
wire _6144_ ;
wire \datapath.alu.b_3_bF$buf7  ;
wire _190_ ;
wire _7769_ ;
wire _7349_ ;
wire _2484_ ;
wire _2064_ ;
wire _8710_ ;
wire _3689_ ;
wire _3269_ ;
wire _4630_ ;
wire _4210_ ;
wire _5835_ ;
wire _5415_ ;
wire _1755_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire _3901_ ;
wire _6793_ ;
wire _6373_ ;
wire _7998_ ;
wire _7578_ ;
wire _7158_ ;
wire _2293_ ;
wire _3498_ ;
wire _3078_ ;
wire _5644_ ;
wire _5224_ ;
wire _6849_ ;
wire _6429_ ;
wire _6009_ ;
wire _1984_ ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _2769_ ;
wire _2349_ ;
wire _3710_ ;
wire _6182_ ;
wire _4915_ ;
wire _7387_ ;
wire [31:0] \datapath.jumptarget  ;
wire _9113_ ;
wire _5873_ ;
wire _5453_ ;
wire _5033_ ;
wire _6658_ ;
wire _6238_ ;
wire _1793_ ;
wire _1373_ ;
wire _284_ ;
wire _2998_ ;
wire _2578_ ;
wire _2158_ ;
wire _8804_ ;
wire [31:0] _0_ ;
wire _4724_ ;
wire _4304_ ;
wire _7196_ ;
wire _5929_ ;
wire _5509_ ;
wire _1849_ ;
wire _1429_ ;
wire _1009_ ;
wire _5682_ ;
wire _5262_ ;
wire _6887_ ;
wire _6467_ ;
wire _6047_ ;
wire _1182_ ;
wire _2387_ ;
wire _8613_ ;
wire _4953_ ;
wire _4533_ ;
wire _4113_ ;
wire _5738_ ;
wire _5318_ ;
wire _9151_ ;
wire _1658_ ;
wire _1238_ ;
wire _5491_ ;
wire _5071_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire CLK_bF$buf100 ;
wire CLK_bF$buf101 ;
wire CLK_bF$buf102 ;
wire CLK_bF$buf103 ;
wire CLK_bF$buf104 ;
wire CLK_bF$buf105 ;
wire \datapath.idinstr_15_bF$buf10  ;
wire CLK_bF$buf106 ;
wire CLK_bF$buf107 ;
wire CLK_bF$buf108 ;
wire _3804_ ;
wire CLK_bF$buf109 ;
wire _6696_ ;
wire _6276_ ;
wire _2196_ ;
wire _8842_ ;
wire _8422_ ;
wire _8002_ ;
wire _4762_ ;
wire _4342_ ;
wire _5967_ ;
wire _5547_ ;
wire _5127_ ;
wire _41_ ;
wire _1887_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _3613_ ;
wire _6085_ ;
wire _4818_ ;
wire _8651_ ;
wire _8231_ ;
wire _9016_ ;
wire _4991_ ;
wire _4571_ ;
wire _4151_ ;
wire _5776_ ;
wire _5356_ ;
wire _1696_ ;
wire _1276_ ;
wire _7922_ ;
wire _7502_ ;
wire _187_ ;
wire _8707_ ;
wire _3842_ ;
wire _3422_ ;
wire _3002_ ;
wire _4627_ ;
wire _4207_ ;
wire [31:0] \datapath._05_  ;
wire _7099_ ;
wire _8880_ ;
wire _8460_ ;
wire _8040_ ;
wire \datapath.idinstr_16_hier0_bF$buf3  ;
wire [31:0] \datapath.csr.csr_pcaddr  ;
wire _4380_ ;
wire _5585_ ;
wire _5165_ ;
wire _1085_ ;
wire _7731_ ;
wire _7311_ ;
wire _8936_ ;
wire _8516_ ;
wire _3651_ ;
wire _3231_ ;
wire _4856_ ;
wire _4436_ ;
wire _4016_ ;
wire _9054_ ;
wire _2922_ ;
wire _2502_ ;
wire _5394_ ;
wire _3707_ ;
wire _6599_ ;
wire _6179_ ;
wire _7960_ ;
wire _7540_ ;
wire _7120_ ;
wire \datapath.idinstr_18_bF$buf0  ;
wire _2099_ ;
wire _8745_ ;
wire _8325_ ;
wire _3880_ ;
wire _3460_ ;
wire _3040_ ;
wire _4665_ ;
wire _4245_ ;
wire _6811_ ;
wire _2731_ ;
wire _2311_ ;
wire _3936_ ;
wire _3516_ ;
wire \datapath.idinstr_22_bF$buf0  ;
wire \datapath.idinstr_16_bF$buf7  ;
wire _8974_ ;
wire _8554_ ;
wire _8134_ ;
wire _4894_ ;
wire _4474_ ;
wire _4054_ ;
wire _913_ ;
wire _5679_ ;
wire _5259_ ;
wire _6620_ ;
wire _6200_ ;
wire _9092_ ;
wire \controlunit.mret_bF$buf2  ;
wire _1599_ ;
wire _1179_ ;
wire _7825_ ;
wire _7405_ ;
wire _2960_ ;
wire _2540_ ;
wire _2120_ ;
wire _3745_ ;
wire _3325_ ;
wire \datapath.idinstr_20_bF$buf7  ;
wire _8783_ ;
wire _8363_ ;
wire _1811_ ;
wire _9148_ ;
wire _4283_ ;
wire _722_ ;
wire _302_ ;
wire _5488_ ;
wire _5068_ ;
wire \datapath.idinstr_22_bF$buf11  ;
wire _7634_ ;
wire _7214_ ;
wire _8839_ ;
wire _8419_ ;
wire _3974_ ;
wire _3554_ ;
wire _3134_ ;
wire [31:0] \datapath.regrs2alu  ;
wire _4759_ ;
wire _4339_ ;
wire _5700_ ;
wire _8592_ ;
wire _8172_ ;
wire \datapath.idinstr_16_bF$buf16  ;
wire _38_ ;
wire _6905_ ;
wire _1620_ ;
wire _1200_ ;
wire _4092_ ;
wire \datapath.idinstr_20_bF$buf31  ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _2825_ ;
wire _2405_ ;
wire _5297_ ;
wire _7863_ ;
wire _7443_ ;
wire _7023_ ;
wire _8648_ ;
wire _8228_ ;
wire _3783_ ;
wire _3363_ ;
wire _4988_ ;
wire _4568_ ;
wire \datapath.idinstr_21_bF$buf40  ;
wire _4148_ ;
wire [31:0] \datapath.idpc_4  ;
wire [31:0] \datapath.meminstr  ;
wire _6714_ ;
wire \datapath.alu.b_0_bF$buf1  ;
wire _9186_ ;
wire _760_ ;
wire _340_ ;
wire _7919_ ;
wire _2634_ ;
wire _2214_ ;
wire \datapath.idinstr_15_bF$buf45  ;
wire _3839_ ;
wire _3419_ ;
wire _7672_ ;
wire _7252_ ;
wire _8877_ ;
wire _8457_ ;
wire _8037_ ;
wire _3592_ ;
wire _3172_ ;
wire _1905_ ;
wire _4797_ ;
wire _4377_ ;
wire _816_ ;
wire _76_ ;
wire _6943_ ;
wire _6523_ ;
wire _6103_ ;
wire _7728_ ;
wire _7308_ ;
wire _2863_ ;
wire _2443_ ;
wire _2023_ ;
wire _3648_ ;
wire _3228_ ;
wire _7481_ ;
wire _7061_ ;
wire _8686_ ;
wire _8266_ ;
wire _1714_ ;
wire _4186_ ;
wire _625_ ;
wire _205_ ;
wire _2919_ ;
wire _6752_ ;
wire _6332_ ;
wire _7957_ ;
wire _7537_ ;
wire _7117_ ;
wire _2672_ ;
wire _2252_ ;
wire _3877_ ;
wire _3457_ ;
wire _3037_ ;
wire _7290_ ;
wire _5603_ ;
wire _8495_ ;
wire _8075_ ;
wire _6808_ ;
wire _1943_ ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire _2728_ ;
wire _2308_ ;
wire _6981_ ;
wire _6561_ ;
wire _6141_ ;
wire \datapath.alu.b_3_bF$buf4  ;
wire _7766_ ;
wire _7346_ ;
wire _2481_ ;
wire _2061_ ;
wire _3686_ ;
wire _3266_ ;
wire _7420__bF$buf10 ;
wire _5832_ ;
wire _5412_ ;
wire _6617_ ;
wire _1752_ ;
wire _1332_ ;
wire _9089_ ;
wire _663_ ;
wire _243_ ;
wire _2957_ ;
wire _2537_ ;
wire _2117_ ;
wire _6790_ ;
wire _6370_ ;
wire _7995_ ;
wire _7575_ ;
wire _7155_ ;
wire _2290_ ;
wire _3495_ ;
wire _3075_ ;
wire _1808_ ;
wire _5641_ ;
wire _5221_ ;
wire _719_ ;
wire _6846_ ;
wire _6426_ ;
wire _6006_ ;
wire _1981_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _2766_ ;
wire _2346_ ;
wire _5152__bF$buf0 ;
wire _5152__bF$buf1 ;
wire _5152__bF$buf2 ;
wire _5152__bF$buf3 ;
wire _5152__bF$buf4 ;
wire _5152__bF$buf5 ;
wire _5152__bF$buf6 ;
wire _5152__bF$buf7 ;
wire _4912_ ;
wire _7384_ ;
wire _8589_ ;
wire _8169_ ;
wire _9110_ ;
wire _1617_ ;
wire _4089_ ;
wire _5870_ ;
wire _5450_ ;
wire _5030_ ;
wire \datapath.idinstr_20_bF$buf28  ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _6655_ ;
wire _6235_ ;
wire _1790_ ;
wire _1370_ ;
wire _281_ ;
wire _2995_ ;
wire _2575_ ;
wire _2155_ ;
wire _8801_ ;
wire _4721_ ;
wire _4301_ ;
wire _7193_ ;
wire \datapath.idinstr_21_bF$buf37  ;
wire _5926_ ;
wire _5506_ ;
wire _8398_ ;
wire _1846_ ;
wire _1426_ ;
wire _1006_ ;
wire _757_ ;
wire _337_ ;
wire _6884_ ;
wire _6464_ ;
wire _6044_ ;
wire \datapath.idinstr_22_hier0_bF$buf3  ;
wire _7669_ ;
wire _7249_ ;
wire _2384_ ;
wire _8610_ ;
wire _3589_ ;
wire _3169_ ;
wire _4950_ ;
wire _4530_ ;
wire _4110_ ;
wire _5735_ ;
wire _5315_ ;
wire _1655_ ;
wire _1235_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire _3801_ ;
wire _6693_ ;
wire _6273_ ;
wire _7898_ ;
wire _7478_ ;
wire _7058_ ;
wire _2193_ ;
wire _5762__bF$buf40 ;
wire _5762__bF$buf41 ;
wire _5762__bF$buf42 ;
wire _5762__bF$buf43 ;
wire _5762__bF$buf44 ;
wire _5762__bF$buf45 ;
wire _5762__bF$buf46 ;
wire _5762__bF$buf47 ;
wire _3398_ ;
wire _5964_ ;
wire _5544_ ;
wire _5124_ ;
wire _6749_ ;
wire _6329_ ;
wire _1884_ ;
wire _1464_ ;
wire _1044_ ;
wire _795_ ;
wire _375_ ;
wire _2669_ ;
wire _2249_ ;
wire _3610_ ;
wire _4839__bF$buf0 ;
wire _6082_ ;
wire _4839__bF$buf1 ;
wire _4839__bF$buf2 ;
wire _4839__bF$buf3 ;
wire _4839__bF$buf4 ;
wire _4815_ ;
wire _7287_ ;
wire _9013_ ;
wire _5773_ ;
wire _5353_ ;
wire [31:0] \datapath.wbpc_4  ;
wire _6978_ ;
wire _6558_ ;
wire _6138_ ;
wire _1693_ ;
wire _1273_ ;
wire _184_ ;
wire _2898_ ;
wire _2478_ ;
wire _2058_ ;
wire _4843__bF$buf0 ;
wire _8704_ ;
wire _4843__bF$buf1 ;
wire _4843__bF$buf2 ;
wire _4843__bF$buf3 ;
wire _4843__bF$buf4 ;
wire _4624_ ;
wire _4204_ ;
wire _7096_ ;
wire _5829_ ;
wire _5409_ ;
wire \datapath.idinstr_16_hier0_bF$buf0  ;
wire _1749_ ;
wire _1329_ ;
wire _5582_ ;
wire _5162_ ;
wire _6787_ ;
wire _6367_ ;
wire _1082_ ;
wire _2287_ ;
wire _8933_ ;
wire _8513_ ;
wire _4853_ ;
wire _4433_ ;
wire _4013_ ;
wire _5638_ ;
wire _5218_ ;
wire _9051_ ;
wire _1978_ ;
wire _1558_ ;
wire _1138_ ;
wire _5391_ ;
wire _889_ ;
wire _469_ ;
wire _3704_ ;
wire _6596_ ;
wire _6176_ ;
wire _4909_ ;
wire _2096_ ;
wire _8742_ ;
wire _8322_ ;
wire _9107_ ;
wire _4662_ ;
wire _4242_ ;
wire _5867_ ;
wire _5447_ ;
wire _5027_ ;
wire _1787_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _3933_ ;
wire _3513_ ;
wire _4718_ ;
wire \datapath.idinstr_16_bF$buf4  ;
wire _8971_ ;
wire _8551_ ;
wire _8131_ ;
wire _4891_ ;
wire _4471_ ;
wire _4051_ ;
wire _910_ ;
wire _5676_ ;
wire _5256_ ;
wire _1596_ ;
wire _1176_ ;
wire _7822_ ;
wire _7402_ ;
wire _8607_ ;
wire _3742_ ;
wire _3322_ ;
wire _4947_ ;
wire \datapath.idinstr_20_bF$buf4  ;
wire _4527_ ;
wire _4107_ ;
wire _8780_ ;
wire _8360_ ;
wire _9145_ ;
wire _4280_ ;
wire _5485_ ;
wire _5065_ ;
wire [31:0] \datapath.programcounter._1_  ;
wire _7631_ ;
wire _7211_ ;
wire _5762__hier0_bF$buf0 ;
wire _5762__hier0_bF$buf1 ;
wire _5762__hier0_bF$buf2 ;
wire _5762__hier0_bF$buf3 ;
wire _5762__hier0_bF$buf4 ;
wire _5762__hier0_bF$buf5 ;
wire _8836_ ;
wire _8416_ ;
wire _3971_ ;
wire _3551_ ;
wire _3131_ ;
wire _4756_ ;
wire _4336_ ;
wire \datapath.idinstr_16_bF$buf13  ;
wire _35_ ;
wire _6902_ ;
wire _2822_ ;
wire _2402_ ;
wire _5294_ ;
wire _3607_ ;
wire _6499_ ;
wire _6079_ ;
wire _7860_ ;
wire _7440_ ;
wire _7020_ ;
wire _8645_ ;
wire _8225_ ;
wire _3780_ ;
wire _3360_ ;
wire _4985_ ;
wire _4565_ ;
wire _4145_ ;
wire _6711_ ;
wire _9183_ ;
wire _7916_ ;
wire _2631_ ;
wire _2211_ ;
wire \datapath.idinstr_15_bF$buf42  ;
wire _3836_ ;
wire _3416_ ;
wire _8874_ ;
wire _8454_ ;
wire _8034_ ;
wire _1902_ ;
wire _4794_ ;
wire _4374_ ;
wire _813_ ;
wire _5999_ ;
wire _5579_ ;
wire _5159_ ;
wire \datapath.idinstr_16_bF$buf51  ;
wire _73_ ;
wire _6940_ ;
wire _6520_ ;
wire _6100_ ;
wire _1499_ ;
wire _1079_ ;
wire _7725_ ;
wire _7305_ ;
wire _2860_ ;
wire _2440_ ;
wire _2020_ ;
wire _3645_ ;
wire _3225_ ;
wire _8683_ ;
wire _8263_ ;
wire _1711_ ;
wire _9048_ ;
wire _4183_ ;
wire _622_ ;
wire _202_ ;
wire _2916_ ;
wire _5388_ ;
wire _7954_ ;
wire _7534_ ;
wire _7114_ ;
wire [31:0] \datapath.registers.838[26]  ;
wire _8739_ ;
wire _8319_ ;
wire _3874_ ;
wire _3454_ ;
wire _3034_ ;
wire _2924__bF$buf0 ;
wire _4659_ ;
wire _2924__bF$buf1 ;
wire _4239_ ;
wire _2924__bF$buf2 ;
wire _2924__bF$buf3 ;
wire _2924__bF$buf4 ;
wire _2924__bF$buf5 ;
wire _2924__bF$buf6 ;
wire _5600_ ;
wire _8492_ ;
wire _8072_ ;
wire _6805_ ;
wire _1940_ ;
wire _1520_ ;
wire _1100_ ;
wire _851_ ;
wire _431_ ;
wire _2725_ ;
wire _2305_ ;
wire _5197_ ;
wire \datapath.alu.b_3_bF$buf1  ;
wire _7763_ ;
wire _7343_ ;
wire _8968_ ;
wire _8548_ ;
wire _8128_ ;
wire \datapath.regwbtrap  ;
wire _3683_ ;
wire _3263_ ;
wire _4888_ ;
wire _4468_ ;
wire _4048_ ;
wire _907_ ;
wire _6614_ ;
wire _9086_ ;
wire _660_ ;
wire _240_ ;
wire _7819_ ;
wire _2954_ ;
wire _2534_ ;
wire _2114_ ;
wire _3739_ ;
wire _3319_ ;
wire _7992_ ;
wire _7572_ ;
wire _7152_ ;
wire _8777_ ;
wire _8357_ ;
wire _3492_ ;
wire _3072_ ;
wire _1805_ ;
wire _4697_ ;
wire _4277_ ;
wire _716_ ;
wire _6843_ ;
wire _6423_ ;
wire _6003_ ;
wire _7628_ ;
wire _7208_ ;
wire _2763_ ;
wire _2343_ ;
wire _3968_ ;
wire _3548_ ;
wire _3128_ ;
wire _7381_ ;
wire _8586_ ;
wire _8166_ ;
wire _1614_ ;
wire _4086_ ;
wire \datapath.idinstr_20_bF$buf25  ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _2819_ ;
wire _6652_ ;
wire _6232_ ;
wire _7857_ ;
wire _7437_ ;
wire _7017_ ;
wire _2992_ ;
wire _2572_ ;
wire _2152_ ;
wire _3777_ ;
wire _3357_ ;
wire _7190_ ;
wire \datapath.idinstr_21_bF$buf34  ;
wire _5923_ ;
wire _5503_ ;
wire _8395_ ;
wire _6708_ ;
wire _1843_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire _2628_ ;
wire _2208_ ;
wire _6881_ ;
wire _6461_ ;
wire _6041_ ;
wire \datapath.idinstr_15_bF$buf39  ;
wire \datapath.idinstr_22_hier0_bF$buf0  ;
wire _7666_ ;
wire _7246_ ;
wire _2381_ ;
wire _3586_ ;
wire _3166_ ;
wire _5732_ ;
wire _5312_ ;
wire \datapath.idinstr_16_bF$buf48  ;
wire _6937_ ;
wire _6517_ ;
wire _1652_ ;
wire _1232_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _2857_ ;
wire _2437_ ;
wire _2017_ ;
wire _6690_ ;
wire _6270_ ;
wire [31:0] \datapath.mempc_4  ;
wire _7895_ ;
wire _7475_ ;
wire _7055_ ;
wire _2190_ ;
wire _5762__bF$buf10 ;
wire _5762__bF$buf11 ;
wire _5762__bF$buf12 ;
wire _5762__bF$buf13 ;
wire _5762__bF$buf14 ;
wire _5762__bF$buf15 ;
wire _5762__bF$buf16 ;
wire _5762__bF$buf17 ;
wire _5762__bF$buf18 ;
wire _5762__bF$buf19 ;
wire _3395_ ;
wire _1708_ ;
wire _5961_ ;
wire _5541_ ;
wire _5121_ ;
wire _619_ ;
wire _6746_ ;
wire _6326_ ;
wire _1881_ ;
wire _1461_ ;
wire _1041_ ;
wire _792_ ;
wire _372_ ;
wire _2666_ ;
wire _2246_ ;
wire _4812_ ;
wire _7284_ ;
wire _8489_ ;
wire _8069_ ;
wire _9010_ ;
wire _1937_ ;
wire _1517_ ;
wire [31:0] \datapath.registers.838[0]  ;
wire _5770_ ;
wire _5350_ ;
wire _848_ ;
wire _428_ ;
wire _6975_ ;
wire _6555_ ;
wire _6135_ ;
wire _1690_ ;
wire _1270_ ;
wire _181_ ;
wire _2895_ ;
wire _2475_ ;
wire _2055_ ;
wire _8701_ ;
wire _4621_ ;
wire _4201_ ;
wire _7093_ ;
wire _5826_ ;
wire _5406_ ;
wire _8298_ ;
wire _1746_ ;
wire _1326_ ;
wire _657_ ;
wire _237_ ;
wire _6784_ ;
wire _6364_ ;
wire _7989_ ;
wire _7569_ ;
wire _7149_ ;
wire _2284_ ;
wire _8930_ ;
wire _8510_ ;
wire _3489_ ;
wire _3069_ ;
wire _4850_ ;
wire _4430_ ;
wire _4010_ ;
wire _5635_ ;
wire _5215_ ;
wire _1975_ ;
wire _1555_ ;
wire _1135_ ;
wire _7425__bF$buf20 ;
wire _7425__bF$buf21 ;
wire _7425__bF$buf22 ;
wire _7425__bF$buf23 ;
wire _7425__bF$buf24 ;
wire _7425__bF$buf25 ;
wire _7425__bF$buf26 ;
wire _7425__bF$buf27 ;
wire _7425__bF$buf28 ;
wire _7425__bF$buf29 ;
wire _886_ ;
wire _466_ ;
wire _3701_ ;
wire _6593_ ;
wire _6173_ ;
wire _4906_ ;
wire _7798_ ;
wire _7378_ ;
wire _2093_ ;
wire _3298_ ;
wire _9104_ ;
wire _5864_ ;
wire _5444_ ;
wire _5024_ ;
wire _6649_ ;
wire _6229_ ;
wire _1784_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _2989_ ;
wire _2569_ ;
wire _2149_ ;
wire _3930_ ;
wire _3510_ ;
wire _4715_ ;
wire _7187_ ;
wire \datapath.idinstr_16_bF$buf1  ;
wire _5673_ ;
wire _5253_ ;
wire _6878_ ;
wire _6458_ ;
wire _6038_ ;
wire _1593_ ;
wire _1173_ ;
wire _2798_ ;
wire _2378_ ;
wire _8604_ ;
wire _4944_ ;
wire \datapath.idinstr_20_bF$buf1  ;
wire _4524_ ;
wire _4104_ ;
wire _5729_ ;
wire _5309_ ;
wire _9142_ ;
wire _1649_ ;
wire _1229_ ;
wire _5482_ ;
wire _5062_ ;
wire [31:0] \datapath.muxbval  ;
wire _6687_ ;
wire _6267_ ;
wire _2187_ ;
wire _8833_ ;
wire _8413_ ;
wire _4753_ ;
wire _4333_ ;
wire _5958_ ;
wire _5538_ ;
wire _5118_ ;
wire \datapath.idinstr_16_bF$buf10  ;
wire _32_ ;
wire _1878_ ;
wire _1458_ ;
wire _1038_ ;
wire _5291_ ;
wire _789_ ;
wire _369_ ;
wire _3604_ ;
wire _6496_ ;
wire _6076_ ;
wire _4809_ ;
wire _8642_ ;
wire _8222_ ;
wire _9007_ ;
wire _4982_ ;
wire _4562_ ;
wire _4142_ ;
wire \datapath.idinstr_19_bF$buf4  ;
wire _5767_ ;
wire _5347_ ;
wire _9180_ ;
wire _1687_ ;
wire _1267_ ;
wire _7913_ ;
wire _598_ ;
wire _178_ ;
wire _3833_ ;
wire _3413_ ;
wire _4618_ ;
wire _8871_ ;
wire _8451_ ;
wire _8031_ ;
wire _4791_ ;
wire _4371_ ;
wire \datapath.idinstr_23_bF$buf4  ;
wire _810_ ;
wire _5996_ ;
wire _5576_ ;
wire _5156_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _7722_ ;
wire _7302_ ;
wire _8927_ ;
wire _8507_ ;
wire _3642_ ;
wire _3222_ ;
wire _4847_ ;
wire _4427_ ;
wire _4007_ ;
wire _8680_ ;
wire _8260_ ;
wire _9045_ ;
wire _4180_ ;
wire _2913_ ;
wire _5385_ ;
wire _7951_ ;
wire _7531_ ;
wire _7111_ ;
wire _8736_ ;
wire _8316_ ;
wire _3871_ ;
wire _3451_ ;
wire _3031_ ;
wire _4656_ ;
wire _4236_ ;
wire _6802_ ;
wire _2722_ ;
wire _2302_ ;
wire _5194_ ;
wire _3927_ ;
wire _3507_ ;
wire _6399_ ;
wire _7760_ ;
wire _7340_ ;
wire _8965_ ;
wire _8545_ ;
wire _8125_ ;
wire _3680_ ;
wire _3260_ ;
wire _4885_ ;
wire _4465_ ;
wire _4045_ ;
wire _904_ ;
wire _6611_ ;
wire _9083_ ;
wire \datapath.regcondt  ;
wire _7816_ ;
wire _2951_ ;
wire _2531_ ;
wire _2111_ ;
wire _3736_ ;
wire _3316_ ;
wire \datapath.alu.b_1_bF$buf5  ;
wire _8774_ ;
wire _8354_ ;
wire _1802_ ;
wire _9139_ ;
wire _4694_ ;
wire _4274_ ;
wire _713_ ;
wire _5899_ ;
wire _5479_ ;
wire _5059_ ;
wire _6840_ ;
wire _6420_ ;
wire _6000_ ;
wire [31:0] \datapath.alu.b  ;
wire _1399_ ;
wire _7625_ ;
wire _7205_ ;
wire _2760_ ;
wire _2340_ ;
wire _3965_ ;
wire _3545_ ;
wire _3125_ ;
wire _8583_ ;
wire _8163_ ;
wire _29_ ;
wire _1611_ ;
wire _4083_ ;
wire \datapath.idinstr_20_bF$buf22  ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _2816_ ;
wire _5288_ ;
wire _7854_ ;
wire _7434_ ;
wire _7014_ ;
wire [31:0] \datapath.registers.838[16]  ;
wire _8639_ ;
wire _8219_ ;
wire _3774_ ;
wire _3354_ ;
wire _4979_ ;
wire _4559_ ;
wire \datapath.idinstr_21_bF$buf31  ;
wire _4139_ ;
wire _5920_ ;
wire _5500_ ;
wire _8392_ ;
wire _6705_ ;
wire _1840_ ;
wire _1420_ ;
wire _1000_ ;
wire _9177_ ;
wire _751_ ;
wire _331_ ;
wire _2625_ ;
wire _2205_ ;
wire _5097_ ;
wire \datapath.idinstr_15_bF$buf36  ;
wire \datapath.idinstr_22_bF$buf40  ;
wire _7663_ ;
wire _7243_ ;
wire _8868_ ;
wire _8448_ ;
wire _8028_ ;
wire _3583_ ;
wire _3163_ ;
wire _4788_ ;
wire _4368_ ;
wire _807_ ;
wire \datapath.idinstr_16_bF$buf45  ;
wire _67_ ;
wire _6934_ ;
wire _6514_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _7719_ ;
wire _2854_ ;
wire _2434_ ;
wire _2014_ ;
wire _3639_ ;
wire _3219_ ;
wire _7892_ ;
wire _7472_ ;
wire _7052_ ;
wire _8677_ ;
wire _8257_ ;
wire _3392_ ;
wire _1705_ ;
wire _4597_ ;
wire _4177_ ;
wire _616_ ;
wire _6743_ ;
wire _6323_ ;
wire _7948_ ;
wire _7528_ ;
wire _7108_ ;
wire _2663_ ;
wire _2243_ ;
wire _3868_ ;
wire _3448_ ;
wire _3028_ ;
wire \datapath.csr.csr_irq  ;
wire _7281_ ;
wire _8486_ ;
wire _8066_ ;
wire _1934_ ;
wire _1514_ ;
wire _5375__bF$buf0 ;
wire _5375__bF$buf1 ;
wire _5375__bF$buf2 ;
wire _5375__bF$buf3 ;
wire _845_ ;
wire _5375__bF$buf4 ;
wire _425_ ;
wire _5375__bF$buf5 ;
wire _5375__bF$buf6 ;
wire _5375__bF$buf7 ;
wire _2719_ ;
wire _6972_ ;
wire _6552_ ;
wire _6132_ ;
wire _7757_ ;
wire _7337_ ;
wire _2892_ ;
wire _2472_ ;
wire _2052_ ;
wire _3677_ ;
wire _3257_ ;
wire _7090_ ;
wire _5823_ ;
wire _5403_ ;
wire _8295_ ;
wire _6608_ ;
wire _1743_ ;
wire _1323_ ;
wire _654_ ;
wire _234_ ;
wire _2948_ ;
wire _2528_ ;
wire _2108_ ;
wire _6781_ ;
wire _6361_ ;
wire _4786__bF$buf0 ;
wire _4786__bF$buf1 ;
wire _4786__bF$buf2 ;
wire _4786__bF$buf3 ;
wire _4786__bF$buf4 ;
wire _7986_ ;
wire _7566_ ;
wire _7146_ ;
wire _2281_ ;
wire _3486_ ;
wire _3066_ ;
wire _5632_ ;
wire _5212_ ;
wire _6837_ ;
wire _6417_ ;
wire _1972_ ;
wire _1552_ ;
wire _1132_ ;
wire _883_ ;
wire _463_ ;
wire _2757_ ;
wire _2337_ ;
wire _6590_ ;
wire _6170_ ;
wire _4903_ ;
wire _7795_ ;
wire _7375_ ;
wire _2090_ ;
wire _3295_ ;
wire _9101_ ;
wire _1608_ ;
wire _5861_ ;
wire _5441_ ;
wire _5021_ ;
wire \datapath.idinstr_20_bF$buf19  ;
wire _939_ ;
wire _519_ ;
wire _6646_ ;
wire _6226_ ;
wire _1781_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _2986_ ;
wire _2566_ ;
wire _2146_ ;
wire _4712_ ;
wire _7184_ ;
wire \datapath.idinstr_21_bF$buf28  ;
wire _5917_ ;
wire _8389_ ;
wire _1837_ ;
wire _1417_ ;
wire _5670_ ;
wire _5250_ ;
wire _748_ ;
wire _328_ ;
wire _6875_ ;
wire _6455_ ;
wire _6035_ ;
wire _1590_ ;
wire _1170_ ;
wire \datapath.idinstr_22_bF$buf37  ;
wire _2795_ ;
wire _2375_ ;
wire _8601_ ;
wire _4941_ ;
wire _4521_ ;
wire _4101_ ;
wire _5726_ ;
wire _5306_ ;
wire _8198_ ;
wire _1646_ ;
wire _1226_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire _6684_ ;
wire _6264_ ;
wire [31:0] \datapath.aluinstr  ;
wire _7889_ ;
wire _7469_ ;
wire _7049_ ;
wire _2184_ ;
wire _8830_ ;
wire _8410_ ;
wire _3389_ ;
wire _4750_ ;
wire _4330_ ;
wire _5955_ ;
wire _5535_ ;
wire _5115_ ;
wire _1875_ ;
wire _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire _3601_ ;
wire _6493_ ;
wire _6073_ ;
wire _4806_ ;
wire _7698_ ;
wire _7278_ ;
wire _3198_ ;
wire _5442__bF$buf0 ;
wire _5442__bF$buf1 ;
wire _5442__bF$buf2 ;
wire _5442__bF$buf3 ;
wire _5442__bF$buf4 ;
wire _5442__bF$buf5 ;
wire _5442__bF$buf6 ;
wire _5442__bF$buf7 ;
wire _9004_ ;
wire \datapath.idinstr_19_bF$buf1  ;
wire _5764_ ;
wire _5344_ ;
wire _4849__bF$buf0 ;
wire _4849__bF$buf1 ;
wire _4849__bF$buf2 ;
wire _4849__bF$buf3 ;
wire _4849__bF$buf4 ;
wire _6969_ ;
wire _6549_ ;
wire _6129_ ;
wire _1684_ ;
wire _1264_ ;
wire _7910_ ;
wire _595_ ;
wire _175_ ;
wire _2889_ ;
wire _2469_ ;
wire _2049_ ;
wire _3830_ ;
wire _3410_ ;
wire _4615_ ;
wire _7087_ ;
wire \datapath.idinstr_23_bF$buf1  ;
wire _5993_ ;
wire _5573_ ;
wire _5153_ ;
wire _4853__bF$buf0 ;
wire _4853__bF$buf1 ;
wire _4853__bF$buf2 ;
wire _4853__bF$buf3 ;
wire _4853__bF$buf4 ;
wire _6778_ ;
wire _6358_ ;
wire _1493_ ;
wire _1073_ ;
wire _2698_ ;
wire _2278_ ;
wire _8924_ ;
wire _8504_ ;
wire _4844_ ;
wire _4424_ ;
wire _4004_ ;
wire _5629_ ;
wire _5209_ ;
wire _9042_ ;
wire _1969_ ;
wire _1549_ ;
wire _1129_ ;
wire _2910_ ;
wire _5382_ ;
wire _6587_ ;
wire _6167_ ;
wire _2087_ ;
wire _8733_ ;
wire _8313_ ;
wire _4653_ ;
wire _4233_ ;
wire _5858_ ;
wire _5438_ ;
wire _5018_ ;
wire _1833__bF$buf0 ;
wire _1833__bF$buf1 ;
wire _1833__bF$buf2 ;
wire _1833__bF$buf3 ;
wire _1833__bF$buf4 ;
wire _1833__bF$buf5 ;
wire _1833__bF$buf6 ;
wire _1833__bF$buf7 ;
wire _1778_ ;
wire _1358_ ;
wire _5191_ ;
wire _689_ ;
wire _269_ ;
wire [31:0] \datapath.registers.838[31]  ;
wire _3924_ ;
wire _3504_ ;
wire _6396_ ;
wire _4709_ ;
wire _8962_ ;
wire _8542_ ;
wire _8122_ ;
wire _4882_ ;
wire _4462_ ;
wire _4042_ ;
wire _901_ ;
wire _5667_ ;
wire _5247_ ;
wire _9080_ ;
wire _1587_ ;
wire [31:0] \datapath.registers.838[7]  ;
wire _1167_ ;
wire _7813_ ;
wire _498_ ;
wire _3733_ ;
wire _3313_ ;
wire \datapath.alu.b_1_bF$buf2  ;
wire _288__bF$buf0 ;
wire _288__bF$buf1 ;
wire _288__bF$buf2 ;
wire _288__bF$buf3 ;
wire _288__bF$buf4 ;
wire _4938_ ;
wire _4518_ ;
wire _8771_ ;
wire _8351_ ;
wire _9136_ ;
wire _4691_ ;
wire _4271_ ;
wire _710_ ;
wire _5896_ ;
wire _5476_ ;
wire _5056_ ;
wire _1396_ ;
wire _7622_ ;
wire _7202_ ;
wire _8827_ ;
wire _8407_ ;
wire _3962_ ;
wire _3542_ ;
wire _3122_ ;
wire _4747_ ;
wire _4327_ ;
wire _386__bF$buf0 ;
wire _386__bF$buf1 ;
wire _386__bF$buf2 ;
wire _386__bF$buf3 ;
wire _386__bF$buf4 ;
wire _8580_ ;
wire _8160_ ;
wire _26_ ;
wire _4080_ ;
wire _2813_ ;
wire _5285_ ;
wire _7851_ ;
wire _7431_ ;
wire _7011_ ;
wire _8636_ ;
wire _8216_ ;
wire _3771_ ;
wire _3351_ ;
wire \datapath.idinstr_17_bF$buf13  ;
wire _4976_ ;
wire _4556_ ;
wire _4136_ ;
wire _6702_ ;
wire _9174_ ;
wire _7907_ ;
wire _2622_ ;
wire _2202_ ;
wire _5094_ ;
wire \datapath.idinstr_15_bF$buf33  ;
wire _3827_ ;
wire _3407_ ;
wire _6299_ ;
wire _7660_ ;
wire _7240_ ;
wire _8865_ ;
wire _8445_ ;
wire _8025_ ;
wire _3580_ ;
wire _3160_ ;
wire _4785_ ;
wire _4365_ ;
wire _804_ ;
wire \datapath.idinstr_16_bF$buf42  ;
wire _64_ ;
wire _6931_ ;
wire _6511_ ;
wire _7716_ ;
wire _2851_ ;
wire _2431_ ;
wire _2011_ ;
wire _3636_ ;
wire _3216_ ;
wire _8674_ ;
wire _8254_ ;
wire \controlunit.csrfile_trap_wen  ;
wire _1702_ ;
wire _9039_ ;
wire _4594_ ;
wire _4174_ ;
wire _613_ ;
wire _2907_ ;
wire _5799_ ;
wire _5379_ ;
wire _6740_ ;
wire _6320_ ;
wire _1299_ ;
wire _7945_ ;
wire _7525_ ;
wire _7105_ ;
wire _2660_ ;
wire _2240_ ;
wire _3865_ ;
wire _3445_ ;
wire _3025_ ;
wire _8483_ ;
wire CLK_bF$buf90 ;
wire _8063_ ;
wire CLK_bF$buf91 ;
wire CLK_bF$buf92 ;
wire CLK_bF$buf93 ;
wire CLK_bF$buf94 ;
wire CLK_bF$buf95 ;
wire CLK_bF$buf96 ;
wire CLK_bF$buf97 ;
wire CLK_bF$buf98 ;
wire CLK_bF$buf99 ;
wire _1931_ ;
wire _1511_ ;
wire _842_ ;
wire _422_ ;
wire _2716_ ;
wire _5188_ ;
wire _7754_ ;
wire _7334_ ;
wire _8959_ ;
wire _8539_ ;
wire _8119_ ;
wire _3674_ ;
wire _3254_ ;
wire _4879_ ;
wire _4459_ ;
wire _4039_ ;
wire _5820_ ;
wire _5400_ ;
wire _8292_ ;
wire _4801__bF$buf0 ;
wire _4801__bF$buf1 ;
wire _4801__bF$buf2 ;
wire _4801__bF$buf3 ;
wire _4801__bF$buf4 ;
wire _6605_ ;
wire _1740_ ;
wire _1320_ ;
wire _9077_ ;
wire _651_ ;
wire _231_ ;
wire _2945_ ;
wire _2525_ ;
wire _2105_ ;
wire _7983_ ;
wire _7563_ ;
wire _7143_ ;
wire _8768_ ;
wire _8348_ ;
wire _3483_ ;
wire _3063_ ;
wire _4688_ ;
wire _4268_ ;
wire _707_ ;
wire _6834_ ;
wire _6414_ ;
wire \controlunit.ecall  ;
wire _880_ ;
wire _460_ ;
wire _7619_ ;
wire _2754_ ;
wire _2334_ ;
wire _3959_ ;
wire _3539_ ;
wire _3119_ ;
wire _4900_ ;
wire _7792_ ;
wire _7372_ ;
wire _8997_ ;
wire _8577_ ;
wire _8157_ ;
wire _3292_ ;
wire _1605_ ;
wire _4497_ ;
wire _4077_ ;
wire \datapath.idinstr_20_bF$buf16  ;
wire _936_ ;
wire _516_ ;
wire _6643_ ;
wire _6223_ ;
wire _7848_ ;
wire _7428_ ;
wire _7008_ ;
wire _2983_ ;
wire _2563_ ;
wire _2143_ ;
wire _3768_ ;
wire _3348_ ;
wire _7181_ ;
wire \datapath.idinstr_21_bF$buf25  ;
wire _5914_ ;
wire _8386_ ;
wire _1834_ ;
wire _1414_ ;
wire _745_ ;
wire _325_ ;
wire _2619_ ;
wire _6872_ ;
wire _6452_ ;
wire _6032_ ;
wire \datapath.idinstr_22_bF$buf34  ;
wire _7657_ ;
wire _7237_ ;
wire _2792_ ;
wire _2372_ ;
wire _3997_ ;
wire _3577_ ;
wire _3157_ ;
wire _4935__bF$buf0 ;
wire _4935__bF$buf1 ;
wire _4935__bF$buf2 ;
wire _4935__bF$buf3 ;
wire _4935__bF$buf4 ;
wire _4935__bF$buf5 ;
wire _4935__bF$buf6 ;
wire _4935__bF$buf7 ;
wire _5723_ ;
wire _5303_ ;
wire _8195_ ;
wire \datapath.idinstr_16_bF$buf39  ;
wire _6928_ ;
wire _6508_ ;
wire _1643_ ;
wire _1223_ ;
wire \datapath.idinstr_20_bF$buf54  ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire _2848_ ;
wire _2428_ ;
wire _2008_ ;
wire _6681_ ;
wire _6261_ ;
wire _7886_ ;
wire _7466_ ;
wire _7046_ ;
wire _2181_ ;
wire _3386_ ;
wire _5952_ ;
wire _5532_ ;
wire _5112_ ;
wire _6737_ ;
wire _6317_ ;
wire _1872_ ;
wire _1452_ ;
wire _1032_ ;
wire _783_ ;
wire _363_ ;
wire _2657_ ;
wire _2237_ ;
wire _6490_ ;
wire _6070_ ;
wire _4803_ ;
wire _7695_ ;
wire _7275_ ;
wire _3195_ ;
wire _9001_ ;
wire _1928_ ;
wire _1508_ ;
wire _5761_ ;
wire _5341_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _6966_ ;
wire _6546_ ;
wire _6126_ ;
wire _1681_ ;
wire _1261_ ;
wire _592_ ;
wire _172_ ;
wire _2886_ ;
wire _2466_ ;
wire _2046_ ;
wire _4612_ ;
wire _7084_ ;
wire _5817_ ;
wire _8289_ ;
wire _1737_ ;
wire _1317_ ;
wire _5990_ ;
wire _5570_ ;
wire _5150_ ;
wire _648_ ;
wire _228_ ;
wire _6775_ ;
wire _6355_ ;
wire _1490_ ;
wire _1070_ ;
wire _5756__bF$buf0 ;
wire _5756__bF$buf1 ;
wire _5756__bF$buf2 ;
wire _5756__bF$buf3 ;
wire _5756__bF$buf4 ;
wire _5756__bF$buf5 ;
wire _5756__bF$buf6 ;
wire _5756__bF$buf7 ;
wire _5756__bF$buf8 ;
wire _5756__bF$buf9 ;
wire _2695_ ;
wire _2275_ ;
wire _8921_ ;
wire _8501_ ;
wire _4841_ ;
wire _4421_ ;
wire _4001_ ;
wire _5626_ ;
wire _5206_ ;
wire _8098_ ;
wire _1966_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire _6584_ ;
wire _6164_ ;
wire _5760__bF$buf0 ;
wire _5760__bF$buf1 ;
wire _5760__bF$buf2 ;
wire _5760__bF$buf3 ;
wire _5760__bF$buf4 ;
wire _5760__bF$buf5 ;
wire _5760__bF$buf6 ;
wire _5760__bF$buf7 ;
wire _7789_ ;
wire _7369_ ;
wire _2084_ ;
wire _8730_ ;
wire _8310_ ;
wire \datapath.immediatedecoder._12_  ;
wire _3289_ ;
wire _4650_ ;
wire _4230_ ;
wire _5855_ ;
wire _5435_ ;
wire _5015_ ;
wire _1775_ ;
wire _1355_ ;
wire _686_ ;
wire [31:0] \datapath.imm  ;
wire _266_ ;
wire _3921_ ;
wire _3501_ ;
wire _6393_ ;
wire _4706_ ;
wire _7598_ ;
wire _7178_ ;
wire _3014__bF$buf0 ;
wire _3014__bF$buf1 ;
wire _3014__bF$buf2 ;
wire _3014__bF$buf3 ;
wire _3014__bF$buf4 ;
wire _3014__bF$buf5 ;
wire _3014__bF$buf6 ;
wire _3098_ ;
wire [31:0] \datapath.regimmalu  ;
wire _5664_ ;
wire _5244_ ;
wire \datapath.idinstr_17_bF$buf7  ;
wire _6869_ ;
wire _6449_ ;
wire _6029_ ;
wire _1584_ ;
wire _1164_ ;
wire _7810_ ;
wire CLK ;
wire _495_ ;
wire _2789_ ;
wire _2369_ ;
wire _3730_ ;
wire _3310_ ;
wire _4935_ ;
wire _4515_ ;
wire _9133_ ;
wire \datapath.idinstr_21_bF$buf7  ;
wire _5893_ ;
wire _5473_ ;
wire _5053_ ;
wire _6678_ ;
wire _6258_ ;
wire _1393_ ;
wire _2598_ ;
wire _2178_ ;
wire _8824_ ;
wire _8404_ ;
wire _4744_ ;
wire _4324_ ;
wire _5949_ ;
wire _5529_ ;
wire _5109_ ;
wire _23_ ;
wire _1869_ ;
wire _1449_ ;
wire _1029_ ;
wire _2810_ ;
wire _5282_ ;
wire _6487_ ;
wire _6067_ ;
wire _8633_ ;
wire _8213_ ;
wire \datapath.idinstr_17_bF$buf10  ;
wire _4973_ ;
wire _4553_ ;
wire _4133_ ;
wire _5758_ ;
wire _5338_ ;
wire _9171_ ;
wire _1678_ ;
wire _1258_ ;
wire _7904_ ;
wire _5091_ ;
wire _589_ ;
wire _169_ ;
wire [31:0] \datapath.registers.838[21]  ;
wire \datapath.idinstr_15_bF$buf30  ;
wire _3824_ ;
wire _3404_ ;
wire _6296_ ;
wire _4609_ ;
wire _8862_ ;
wire _8442_ ;
wire _8022_ ;
wire \datapath.alu.b_4_bF$buf2  ;
wire _4782_ ;
wire _4362_ ;
wire _801_ ;
wire _5987_ ;
wire _5567_ ;
wire _5147_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _7713_ ;
wire _398_ ;
wire _8918_ ;
wire _3633_ ;
wire _3213_ ;
wire _4838_ ;
wire _4418_ ;
wire _4899__bF$buf10 ;
wire _4899__bF$buf11 ;
wire _4899__bF$buf12 ;
wire _4899__bF$buf13 ;
wire _8671_ ;
wire _8251_ ;
wire _9036_ ;
wire _4591_ ;
wire _4171_ ;
wire _610_ ;
wire _2904_ ;
wire _5796_ ;
wire _5376_ ;
wire _1296_ ;
wire _7942_ ;
wire _7522_ ;
wire _7102_ ;
wire _8727_ ;
wire _8307_ ;
wire _3862_ ;
wire _3442_ ;
wire _3022_ ;
wire _4647_ ;
wire _4227_ ;
wire _8480_ ;
wire CLK_bF$buf60 ;
wire _8060_ ;
wire CLK_bF$buf61 ;
wire CLK_bF$buf62 ;
wire CLK_bF$buf63 ;
wire CLK_bF$buf64 ;
wire CLK_bF$buf65 ;
wire CLK_bF$buf66 ;
wire CLK_bF$buf67 ;
wire CLK_bF$buf68 ;
wire CLK_bF$buf69 ;
wire _2713_ ;
wire _5185_ ;
wire [31:0] \datapath.rd  ;
wire _3918_ ;
wire _7751_ ;
wire _7331_ ;
wire _8956_ ;
wire _8536_ ;
wire _8116_ ;
wire _3671_ ;
wire _3251_ ;
wire _4876_ ;
wire _4456_ ;
wire _4036_ ;
wire _6602_ ;
wire _9074_ ;
wire _7807_ ;
wire _2942_ ;
wire _2522_ ;
wire _2102_ ;
wire _3727_ ;
wire _3307_ ;
wire _6199_ ;
wire _7980_ ;
wire _7560_ ;
wire _7140_ ;
wire _8765_ ;
wire _8345_ ;
wire _3480_ ;
wire _3060_ ;
wire _4685_ ;
wire _4265_ ;
wire _704_ ;
wire _6831_ ;
wire _6411_ ;
wire _7616_ ;
wire _2751_ ;
wire _2331_ ;
wire _3956_ ;
wire _3536_ ;
wire _3116_ ;
wire _8994_ ;
wire _8574_ ;
wire _8154_ ;
wire _1602_ ;
wire _4494_ ;
wire _4074_ ;
wire \datapath.idinstr_20_bF$buf13  ;
wire _933_ ;
wire _513_ ;
wire _2807_ ;
wire _5699_ ;
wire _5279_ ;
wire _6640_ ;
wire _6220_ ;
wire _1199_ ;
wire _7845_ ;
wire _7425_ ;
wire _7005_ ;
wire _2980_ ;
wire _2560_ ;
wire _2140_ ;
wire _3765_ ;
wire _3345_ ;
wire \datapath.idinstr_21_bF$buf22  ;
wire _5911_ ;
wire _8383_ ;
wire _5757__bF$buf10 ;
wire _1831_ ;
wire _1411_ ;
wire _9168_ ;
wire _742_ ;
wire _322_ ;
wire _2616_ ;
wire _5088_ ;
wire \datapath.idinstr_15_bF$buf27  ;
wire \datapath.idinstr_22_bF$buf31  ;
wire _7654_ ;
wire _7234_ ;
wire _8859_ ;
wire _8439_ ;
wire _8019_ ;
wire _3994_ ;
wire _3574_ ;
wire _3154_ ;
wire [31:0] IMEM_ADDR ;
wire _2133__bF$buf0 ;
wire _2133__bF$buf1 ;
wire _2133__bF$buf2 ;
wire _2133__bF$buf3 ;
wire _4779_ ;
wire _4359_ ;
wire _5720_ ;
wire _5300_ ;
wire _8192_ ;
wire \datapath.idinstr_16_bF$buf36  ;
wire _58_ ;
wire _6925_ ;
wire _6505_ ;
wire _1640_ ;
wire _1220_ ;
wire \datapath.idinstr_20_bF$buf51  ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _2845_ ;
wire _2425_ ;
wire _2005_ ;
wire _7883_ ;
wire _7463_ ;
wire _7043_ ;
wire _8668_ ;
wire _8248_ ;
wire _3383_ ;
wire _4588_ ;
wire _4168_ ;
wire _607_ ;
wire _6734_ ;
wire _6314_ ;
wire _780_ ;
wire _360_ ;
wire _7939_ ;
wire _7519_ ;
wire _2654_ ;
wire _2234_ ;
wire _3859_ ;
wire _3439_ ;
wire _3019_ ;
wire _4800_ ;
wire _7692_ ;
wire _7272_ ;
wire _8897_ ;
wire _8477_ ;
wire _8057_ ;
wire _3192_ ;
wire _1925_ ;
wire _1505_ ;
wire _4397_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _6963_ ;
wire _6543_ ;
wire _6123_ ;
wire _7748_ ;
wire _7328_ ;
wire _2883_ ;
wire _2463_ ;
wire _2043_ ;
wire _3668_ ;
wire _3248_ ;
wire _7081_ ;
wire _5814_ ;
wire _8286_ ;
wire _1734_ ;
wire _1314_ ;
wire _645_ ;
wire _225_ ;
wire _2939_ ;
wire _2519_ ;
wire _6772_ ;
wire _6352_ ;
wire _7977_ ;
wire _7557_ ;
wire _7137_ ;
wire _2692_ ;
wire _2272_ ;
wire _3897_ ;
wire _3477_ ;
wire _3057_ ;
wire _5623_ ;
wire _5203_ ;
wire _8095_ ;
wire _6828_ ;
wire _6408_ ;
wire _1963_ ;
wire _1543_ ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _2748_ ;
wire _2328_ ;
wire _6581_ ;
wire _6161_ ;
wire _7786_ ;
wire _7366_ ;
wire _2081_ ;
wire _3286_ ;
wire _5852_ ;
wire _5432_ ;
wire _5012_ ;
wire _6637_ ;
wire _6217_ ;
wire _1772_ ;
wire _1352_ ;
wire _683_ ;
wire _263_ ;
wire _2977_ ;
wire _2557_ ;
wire _2137_ ;
wire _6390_ ;
wire _4703_ ;
wire _7595_ ;
wire _7175_ ;
wire \datapath.idinstr_21_bF$buf19  ;
wire _5908_ ;
wire _3095_ ;
wire _1828_ ;
wire _1408_ ;
wire _5661_ ;
wire _5241_ ;
wire _739_ ;
wire _319_ ;
wire \datapath.idinstr_17_bF$buf4  ;
wire _6866_ ;
wire _6446_ ;
wire _6026_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire \datapath.idinstr_22_bF$buf28  ;
wire _2786_ ;
wire _2366_ ;
wire _4932_ ;
wire _4512_ ;
wire _5717_ ;
wire _8189_ ;
wire _9130_ ;
wire _1637_ ;
wire _1217_ ;
wire \datapath.idinstr_21_bF$buf4  ;
wire _5890_ ;
wire _5470_ ;
wire _5050_ ;
wire \datapath.idinstr_20_bF$buf48  ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _6675_ ;
wire _6255_ ;
wire _1390_ ;
wire _2595_ ;
wire _2175_ ;
wire _8821_ ;
wire _8401_ ;
wire _4741_ ;
wire _4321_ ;
wire _5946_ ;
wire _5526_ ;
wire _5106_ ;
wire _20_ ;
wire _1866_ ;
wire _1446_ ;
wire _1026_ ;
wire _777_ ;
wire _357_ ;
wire _6484_ ;
wire _6064_ ;
wire _7689_ ;
wire _7269_ ;
wire _8630_ ;
wire _8210_ ;
wire _3189_ ;
wire _4970_ ;
wire _4550_ ;
wire _4130_ ;
wire _5755_ ;
wire _5335_ ;
wire _3017__bF$buf0 ;
wire _3017__bF$buf1 ;
wire _3017__bF$buf2 ;
wire _3017__bF$buf3 ;
wire _3017__bF$buf4 ;
wire _1675_ ;
wire _1255_ ;
wire _7901_ ;
wire _586_ ;
wire _166_ ;
wire _3821_ ;
wire _3401_ ;
wire _6293_ ;
wire _4606_ ;
wire _7498_ ;
wire _7078_ ;
wire _4859__bF$buf0 ;
wire _4859__bF$buf1 ;
wire _4859__bF$buf2 ;
wire _4859__bF$buf3 ;
wire _4859__bF$buf4 ;
wire _5984_ ;
wire _5564_ ;
wire _5144_ ;
wire _6769_ ;
wire _6349_ ;
wire _1484_ ;
wire _1064_ ;
wire _7710_ ;
wire _395_ ;
wire _2689_ ;
wire _2269_ ;
wire _8915_ ;
wire [31:0] \datapath.programcounter.jumps  ;
wire _3630_ ;
wire _3210_ ;
wire _4835_ ;
wire _4415_ ;
wire _4863__bF$buf0 ;
wire _4863__bF$buf1 ;
wire _4863__bF$buf2 ;
wire _4863__bF$buf3 ;
wire _4863__bF$buf4 ;
wire _4863__bF$buf5 ;
wire _4863__bF$buf6 ;
wire _4863__bF$buf7 ;
wire _9033_ ;
wire \datapath.alu.b_2_bF$buf6  ;
wire _2901_ ;
wire _5793_ ;
wire _5373_ ;
wire _6998_ ;
wire _6578_ ;
wire _6158_ ;
wire _1293_ ;
wire _2498_ ;
wire _2078_ ;
wire _8724_ ;
wire _8304_ ;
wire _1839__bF$buf0 ;
wire _1839__bF$buf1 ;
wire _1839__bF$buf2 ;
wire _1839__bF$buf3 ;
wire _1839__bF$buf4 ;
wire _1839__bF$buf5 ;
wire _1839__bF$buf6 ;
wire _4644_ ;
wire _4224_ ;
wire CLK_bF$buf30 ;
wire CLK_bF$buf31 ;
wire CLK_bF$buf32 ;
wire CLK_bF$buf33 ;
wire CLK_bF$buf34 ;
wire CLK_bF$buf35 ;
wire CLK_bF$buf36 ;
wire CLK_bF$buf37 ;
wire CLK_bF$buf38 ;
wire CLK_bF$buf39 ;
wire _5849_ ;
wire _5429_ ;
wire _5009_ ;
wire _1769_ ;
wire _1349_ ;
wire _2710_ ;
wire _5182_ ;
wire _3915_ ;
wire _6387_ ;
wire _8953_ ;
wire _8533_ ;
wire _8113_ ;
wire _4873_ ;
wire _4453_ ;
wire _4033_ ;
wire _5658_ ;
wire _5238_ ;
wire _9071_ ;
wire _1998_ ;
wire _1578_ ;
wire _1158_ ;
wire _7804_ ;
wire _489_ ;
wire [31:0] \datapath.registers.838[11]  ;
wire _3724_ ;
wire _3304_ ;
wire _6196_ ;
wire _4929_ ;
wire _4509_ ;
wire _8762_ ;
wire _8342_ ;
wire _9127_ ;
wire _4682_ ;
wire _4262_ ;
wire _701_ ;
wire _5887_ ;
wire _5467_ ;
wire _5047_ ;
wire _1387_ ;
wire _7613_ ;
wire _298_ ;
wire \datapath.idinstr_20_hier0_bF$buf5  ;
wire _8818_ ;
wire _3953_ ;
wire _3533_ ;
wire _3113_ ;
wire _4738_ ;
wire _4318_ ;
wire _8991_ ;
wire _8571_ ;
wire _8151_ ;
wire _17_ ;
wire _4491_ ;
wire _4071_ ;
wire \datapath.idinstr_20_bF$buf10  ;
wire _930_ ;
wire _510_ ;
wire _2804_ ;
wire _5696_ ;
wire _5276_ ;
wire _1196_ ;
wire _7842_ ;
wire _7422_ ;
wire _7002_ ;
wire _8627_ ;
wire _8207_ ;
wire _3762_ ;
wire _3342_ ;
wire _4967_ ;
wire _4547_ ;
wire _4127_ ;
wire _8380_ ;
wire _9165_ ;
wire _2613_ ;
wire _5085_ ;
wire \datapath.idinstr_15_bF$buf24  ;
wire _3818_ ;
wire _7651_ ;
wire _7231_ ;
wire _8856_ ;
wire _8436_ ;
wire _8016_ ;
wire _3991_ ;
wire _3571_ ;
wire _3151_ ;
wire _4776_ ;
wire _4356_ ;
wire \datapath.idinstr_16_bF$buf33  ;
wire _55_ ;
wire _6922_ ;
wire _6502_ ;
wire _7707_ ;
wire _2842_ ;
wire _2422_ ;
wire _2002_ ;
wire _3627_ ;
wire _3207_ ;
wire _6099_ ;
wire _7880_ ;
wire _7460_ ;
wire _7040_ ;
wire _8665_ ;
wire _8245_ ;
wire _3380_ ;
wire _4585_ ;
wire _4165_ ;
wire _604_ ;
wire _6731_ ;
wire _6311_ ;
wire _7936_ ;
wire _7516_ ;
wire _2651_ ;
wire _2231_ ;
wire _3856_ ;
wire _3436_ ;
wire _3016_ ;
wire _8894_ ;
wire _8474_ ;
wire _8054_ ;
wire _1922_ ;
wire _1502_ ;
wire _4394_ ;
wire _833_ ;
wire _413_ ;
wire _2707_ ;
wire _5599_ ;
wire _5179_ ;
wire _93_ ;
wire _6960_ ;
wire _6540_ ;
wire _6120_ ;
wire _1099_ ;
wire _7745_ ;
wire _7325_ ;
wire _2880_ ;
wire _2460_ ;
wire _2040_ ;
wire _3665_ ;
wire _3245_ ;
wire _4807__bF$buf0 ;
wire _4807__bF$buf1 ;
wire _4807__bF$buf2 ;
wire _4807__bF$buf3 ;
wire _4807__bF$buf4 ;
wire _5811_ ;
wire _8283_ ;
wire _1731_ ;
wire _1311_ ;
wire _9068_ ;
wire _642_ ;
wire _222_ ;
wire _2936_ ;
wire _2516_ ;
wire _7974_ ;
wire _7554_ ;
wire _7134_ ;
wire _4811__bF$buf0 ;
wire _4811__bF$buf1 ;
wire [31:0] \datapath.registers.838[28]  ;
wire _4811__bF$buf2 ;
wire _4811__bF$buf3 ;
wire _4811__bF$buf4 ;
wire _8759_ ;
wire _8339_ ;
wire _3894_ ;
wire _3474_ ;
wire _3054_ ;
wire _4679_ ;
wire _4259_ ;
wire _5620_ ;
wire _5200_ ;
wire _8092_ ;
wire _6825_ ;
wire _6405_ ;
wire _1960_ ;
wire _1540_ ;
wire _1120_ ;
wire _871_ ;
wire _451_ ;
wire _2745_ ;
wire _2325_ ;
wire _7783_ ;
wire _7363_ ;
wire _8988_ ;
wire _8568_ ;
wire _8148_ ;
wire _3283_ ;
wire _4488_ ;
wire _4068_ ;
wire _927_ ;
wire _507_ ;
wire _6634_ ;
wire _6214_ ;
wire _680_ ;
wire _260_ ;
wire _7839_ ;
wire _7419_ ;
wire _2974_ ;
wire _2554_ ;
wire _2134_ ;
wire _3759_ ;
wire _3339_ ;
wire _4700_ ;
wire _7592_ ;
wire _7172_ ;
wire \datapath.idinstr_21_bF$buf16  ;
wire _5905_ ;
wire _8797_ ;
wire _8377_ ;
wire _3092_ ;
wire _1825_ ;
wire _1405_ ;
wire _4297_ ;
wire _736_ ;
wire _316_ ;
wire \datapath.idinstr_17_bF$buf1  ;
wire _6863_ ;
wire _6443_ ;
wire _6023_ ;
wire \datapath.idinstr_22_bF$buf25  ;
wire _7648_ ;
wire _7228_ ;
wire _2783_ ;
wire _2363_ ;
wire _3988_ ;
wire _3568_ ;
wire _3148_ ;
wire _5714_ ;
wire _8186_ ;
wire _6919_ ;
wire _1634_ ;
wire _1214_ ;
wire \datapath.idinstr_21_bF$buf1  ;
wire \datapath.idinstr_20_bF$buf45  ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _2839_ ;
wire \datapath.idinstr_15_bF$buf8  ;
wire _2419_ ;
wire _6672_ ;
wire _6252_ ;
wire _4799__bF$buf0 ;
wire _4799__bF$buf1 ;
wire _4799__bF$buf2 ;
wire _4799__bF$buf3 ;
wire _4799__bF$buf4 ;
wire _4799__bF$buf5 ;
wire _4799__bF$buf6 ;
wire _4799__bF$buf7 ;
wire _7877_ ;
wire _7457_ ;
wire _7037_ ;
wire _2592_ ;
wire _2172_ ;
wire _3797_ ;
wire _3377_ ;
wire _5943_ ;
wire _5523_ ;
wire _5103_ ;
wire _6728_ ;
wire _6308_ ;
wire _1863_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _2648_ ;
wire _2228_ ;
wire _6481_ ;
wire _6061_ ;
wire _7686_ ;
wire _7266_ ;
wire _3186_ ;
wire _1919_ ;
wire _5752_ ;
wire _5332_ ;
wire _6957_ ;
wire _6537_ ;
wire _6117_ ;
wire _1672_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _2877_ ;
wire _2457_ ;
wire _2037_ ;
wire _6290_ ;
wire _4603_ ;
wire _7495_ ;
wire _7075_ ;
wire _5808_ ;
wire _1728_ ;
wire _1308_ ;
wire _5981_ ;
wire _5561_ ;
wire _5141_ ;
wire _639_ ;
wire _219_ ;
wire [31:0] DMEM_ADDR ;
wire _6766_ ;
wire _6346_ ;
wire _1481_ ;
wire _1061_ ;
wire _392_ ;
wire \datapath.idinstr_24_bF$buf4  ;
wire _2686_ ;
wire _2266_ ;
wire _8912_ ;
wire _4832_ ;
wire _4412_ ;
wire _5617_ ;
wire _8089_ ;
wire _9030_ ;
wire \datapath.alu.b_2_bF$buf3  ;
wire _1957_ ;
wire _1537_ ;
wire [31:0] \datapath.registers.838[2]  ;
wire _1117_ ;
wire _5790_ ;
wire _5370_ ;
wire _868_ ;
wire _448_ ;
wire _6995_ ;
wire _6575_ ;
wire _6155_ ;
wire _1290_ ;
wire _2495_ ;
wire _2075_ ;
wire _8721_ ;
wire _8301_ ;
wire _4641_ ;
wire _4221_ ;
wire _5846_ ;
wire _5426_ ;
wire _5006_ ;
wire _1766_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire _3912_ ;
wire _6384_ ;
wire _7589_ ;
wire _7169_ ;
wire _8950_ ;
wire _8530_ ;
wire _8110_ ;
wire _3089_ ;
wire _4870_ ;
wire _4450_ ;
wire _4030_ ;
wire _5655_ ;
wire _5235_ ;
wire _1995_ ;
wire _1575_ ;
wire _1155_ ;
wire _7801_ ;
wire _486_ ;
wire _3721_ ;
wire _3301_ ;
wire _6193_ ;
wire _4926_ ;
wire _4506_ ;
wire _7398_ ;
wire _9124_ ;
wire _5884_ ;
wire _5464_ ;
wire _5044_ ;
wire _6669_ ;
wire _6249_ ;
wire _1384_ ;
wire _7610_ ;
wire _295_ ;
wire _2589_ ;
wire _2169_ ;
wire \datapath.idinstr_20_hier0_bF$buf2  ;
wire _8815_ ;
wire _3950_ ;
wire _3530_ ;
wire _3110_ ;
wire _4735_ ;
wire _4315_ ;
wire _14_ ;
wire _2801_ ;
wire _5693_ ;
wire _5273_ ;
wire _6898_ ;
wire _6478_ ;
wire _6058_ ;
wire _1193_ ;
wire _2398_ ;
wire _8624_ ;
wire _8204_ ;
wire _4964_ ;
wire _4544_ ;
wire _4124_ ;
wire _5749_ ;
wire _5329_ ;
wire _9162_ ;
wire _1669_ ;
wire _1249_ ;
wire _2610_ ;
wire _5082_ ;
wire \datapath.idinstr_15_bF$buf21  ;
wire _3815_ ;
wire _6287_ ;
wire _8853_ ;
wire _8433_ ;
wire _8013_ ;
wire _4773_ ;
wire _4353_ ;
wire _5978_ ;
wire _5558_ ;
wire _5138_ ;
wire \datapath.idinstr_16_bF$buf30  ;
wire _52_ ;
wire _1898_ ;
wire _1478_ ;
wire _1058_ ;
wire _7704_ ;
wire _389_ ;
wire _8909_ ;
wire _3624_ ;
wire _3204_ ;
wire _6096_ ;
wire _4829_ ;
wire _4409_ ;
wire _8662_ ;
wire _8242_ ;
wire _5687__bF$buf0 ;
wire _5687__bF$buf1 ;
wire _5687__bF$buf2 ;
wire _5687__bF$buf3 ;
wire _5687__bF$buf4 ;
wire _5687__bF$buf5 ;
wire _5687__bF$buf6 ;
wire _5687__bF$buf7 ;
wire _5687__bF$buf8 ;
wire _9027_ ;
wire _4582_ ;
wire _4162_ ;
wire _601_ ;
wire _5787_ ;
wire _5367_ ;
wire _1287_ ;
wire _7933_ ;
wire _7513_ ;
wire _198_ ;
wire _8718_ ;
wire _3853_ ;
wire _3433_ ;
wire _3013_ ;
wire _4638_ ;
wire _4218_ ;
wire _8891_ ;
wire _8471_ ;
wire _8051_ ;
wire _4391_ ;
wire _830_ ;
wire _410_ ;
wire _2704_ ;
wire _5596_ ;
wire _5176_ ;
wire _90_ ;
wire _3909_ ;
wire _1096_ ;
wire _7742_ ;
wire _7322_ ;
wire _8947_ ;
wire _8527_ ;
wire _8107_ ;
wire _3662_ ;
wire _3242_ ;
wire _4867_ ;
wire _4447_ ;
wire _4027_ ;
wire _8280_ ;
wire \datapath.immediatedecoder._09_  ;
wire _9065_ ;
wire _2933_ ;
wire _2513_ ;
wire _3718_ ;
wire _7971_ ;
wire _7551_ ;
wire _7131_ ;
wire _8756_ ;
wire _8336_ ;
wire _5620__bF$buf0 ;
wire _3891_ ;
wire _5620__bF$buf1 ;
wire _3471_ ;
wire _5620__bF$buf2 ;
wire _3051_ ;
wire _5620__bF$buf3 ;
wire _5620__bF$buf4 ;
wire _4676_ ;
wire _4256_ ;
wire _6822_ ;
wire _6402_ ;
wire _7607_ ;
wire _2742_ ;
wire _2322_ ;
wire _3947_ ;
wire _3527_ ;
wire _3107_ ;
wire _8_ ;
wire _7780_ ;
wire _7360_ ;
wire _8985_ ;
wire _8565_ ;
wire _8145_ ;
wire _3280_ ;
wire _4485_ ;
wire _4065_ ;
wire _924_ ;
wire _504_ ;
wire _6631_ ;
wire _6211_ ;
wire _7836_ ;
wire _7416_ ;
wire _2971_ ;
wire _2551_ ;
wire _2131_ ;
wire _3756_ ;
wire _3336_ ;
wire \datapath.idinstr_21_bF$buf13  ;
wire _5902_ ;
wire _8794_ ;
wire _8374_ ;
wire _1822_ ;
wire _1402_ ;
wire _9159_ ;
wire _4294_ ;
wire _733_ ;
wire _313_ ;
wire _2607_ ;
wire _5499_ ;
wire _5079_ ;
wire _6860_ ;
wire _6440_ ;
wire _6020_ ;
wire \datapath.idinstr_15_bF$buf18  ;
wire \datapath.idinstr_15_hier0_bF$buf6  ;
wire \datapath.idinstr_22_bF$buf22  ;
wire _7645_ ;
wire _7225_ ;
wire _2780_ ;
wire _2360_ ;
wire _3985_ ;
wire _3565_ ;
wire _3145_ ;
wire _5711_ ;
wire _8183_ ;
wire \datapath.idinstr_16_bF$buf27  ;
wire _49_ ;
wire _6916_ ;
wire _1631_ ;
wire _1211_ ;
wire \datapath.idinstr_20_bF$buf42  ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _2836_ ;
wire \datapath.idinstr_15_bF$buf5  ;
wire _2416_ ;
wire _7874_ ;
wire _7454_ ;
wire _7034_ ;
wire [31:0] \datapath.registers.838[18]  ;
wire _8659_ ;
wire _8239_ ;
wire _3794_ ;
wire _3374_ ;
wire _4999_ ;
wire _4579_ ;
wire \datapath.idinstr_21_bF$buf51  ;
wire _4159_ ;
wire _5940_ ;
wire _5520_ ;
wire _5100_ ;
wire _6725_ ;
wire _6305_ ;
wire _1860_ ;
wire _1440_ ;
wire _1020_ ;
wire _771_ ;
wire _351_ ;
wire _2645_ ;
wire _2225_ ;
wire _7683_ ;
wire _7263_ ;
wire _8888_ ;
wire _8468_ ;
wire _8048_ ;
wire _3183_ ;
wire _1916_ ;
wire _4388_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _6954_ ;
wire _6534_ ;
wire _6114_ ;
wire _580_ ;
wire _160_ ;
wire _7739_ ;
wire _7319_ ;
wire _2874_ ;
wire _2454_ ;
wire _2034_ ;
wire _3659_ ;
wire _3239_ ;
wire _4600_ ;
wire _7492_ ;
wire _7072_ ;
wire _5805_ ;
wire _8697_ ;
wire _8277_ ;
wire _1725_ ;
wire _1305_ ;
wire _4197_ ;
wire _636_ ;
wire _216_ ;
wire _6763_ ;
wire _6343_ ;
wire _7968_ ;
wire _7548_ ;
wire _7128_ ;
wire \datapath.idinstr_24_bF$buf1  ;
wire _2683_ ;
wire _2263_ ;
wire _3888_ ;
wire _3468_ ;
wire _3048_ ;
wire _5614_ ;
wire _8086_ ;
wire [31:0] \datapath.csr._13_  ;
wire \datapath.alu.b_2_bF$buf0  ;
wire _6819_ ;
wire _1954_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire _2739_ ;
wire _2319_ ;
wire _6992_ ;
wire _6572_ ;
wire _6152_ ;
wire \controlunit.csrfile_trap_wen_bF$buf6  ;
wire _7777_ ;
wire _7357_ ;
wire _2492_ ;
wire _2072_ ;
wire \datapath.idinstr_22_bF$buf8  ;
wire _3697_ ;
wire _3277_ ;
wire _5843_ ;
wire _5423_ ;
wire _5003_ ;
wire _6628_ ;
wire _6208_ ;
wire _1763_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _2968_ ;
wire _2548_ ;
wire _2128_ ;
wire _6381_ ;
wire _7586_ ;
wire _7166_ ;
wire _3086_ ;
wire _1819_ ;
wire _5652_ ;
wire _5232_ ;
wire _6857_ ;
wire _6437_ ;
wire _6017_ ;
wire _1992_ ;
wire _1572_ ;
wire _1152_ ;
wire _483_ ;
wire \datapath.idinstr_22_bF$buf19  ;
wire _2777_ ;
wire _2357_ ;
wire _6190_ ;
wire _4923_ ;
wire _4503_ ;
wire _7395_ ;
wire _5708_ ;
wire _9121_ ;
wire _1628_ ;
wire _1208_ ;
wire _5881_ ;
wire _5461_ ;
wire _5041_ ;
wire \datapath.idinstr_20_bF$buf39  ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _6666_ ;
wire _6246_ ;
wire _1381_ ;
wire _292_ ;
wire _2586_ ;
wire _2166_ ;
wire _8812_ ;
wire _4732_ ;
wire _4312_ ;
wire \datapath.idinstr_21_bF$buf48  ;
wire _5937_ ;
wire _5517_ ;
wire _11_ ;
wire \datapath.alu.b_0_bF$buf9  ;
wire _1857_ ;
wire _1437_ ;
wire _1017_ ;
wire _5690_ ;
wire _387__bF$buf0 ;
wire _5270_ ;
wire _387__bF$buf1 ;
wire _387__bF$buf2 ;
wire _387__bF$buf3 ;
wire _387__bF$buf4 ;
wire _768_ ;
wire _348_ ;
wire _6895_ ;
wire _6475_ ;
wire _6055_ ;
wire _1190_ ;
wire _2395_ ;
wire _8621_ ;
wire _8201_ ;
wire _4961_ ;
wire _4541_ ;
wire _4121_ ;
wire [1:0] \datapath.csr.mstatus  ;
wire _5746_ ;
wire _5326_ ;
wire \controlunit.ill_op  ;
wire _1666_ ;
wire _1246_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _3812_ ;
wire _6284_ ;
wire _7489_ ;
wire _7069_ ;
wire _8850_ ;
wire _8430_ ;
wire _8010_ ;
wire _4770_ ;
wire _4350_ ;
wire \datapath.idinstr_21_hier0_bF$buf4  ;
wire _5975_ ;
wire _5555_ ;
wire _5135_ ;
wire _1895_ ;
wire _1475_ ;
wire _1055_ ;
wire _7701_ ;
wire _386_ ;
wire _8906_ ;
wire _3621_ ;
wire _3201_ ;
wire _6093_ ;
wire _4826_ ;
wire _4406_ ;
wire _7298_ ;
wire _9024_ ;
wire _5784_ ;
wire _5364_ ;
wire _6989_ ;
wire _6569_ ;
wire _6149_ ;
wire _1284_ ;
wire _7930_ ;
wire _7510_ ;
wire _195_ ;
wire _2489_ ;
wire _2069_ ;
wire _8715_ ;
wire _3850_ ;
wire _3430_ ;
wire _3010_ ;
wire _4635_ ;
wire _4215_ ;
wire _2701_ ;
wire _5593_ ;
wire _5173_ ;
wire _3906_ ;
wire _6798_ ;
wire _6378_ ;
wire _1093_ ;
wire _2298_ ;
wire _8944_ ;
wire _8524_ ;
wire _8104_ ;
wire _4864_ ;
wire _4444_ ;
wire _4024_ ;
wire _5649_ ;
wire _5229_ ;
wire _9062_ ;
wire _1989_ ;
wire _1569_ ;
wire _1149_ ;
wire _2930_ ;
wire _2510_ ;
wire _3715_ ;
wire _6187_ ;
wire _8753_ ;
wire _8333_ ;
wire _9118_ ;
wire _4673_ ;
wire _4253_ ;
wire _5878_ ;
wire _5458_ ;
wire _5038_ ;
wire _1798_ ;
wire _1378_ ;
wire _7604_ ;
wire _289_ ;
wire _8809_ ;
wire _3944_ ;
wire _3524_ ;
wire _3104_ ;
wire _5_ ;
wire _4729_ ;
wire _4309_ ;
wire _8982_ ;
wire _8562_ ;
wire _8142_ ;
wire _4482_ ;
wire _4062_ ;
wire [31:0] \datapath.muxaval  ;
wire _921_ ;
wire _501_ ;
wire _5687_ ;
wire _5267_ ;
wire [31:0] \datapath.registers.838[9]  ;
wire _1187_ ;
wire _7833_ ;
wire _7413_ ;
wire _8618_ ;
wire _3753_ ;
wire _3333_ ;
wire _4958_ ;
wire _4538_ ;
wire \datapath.idinstr_21_bF$buf10  ;
wire _4118_ ;
wire _8791_ ;
wire _8371_ ;
wire _9156_ ;
wire _4291_ ;
wire _730_ ;
wire _310_ ;
wire _2604_ ;
wire _5496_ ;
wire _5076_ ;
wire CLK_bF$buf150 ;
wire CLK_bF$buf151 ;
wire \datapath.idinstr_15_bF$buf15  ;
wire _3809_ ;
wire \datapath.idinstr_15_hier0_bF$buf3  ;
wire _7642_ ;
wire _7222_ ;
wire _8847_ ;
wire _8427_ ;
wire _8007_ ;
wire _3982_ ;
wire _3562_ ;
wire _3142_ ;
wire _4767_ ;
wire _4347_ ;
wire _8180_ ;
wire \datapath.idinstr_16_bF$buf24  ;
wire _46_ ;
wire _5477__bF$buf0 ;
wire _6913_ ;
wire _5477__bF$buf1 ;
wire _5477__bF$buf2 ;
wire _5477__bF$buf3 ;
wire _5477__bF$buf4 ;
wire _5477__bF$buf5 ;
wire _5477__bF$buf6 ;
wire _5477__bF$buf7 ;
wire _2833_ ;
wire \datapath.idinstr_15_bF$buf2  ;
wire _2413_ ;
wire _3618_ ;
wire _7871_ ;
wire _7451_ ;
wire _7031_ ;
wire _8656_ ;
wire _8236_ ;
wire _3791_ ;
wire _3371_ ;
wire _5308__bF$buf0 ;
wire _5308__bF$buf1 ;
wire _5308__bF$buf2 ;
wire _5308__bF$buf3 ;
wire _5308__bF$buf4 ;
wire _5308__bF$buf5 ;
wire _5308__bF$buf6 ;
wire _5308__bF$buf7 ;
wire \datapath.regmret  ;
wire _4996_ ;
wire _4576_ ;
wire _4156_ ;
wire _6722_ ;
wire _6302_ ;
wire _4794__bF$buf0 ;
wire _4794__bF$buf1 ;
wire _4794__bF$buf2 ;
wire _4794__bF$buf3 ;
wire _4794__bF$buf4 ;
wire _4794__bF$buf5 ;
wire _4794__bF$buf6 ;
wire _4794__bF$buf7 ;
wire _7927_ ;
wire _7507_ ;
wire _2642_ ;
wire _2222_ ;
wire \datapath.idinstr_15_bF$buf53  ;
wire _3847_ ;
wire _3427_ ;
wire _3007_ ;
wire _7680_ ;
wire _7260_ ;
wire _8885_ ;
wire _8465_ ;
wire _8045_ ;
wire _3180_ ;
wire _1913_ ;
wire _4385_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _6951_ ;
wire _6531_ ;
wire _6111_ ;
wire _7736_ ;
wire _7316_ ;
wire _2871_ ;
wire _2451_ ;
wire _2031_ ;
wire _3656_ ;
wire _3236_ ;
wire _5802_ ;
wire _8694_ ;
wire _8274_ ;
wire _5264__bF$buf0 ;
wire _5264__bF$buf1 ;
wire _5264__bF$buf2 ;
wire _5264__bF$buf3 ;
wire _5264__bF$buf4 ;
wire _1722_ ;
wire _5264__bF$buf5 ;
wire _1302_ ;
wire _5264__bF$buf6 ;
wire _5264__bF$buf7 ;
wire _9059_ ;
wire _4194_ ;
wire _633_ ;
wire _213_ ;
wire _2927_ ;
wire _2507_ ;
wire _5399_ ;
wire _6760_ ;
wire _6340_ ;
wire _4817__bF$buf0 ;
wire _4817__bF$buf1 ;
wire _4817__bF$buf2 ;
wire _4817__bF$buf3 ;
wire _4817__bF$buf4 ;
wire _7965_ ;
wire _7545_ ;
wire _7125_ ;
wire _2680_ ;
wire _2260_ ;
wire \datapath.idinstr_18_bF$buf5  ;
wire _3885_ ;
wire _3465_ ;
wire _3045_ ;
wire _5757__bF$buf0 ;
wire _5757__bF$buf1 ;
wire _5757__bF$buf2 ;
wire _5757__bF$buf3 ;
wire _5757__bF$buf4 ;
wire _5757__bF$buf5 ;
wire _5757__bF$buf6 ;
wire _5757__bF$buf7 ;
wire _5757__bF$buf8 ;
wire _5757__bF$buf9 ;
wire _5611_ ;
wire _8083_ ;
wire _6816_ ;
wire _1951_ ;
wire _1531_ ;
wire _1111_ ;
wire _862_ ;
wire _442_ ;
wire _2736_ ;
wire _2316_ ;
wire _4821__bF$buf0 ;
wire _4821__bF$buf1 ;
wire _4821__bF$buf2 ;
wire _4821__bF$buf3 ;
wire _4821__bF$buf4 ;
wire \controlunit.csrfile_trap_wen_bF$buf3  ;
wire _7774_ ;
wire _7354_ ;
wire \datapath.idinstr_22_bF$buf5  ;
wire _8979_ ;
wire _8559_ ;
wire _8139_ ;
wire _3694_ ;
wire _3274_ ;
wire _4899_ ;
wire _4479_ ;
wire _4059_ ;
wire _5840_ ;
wire _5420_ ;
wire _5000_ ;
wire _918_ ;
wire _6625_ ;
wire _6205_ ;
wire _1760_ ;
wire _1340_ ;
wire _9097_ ;
wire _671_ ;
wire _251_ ;
wire _2965_ ;
wire _2545_ ;
wire _2125_ ;
wire _7583_ ;
wire _7163_ ;
wire _8788_ ;
wire _8368_ ;
wire _3083_ ;
wire _5051__bF$buf0 ;
wire _5051__bF$buf1 ;
wire _5051__bF$buf2 ;
wire _5051__bF$buf3 ;
wire _1816_ ;
wire _5051__bF$buf4 ;
wire _5051__bF$buf5 ;
wire _4288_ ;
wire _727_ ;
wire _307_ ;
wire _6854_ ;
wire _6434_ ;
wire _6014_ ;
wire _480_ ;
wire \datapath.idinstr_22_bF$buf16  ;
wire _7639_ ;
wire _7219_ ;
wire _2774_ ;
wire _2354_ ;
wire _3979_ ;
wire _3559_ ;
wire _3139_ ;
wire _4920_ ;
wire _4500_ ;
wire _7392_ ;
wire _5705_ ;
wire _8597_ ;
wire _8177_ ;
wire _1625_ ;
wire _1205_ ;
wire _4097_ ;
wire \datapath.idinstr_20_bF$buf36  ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _6663_ ;
wire _6243_ ;
wire _7868_ ;
wire _7448_ ;
wire _7028_ ;
wire _2583_ ;
wire _2163_ ;
wire _3788_ ;
wire _3368_ ;
wire \datapath.idinstr_21_bF$buf45  ;
wire _5934_ ;
wire _5514_ ;
wire _6719_ ;
wire \datapath.alu.b_0_bF$buf6  ;
wire _1854_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _2639_ ;
wire _2219_ ;
wire _6892_ ;
wire _6472_ ;
wire _6052_ ;
wire _7677_ ;
wire _7257_ ;
wire _2392_ ;
wire _3597_ ;
wire _3177_ ;
wire _5743_ ;
wire _5323_ ;
wire _6948_ ;
wire _6528_ ;
wire _6108_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _3558__bF$buf0 ;
wire _2868_ ;
wire _3558__bF$buf1 ;
wire _2448_ ;
wire _3558__bF$buf2 ;
wire _2028_ ;
wire _3558__bF$buf3 ;
wire _3558__bF$buf4 ;
wire _6281_ ;
wire _7486_ ;
wire _7066_ ;
wire _5185__bF$buf0 ;
wire _5185__bF$buf1 ;
wire _5185__bF$buf2 ;
wire _5185__bF$buf3 ;
wire _5185__bF$buf4 ;
wire _5185__bF$buf5 ;
wire _1719_ ;
wire \datapath.idinstr_21_hier0_bF$buf1  ;
wire _5972_ ;
wire _5552_ ;
wire _5132_ ;
wire _6757_ ;
wire _6337_ ;
wire _1892_ ;
wire _1472_ ;
wire _1052_ ;
wire _383_ ;
wire _2677_ ;
wire _2257_ ;
wire _8903_ ;
wire _6090_ ;
wire \controlunit.regfile_wen  ;
wire _4823_ ;
wire _4403_ ;
wire _7295_ ;
wire _5608_ ;
wire _9021_ ;
wire _1948_ ;
wire _1528_ ;
wire _1108_ ;
wire [31:0] \datapath.csr.csr_wdata  ;
wire _5781_ ;
wire _5361_ ;
wire _859_ ;
wire _439_ ;
wire _6986_ ;
wire _6566_ ;
wire _6146_ ;
wire _1281_ ;
wire _192_ ;
wire _2486_ ;
wire _2066_ ;
wire _8712_ ;
wire _4632_ ;
wire _4212_ ;
wire _5837_ ;
wire _5417_ ;
wire _1757_ ;
wire _1337_ ;
wire _5590_ ;
wire _5170_ ;
wire _668_ ;
wire _248_ ;
wire _3903_ ;
wire _6795_ ;
wire _6375_ ;
wire _1090_ ;
wire _2295_ ;
wire _8941_ ;
wire _8521_ ;
wire _8101_ ;
wire _4861_ ;
wire _4441_ ;
wire _4021_ ;
wire _5646_ ;
wire _5226_ ;
wire _1986_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _3712_ ;
wire _6184_ ;
wire _4917_ ;
wire \datapath._34_  ;
wire _7389_ ;
wire _8750_ ;
wire _8330_ ;
wire _9115_ ;
wire _4670_ ;
wire _4250_ ;
wire _5875_ ;
wire _5455_ ;
wire _5035_ ;
wire _1795_ ;
wire _1375_ ;
wire _7601_ ;
wire _286_ ;
wire [31:0] \datapath.csr.mcause  ;
wire _8806_ ;
wire _3941_ ;
wire _3521_ ;
wire _3101_ ;
wire _2_ ;
wire _4726_ ;
wire _4306_ ;
wire _7198_ ;
wire _5684_ ;
wire _5264_ ;
wire _3132__bF$buf0 ;
wire _3132__bF$buf1 ;
wire _3132__bF$buf2 ;
wire _3132__bF$buf3 ;
wire _3132__bF$buf4 ;
wire _3132__bF$buf5 ;
wire _6889_ ;
wire _6469_ ;
wire _6049_ ;
wire _1184_ ;
wire _7830_ ;
wire _7410_ ;
wire _2389_ ;
wire _8615_ ;
wire _3750_ ;
wire _3330_ ;
wire _4955_ ;
wire _4535_ ;
wire _4115_ ;
wire _9153_ ;
wire _2601_ ;
wire _5493_ ;
wire _5073_ ;
wire CLK_bF$buf120 ;
wire CLK_bF$buf121 ;
wire CLK_bF$buf122 ;
wire CLK_bF$buf123 ;
wire CLK_bF$buf124 ;
wire CLK_bF$buf125 ;
wire \datapath.idinstr_15_bF$buf12  ;
wire CLK_bF$buf126 ;
wire CLK_bF$buf127 ;
wire CLK_bF$buf128 ;
wire _3806_ ;
wire CLK_bF$buf129 ;
wire \datapath.idinstr_15_hier0_bF$buf0  ;
wire _6698_ ;
wire _6278_ ;
wire _2198_ ;
wire _8844_ ;
wire _8424_ ;
wire _8004_ ;
wire _4805__bF$buf0 ;
wire _4805__bF$buf1 ;
wire _4805__bF$buf2 ;
wire _4805__bF$buf3 ;
wire _4805__bF$buf4 ;
wire _4764_ ;
wire _4344_ ;
wire _5969_ ;
wire _5549_ ;
wire _5129_ ;
wire \datapath.idinstr_16_bF$buf21  ;
wire _43_ ;
wire _6910_ ;
wire _1889_ ;
wire _1469_ ;
wire _1049_ ;
wire _2830_ ;
wire _2410_ ;
wire _3615_ ;
wire _6087_ ;
wire _8653_ ;
wire _8233_ ;
wire _9018_ ;
wire _4993_ ;
wire _4573_ ;
wire _4153_ ;
wire _5778_ ;
wire _5358_ ;
wire _1698_ ;
wire _1278_ ;
wire _7924_ ;
wire _7504_ ;
wire _189_ ;
wire [31:0] \datapath.registers.838[23]  ;
wire _8709_ ;
wire \datapath.idinstr_15_bF$buf50  ;
wire _3844_ ;
wire _3424_ ;
wire _3004_ ;
wire _4629_ ;
wire _4209_ ;
wire _8882_ ;
wire _8462_ ;
wire _8042_ ;
wire \datapath.idinstr_16_hier0_bF$buf5  ;
wire _1910_ ;
wire _4382_ ;
wire _821_ ;
wire _401_ ;
wire _5587_ ;
wire _5167_ ;
wire _81_ ;
wire _1087_ ;
wire _7733_ ;
wire _7313_ ;
wire _8938_ ;
wire _8518_ ;
wire _3653_ ;
wire _3233_ ;
wire _4858_ ;
wire _4438_ ;
wire _4018_ ;
wire _8691_ ;
wire _8271_ ;
wire _9056_ ;
wire _4191_ ;
wire _630_ ;
wire _210_ ;
wire _2924_ ;
wire _2504_ ;
wire _5396_ ;
wire _3709_ ;
wire _7962_ ;
wire _7542_ ;
wire _7122_ ;
wire \datapath.idinstr_18_bF$buf2  ;
wire _8747_ ;
wire _8327_ ;
wire _3882_ ;
wire _3462_ ;
wire _3042_ ;
wire [31:0] \datapath.regcsrwb  ;
wire _4667_ ;
wire _4247_ ;
wire _8080_ ;
wire _6813_ ;
wire _2733_ ;
wire _2313_ ;
wire _3938_ ;
wire _3518_ ;
wire \controlunit.csrfile_trap_wen_bF$buf0  ;
wire _7771_ ;
wire _7351_ ;
wire \datapath.idinstr_22_bF$buf2  ;
wire \datapath.idinstr_16_bF$buf9  ;
wire _8976_ ;
wire _8556_ ;
wire _8136_ ;
wire _3691_ ;
wire _3271_ ;
wire _4896_ ;
wire _4476_ ;
wire _4056_ ;
wire _915_ ;
wire _6622_ ;
wire _6202_ ;
wire _9094_ ;
wire \controlunit.mret_bF$buf4  ;
wire _7827_ ;
wire _7407_ ;
wire _2962_ ;
wire _2542_ ;
wire _2122_ ;
wire _3747_ ;
wire _3327_ ;
wire _7580_ ;
wire _7160_ ;
wire \datapath.idinstr_20_bF$buf9  ;
wire _8785_ ;
wire _8365_ ;
wire _3080_ ;
wire _1813_ ;
wire _4285_ ;
wire _724_ ;
wire _304_ ;
wire _6851_ ;
wire _6431_ ;
wire _6011_ ;
wire \datapath.idinstr_22_bF$buf13  ;
wire _7636_ ;
wire _7216_ ;
wire _2771_ ;
wire _2351_ ;
wire _3976_ ;
wire _3556_ ;
wire _3136_ ;
wire _5702_ ;
wire _8594_ ;
wire _8174_ ;
wire \datapath.idinstr_16_bF$buf18  ;
wire _6907_ ;
wire _1622_ ;
wire _1202_ ;
wire _4094_ ;
wire \datapath.idinstr_20_bF$buf33  ;
wire _953_ ;
wire _533_ ;
wire _113_ ;
wire _2827_ ;
wire _2407_ ;
wire _5299_ ;
wire _6660_ ;
wire _6240_ ;
wire _7865_ ;
wire _7445_ ;
wire _7025_ ;
wire _2580_ ;
wire _2160_ ;
wire _3785_ ;
wire _3365_ ;
wire \datapath.idinstr_21_bF$buf42  ;
wire _5931_ ;
wire _5511_ ;
wire _6716_ ;
wire \datapath.alu.b_0_bF$buf3  ;
wire _1851_ ;
wire _1431_ ;
wire _1011_ ;
wire _9188_ ;
wire _762_ ;
wire _342_ ;
wire _2636_ ;
wire _2216_ ;
wire \datapath.idinstr_15_bF$buf47  ;
wire _7674_ ;
wire _7254_ ;
wire _8879_ ;
wire _8459_ ;
wire _8039_ ;
wire _3594_ ;
wire _3174_ ;
wire _1907_ ;
wire _4799_ ;
wire _4379_ ;
wire _5740_ ;
wire _5320_ ;
wire _818_ ;
wire _78_ ;
wire _6945_ ;
wire _6525_ ;
wire _6105_ ;
wire _1660_ ;
wire _1240_ ;
wire _2251__bF$buf0 ;
wire _2251__bF$buf1 ;
wire _2251__bF$buf2 ;
wire _2251__bF$buf3 ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _2865_ ;
wire _2445_ ;
wire _2025_ ;
wire _7483_ ;
wire _7063_ ;
wire _8688_ ;
wire _8268_ ;
wire _1716_ ;
wire _4188_ ;
wire _627_ ;
wire _207_ ;
wire _6754_ ;
wire _6334_ ;
wire _380_ ;
wire _7959_ ;
wire _7539_ ;
wire _7119_ ;
wire _2674_ ;
wire _2254_ ;
wire _8900_ ;
wire _3879_ ;
wire _3459_ ;
wire _3039_ ;
wire _4820_ ;
wire _4400_ ;
wire _7292_ ;
wire _5605_ ;
wire _8497_ ;
wire _8077_ ;
wire _1945_ ;
wire _1525_ ;
wire _1105_ ;
wire _5551__bF$buf0 ;
wire _5551__bF$buf1 ;
wire _5551__bF$buf2 ;
wire _5551__bF$buf3 ;
wire _5551__bF$buf4 ;
wire _5551__bF$buf5 ;
wire _5551__bF$buf6 ;
wire _5551__bF$buf7 ;
wire _856_ ;
wire _436_ ;
wire _6983_ ;
wire _6563_ ;
wire _6143_ ;
wire \datapath.alu.b_3_bF$buf6  ;
wire _7768_ ;
wire _7348_ ;
wire _2483_ ;
wire _2063_ ;
wire _3688_ ;
wire _3268_ ;
wire _5834_ ;
wire _5414_ ;
wire _6619_ ;
wire _1754_ ;
wire _1334_ ;
wire _665_ ;
wire _245_ ;
wire _2959_ ;
wire _2539_ ;
wire _2119_ ;
wire [29:0] \datapath.csr.mepc  ;
wire _3900_ ;
wire _6792_ ;
wire _6372_ ;
wire _7997_ ;
wire _7577_ ;
wire _7157_ ;
wire _2292_ ;
wire _3497_ ;
wire _3077_ ;
wire _5643_ ;
wire _5223_ ;
wire _6848_ ;
wire _6428_ ;
wire _6008_ ;
wire _1983_ ;
wire _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _2768_ ;
wire _2348_ ;
wire _6181_ ;
wire _4914_ ;
wire _7386_ ;
wire _9112_ ;
wire _1619_ ;
wire _5872_ ;
wire _5452_ ;
wire _5032_ ;
wire _6657_ ;
wire _6237_ ;
wire _1792_ ;
wire _1372_ ;
wire CLK_hier0_bF$buf0 ;
wire CLK_hier0_bF$buf1 ;
wire CLK_hier0_bF$buf2 ;
wire CLK_hier0_bF$buf3 ;
wire CLK_hier0_bF$buf4 ;
wire CLK_hier0_bF$buf5 ;
wire CLK_hier0_bF$buf6 ;
wire CLK_hier0_bF$buf7 ;
wire CLK_hier0_bF$buf8 ;
wire CLK_hier0_bF$buf9 ;
wire _283_ ;
wire _2997_ ;
wire _2577_ ;
wire _2157_ ;
wire _8803_ ;
wire _4723_ ;
wire _4303_ ;
wire _7195_ ;
wire \datapath.idinstr_21_bF$buf39  ;
wire _5928_ ;
wire _5508_ ;
wire _1848_ ;
wire _1428_ ;
wire _1008_ ;
wire _5681_ ;
wire _5261_ ;
wire _759_ ;
wire _339_ ;
wire _6886_ ;
wire _6466_ ;
wire _6046_ ;
wire _1181_ ;
wire \datapath.idinstr_22_hier0_bF$buf5  ;
wire _2386_ ;
wire _8612_ ;
wire _4952_ ;
wire _4532_ ;
wire _4112_ ;
wire _5737_ ;
wire _5317_ ;
wire _9150_ ;
wire _1657_ ;
wire _1237_ ;
wire _5490_ ;
wire _5070_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _3803_ ;
wire _6695_ ;
wire _6275_ ;
wire _2195_ ;
wire _8841_ ;
wire _8421_ ;
wire _8001_ ;
wire _4761_ ;
wire _4341_ ;
wire _5966_ ;
wire _5546_ ;
wire _5126_ ;
wire _40_ ;
wire _1886_ ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire _3612_ ;
wire _6084_ ;
wire _4817_ ;
wire _7289_ ;
wire _8650_ ;
wire _8230_ ;
wire _9015_ ;
wire _4990_ ;
wire _4570_ ;
wire _4150_ ;
wire _5775_ ;
wire _5355_ ;
wire _1695_ ;
wire _1275_ ;
wire _7921_ ;
wire _7501_ ;
wire _186_ ;
wire _8706_ ;
wire _3841_ ;
wire _3421_ ;
wire _3001_ ;
wire _4626_ ;
wire _4206_ ;
wire _7098_ ;
wire _184__bF$buf0 ;
wire _184__bF$buf1 ;
wire _184__bF$buf2 ;
wire _184__bF$buf3 ;
wire _184__bF$buf4 ;
wire \datapath.idinstr_16_hier0_bF$buf2  ;
wire _5584_ ;
wire _5164_ ;
wire _6789_ ;
wire _6369_ ;
wire _1084_ ;
wire _7730_ ;
wire _7310_ ;
wire _2289_ ;
wire _8935_ ;
wire _8515_ ;
wire _3650_ ;
wire _3230_ ;
wire _4855_ ;
wire _4435_ ;
wire _4015_ ;
wire _9053_ ;
wire _2921_ ;
wire _2501_ ;
wire _5393_ ;
wire _3706_ ;
wire _6598_ ;
wire _6178_ ;
wire _2098_ ;
wire _8744_ ;
wire _8324_ ;
wire _9109_ ;
wire _4664_ ;
wire _4244_ ;
wire _5869_ ;
wire _5449_ ;
wire _5029_ ;
wire _6810_ ;
wire _1789_ ;
wire _1369_ ;
wire _2730_ ;
wire _2310_ ;
wire _3935_ ;
wire _3515_ ;
wire \datapath.idinstr_16_bF$buf6  ;
wire _8973_ ;
wire _8553_ ;
wire _8133_ ;
wire _4893_ ;
wire _4473_ ;
wire _4053_ ;
wire _912_ ;
wire _5678_ ;
wire _5258_ ;
wire _9091_ ;
wire \controlunit.mret_bF$buf1  ;
wire _1598_ ;
wire _1178_ ;
wire _7824_ ;
wire _7404_ ;
wire [31:0] \datapath.registers.838[13]  ;
wire _8609_ ;
wire _3744_ ;
wire _3324_ ;
wire _4949_ ;
wire \datapath.idinstr_20_bF$buf6  ;
wire _4529_ ;
wire _4109_ ;
wire _8782_ ;
wire _8362_ ;
wire _1810_ ;
wire _9147_ ;
wire _4282_ ;
wire _721_ ;
wire _301_ ;
wire _5487_ ;
wire _5067_ ;
wire _9025__bF$buf0 ;
wire _9025__bF$buf1 ;
wire _9025__bF$buf2 ;
wire \datapath.idinstr_22_bF$buf10  ;
wire _9025__bF$buf3 ;
wire _7633_ ;
wire _9025__bF$buf4 ;
wire _7213_ ;
wire _8838_ ;
wire _8418_ ;
wire _3973_ ;
wire _3553_ ;
wire _3133_ ;
wire _4758_ ;
wire _4338_ ;
wire _8591_ ;
wire _8171_ ;
wire \datapath.idinstr_16_bF$buf15  ;
wire _37_ ;
wire _6904_ ;
wire _4091_ ;
wire \datapath.idinstr_20_bF$buf30  ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _2824_ ;
wire _2404_ ;
wire _5296_ ;
wire _3609_ ;
wire _7862_ ;
wire _7442_ ;
wire _7022_ ;
wire _8647_ ;
wire _8227_ ;
wire _3782_ ;
wire _3362_ ;
wire _4987_ ;
wire _4567_ ;
wire _4147_ ;
wire _6713_ ;
wire \datapath.alu.b_0_bF$buf0  ;
wire _9185_ ;
wire _7918_ ;
wire _2633_ ;
wire _2213_ ;
wire \datapath.idinstr_15_bF$buf44  ;
wire _3838_ ;
wire _3418_ ;
wire _7671_ ;
wire _7251_ ;
wire _8876_ ;
wire _8456_ ;
wire _8036_ ;
wire _3591_ ;
wire _3171_ ;
wire _1904_ ;
wire _4796_ ;
wire _4376_ ;
wire _815_ ;
wire _75_ ;
wire _6942_ ;
wire _6522_ ;
wire _6102_ ;
wire _7727_ ;
wire _7307_ ;
wire _2862_ ;
wire _2442_ ;
wire _2022_ ;
wire _3647_ ;
wire _3227_ ;
wire _7480_ ;
wire _7060_ ;
wire _8685_ ;
wire _8265_ ;
wire _1713_ ;
wire _4185_ ;
wire _624_ ;
wire _204_ ;
wire _2918_ ;
wire _6751_ ;
wire _6331_ ;
wire _7956_ ;
wire _7536_ ;
wire _7116_ ;
wire _2671_ ;
wire _2251_ ;
wire _3876_ ;
wire _3456_ ;
wire _3036_ ;
wire _5602_ ;
wire _8494_ ;
wire _8074_ ;
wire _4827__bF$buf0 ;
wire _4827__bF$buf1 ;
wire _4827__bF$buf2 ;
wire _4827__bF$buf3 ;
wire _4827__bF$buf4 ;
wire _6807_ ;
wire _1942_ ;
wire _1522_ ;
wire _1102_ ;
wire _853_ ;
wire _433_ ;
wire _2727_ ;
wire _2307_ ;
wire _5199_ ;
wire _6980_ ;
wire _6560_ ;
wire _6140_ ;
wire \datapath.alu.b_3_bF$buf3  ;
wire _7765_ ;
wire _7345_ ;
wire _2480_ ;
wire _2060_ ;
wire [31:0] \datapath.programcounter.pc  ;
wire _3685_ ;
wire _3265_ ;
wire _5831_ ;
wire _5411_ ;
wire _909_ ;
wire _4831__bF$buf0 ;
wire _4831__bF$buf1 ;
wire _4831__bF$buf2 ;
wire _4831__bF$buf3 ;
wire _4831__bF$buf4 ;
wire _6616_ ;
wire _1751_ ;
wire _1331_ ;
wire _9088_ ;
wire _662_ ;
wire _242_ ;
wire _2956_ ;
wire _2536_ ;
wire _2116_ ;
wire _7994_ ;
wire _7574_ ;
wire _7154_ ;
wire _8779_ ;
wire _8359_ ;
wire _3494_ ;
wire _3074_ ;
wire _1807_ ;
wire _4699_ ;
wire _4279_ ;
wire _5640_ ;
wire _5220_ ;
wire _718_ ;
wire _6845_ ;
wire _6425_ ;
wire _6005_ ;
wire _1980_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _2765_ ;
wire _2345_ ;
wire _4911_ ;
wire _7383_ ;
wire _8588_ ;
wire _8168_ ;
wire _1616_ ;
wire _4088_ ;
wire \datapath.idinstr_20_bF$buf27  ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _6654_ ;
wire _6234_ ;
wire _280_ ;
wire _7859_ ;
wire _7439_ ;
wire _7019_ ;
wire _2994_ ;
wire _2574_ ;
wire _2154_ ;
wire _8800_ ;
wire _3779_ ;
wire _3359_ ;
wire _4720_ ;
wire _4300_ ;
wire _7192_ ;
wire \datapath.idinstr_21_bF$buf36  ;
wire _5925_ ;
wire _5505_ ;
wire _8397_ ;
wire _1845_ ;
wire _1425_ ;
wire _1005_ ;
wire _756_ ;
wire _336_ ;
wire _6883_ ;
wire _6463_ ;
wire _6043_ ;
wire \datapath.idinstr_22_hier0_bF$buf2  ;
wire _7668_ ;
wire _7248_ ;
wire _2383_ ;
wire _3588_ ;
wire _3168_ ;
wire _5734_ ;
wire _5314_ ;
wire _6939_ ;
wire _6519_ ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _2859_ ;
wire _2439_ ;
wire _2019_ ;
wire _3800_ ;
wire _6692_ ;
wire _6272_ ;
wire _7897_ ;
wire _7477_ ;
wire _7057_ ;
wire _2192_ ;
wire _5762__bF$buf30 ;
wire _5762__bF$buf31 ;
wire _5762__bF$buf32 ;
wire _5762__bF$buf33 ;
wire _5762__bF$buf34 ;
wire _5762__bF$buf35 ;
wire _5762__bF$buf36 ;
wire _5762__bF$buf37 ;
wire _5762__bF$buf38 ;
wire _5762__bF$buf39 ;
wire _3397_ ;
wire _5963_ ;
wire _5543_ ;
wire _5123_ ;
wire _6748_ ;
wire _6328_ ;
wire _1883_ ;
wire _1463_ ;
wire _1043_ ;
wire _794_ ;
wire _5341__bF$buf0 ;
wire _374_ ;
wire _5341__bF$buf1 ;
wire _5341__bF$buf2 ;
wire _5341__bF$buf3 ;
wire _5341__bF$buf4 ;
wire _5341__bF$buf5 ;
wire _2668_ ;
wire _2248_ ;
wire _6081_ ;
wire _4814_ ;
wire _7286_ ;
wire _9012_ ;
wire _1939_ ;
wire _1519_ ;
wire _5772_ ;
wire _5352_ ;
wire _6977_ ;
wire _6557_ ;
wire _6137_ ;
wire _1692_ ;
wire _1272_ ;
wire _183_ ;
wire _2897_ ;
wire _2477_ ;
wire _2057_ ;
wire _8703_ ;
wire _4623_ ;
wire _4203_ ;
wire _7095_ ;
wire _5828_ ;
wire _5408_ ;
wire _1748_ ;
wire _1328_ ;
wire _5581_ ;
wire _5161_ ;
wire _659_ ;
wire _239_ ;
wire [31:0] \datapath.memoryinterface.data_store  ;
wire _6786_ ;
wire _6366_ ;
wire _1081_ ;
wire _2286_ ;
wire _8932_ ;
wire _8512_ ;
wire _4852_ ;
wire _4432_ ;
wire _4012_ ;
wire _5637_ ;
wire _5217_ ;
wire _9050_ ;
wire _1977_ ;
wire _1557_ ;
wire [31:0] \datapath.registers.838[4]  ;
wire _1137_ ;
wire _7425__bF$buf40 ;
wire _7425__bF$buf41 ;
wire _7425__bF$buf42 ;
wire _7425__bF$buf43 ;
wire _7425__bF$buf44 ;
wire _7425__bF$buf45 ;
wire _7425__bF$buf46 ;
wire _7425__bF$buf47 ;
wire _5390_ ;
wire _888_ ;
wire _468_ ;
wire _3703_ ;
wire _6595_ ;
wire _6175_ ;
wire _4908_ ;
wire _2095_ ;
wire _8741_ ;
wire _8321_ ;
wire _9106_ ;
wire _4661_ ;
wire _4241_ ;
wire _5866_ ;
wire _5446_ ;
wire _5026_ ;
wire _1786_ ;
wire _1366_ ;
wire _697_ ;
wire _277_ ;
wire _3932_ ;
wire _3512_ ;
wire _4717_ ;
wire _7189_ ;
wire \datapath.idinstr_16_bF$buf3  ;
wire _8970_ ;
wire _8550_ ;
wire _8130_ ;
wire _3138__bF$buf0 ;
wire _3138__bF$buf1 ;
wire _3138__bF$buf2 ;
wire _3138__bF$buf3 ;
wire _3138__bF$buf4 ;
wire _3138__bF$buf5 ;
wire _3138__bF$buf6 ;
wire _4890_ ;
wire _4470_ ;
wire _4050_ ;
wire _0__0_bF$buf0 ;
wire _5675_ ;
wire _0__0_bF$buf1 ;
wire _5255_ ;
wire _0__0_bF$buf2 ;
wire _0__0_bF$buf3 ;
wire _0__0_bF$buf4 ;
wire _187__bF$buf0 ;
wire _187__bF$buf1 ;
wire _187__bF$buf2 ;
wire _187__bF$buf3 ;
wire _187__bF$buf4 ;
wire _1595_ ;
wire _1175_ ;
wire _7821_ ;
wire _7401_ ;
wire _8606_ ;
wire _3741_ ;
wire _3321_ ;
wire _4946_ ;
wire \datapath.idinstr_20_bF$buf3  ;
wire _4526_ ;
wire _4106_ ;
wire _9144_ ;
wire \datapath.allowcsrwrite  ;
wire _5484_ ;
wire _5064_ ;
wire _6689_ ;
wire _6269_ ;
wire _7630_ ;
wire _7210_ ;
wire _2189_ ;
wire _8835_ ;
wire _8415_ ;
wire _3970_ ;
wire _3550_ ;
wire _3130_ ;
wire _4755_ ;
wire _4335_ ;
wire \datapath.idinstr_16_bF$buf12  ;
wire _34_ ;
wire _6901_ ;
wire _2821_ ;
wire _2401_ ;
wire _5293_ ;
wire [3:0] \datapath.csr.csr_mcause  ;
wire _4815__bF$buf0 ;
wire _4815__bF$buf1 ;
wire _3606_ ;
wire _4815__bF$buf2 ;
wire _4815__bF$buf3 ;
wire _4815__bF$buf4 ;
wire _6498_ ;
wire _6078_ ;
wire _8644_ ;
wire _8224_ ;
wire _9009_ ;
wire _4984_ ;
wire _4564_ ;
wire _4144_ ;
wire _5769_ ;
wire _5349_ ;
wire _6710_ ;
wire _9182_ ;
wire _1689_ ;
wire _1269_ ;
wire _7915_ ;
wire _2630_ ;
wire _2210_ ;
wire \datapath.idinstr_15_bF$buf41  ;
wire _3835_ ;
wire _3415_ ;
wire _8873_ ;
wire _8453_ ;
wire _8033_ ;
wire _1901_ ;
wire _4793_ ;
wire _4373_ ;
wire \datapath.idinstr_23_bF$buf6  ;
wire _812_ ;
wire _5998_ ;
wire _5578_ ;
wire _5158_ ;
wire \datapath.idinstr_16_bF$buf50  ;
wire _72_ ;
wire _1498_ ;
wire _1078_ ;
wire _7724_ ;
wire _7304_ ;
wire _8929_ ;
wire _8509_ ;
wire _3644_ ;
wire _3224_ ;
wire _4849_ ;
wire _4429_ ;
wire _4009_ ;
wire _8682_ ;
wire _8262_ ;
wire _1710_ ;
wire _9047_ ;
wire _4182_ ;
wire _621_ ;
wire _201_ ;
wire _2915_ ;
wire _5387_ ;
wire _7953_ ;
wire _7533_ ;
wire _7113_ ;
wire _8738_ ;
wire _8318_ ;
wire _3873_ ;
wire _3453_ ;
wire _3033_ ;
wire _4658_ ;
wire _4238_ ;
wire _8491_ ;
wire _8071_ ;
wire _6804_ ;
wire _850_ ;
wire _430_ ;
wire _2724_ ;
wire _2304_ ;
wire _5196_ ;
wire _3929_ ;
wire _3509_ ;
wire \datapath.alu.b_3_bF$buf0  ;
wire _7762_ ;
wire _7342_ ;
wire _8967_ ;
wire _8547_ ;
wire _8127_ ;
wire _3682_ ;
wire _3262_ ;
wire _4887_ ;
wire _4467_ ;
wire _4047_ ;
wire _906_ ;
wire _6613_ ;
wire _9085_ ;
wire _7818_ ;
wire _2953_ ;
wire _2533_ ;
wire _2113_ ;
wire _3738_ ;
wire _3318_ ;
wire _7991_ ;
wire _7571_ ;
wire _7151_ ;
wire _8776_ ;
wire _8356_ ;
wire _3491_ ;
wire _3071_ ;
wire _1804_ ;
wire _4696_ ;
wire _4276_ ;
wire _715_ ;
wire _6842_ ;
wire _6422_ ;
wire _6002_ ;
wire _7627_ ;
wire _7207_ ;
wire _2762_ ;
wire _2342_ ;
wire _3967_ ;
wire _3547_ ;
wire _3127_ ;
wire _7380_ ;
wire _8585_ ;
wire _8165_ ;
wire _1613_ ;
wire _4085_ ;
wire \datapath.idinstr_20_bF$buf24  ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire _2818_ ;
wire _6651_ ;
wire _6231_ ;
wire _7856_ ;
wire _7436_ ;
wire _7016_ ;
wire _2991_ ;
wire _2571_ ;
wire _2151_ ;
wire _3776_ ;
wire _3356_ ;
wire \datapath.idinstr_21_bF$buf33  ;
wire _5922_ ;
wire _5502_ ;
wire _8394_ ;
wire _6707_ ;
wire _1842_ ;
wire _1422_ ;
wire _1002_ ;
wire _9179_ ;
wire _753_ ;
wire _333_ ;
wire _2627_ ;
wire _2207_ ;
wire _5099_ ;
wire _6880_ ;
wire _6460_ ;
wire _6040_ ;
wire \datapath.idinstr_15_bF$buf38  ;
wire _7665_ ;
wire _7245_ ;
wire _2380_ ;
wire _3585_ ;
wire _3165_ ;
wire _5731_ ;
wire _5311_ ;
wire [31:0] \datapath.registers.rega_data  ;
wire _809_ ;
wire \datapath.idinstr_16_bF$buf47  ;
wire _69_ ;
wire _6936_ ;
wire _6516_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _2856_ ;
wire _2436_ ;
wire _2016_ ;
wire _7894_ ;
wire _7474_ ;
wire _7054_ ;
wire _8679_ ;
wire _8259_ ;
wire _3394_ ;
wire _1707_ ;
wire _4599_ ;
wire _4179_ ;
wire _5960_ ;
wire _5540_ ;
wire _5120_ ;
wire _618_ ;
wire _6745_ ;
wire _6325_ ;
wire _1880_ ;
wire _1460_ ;
wire _1040_ ;
wire _791_ ;
wire _371_ ;
wire _2665_ ;
wire _2245_ ;
wire _4811_ ;
wire _7283_ ;
wire _8488_ ;
wire _8068_ ;
wire _1936_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire _6974_ ;
wire _6554_ ;
wire _6134_ ;
wire _180_ ;
wire _7759_ ;
wire _7339_ ;
wire _2894_ ;
wire _2474_ ;
wire _2054_ ;
wire _8700_ ;
wire _3679_ ;
wire _3259_ ;
wire _4620_ ;
wire _4200_ ;
wire _7092_ ;
wire _5825_ ;
wire _5405_ ;
wire _8297_ ;
wire _1745_ ;
wire _4968__bF$buf0 ;
wire _1325_ ;
wire _4968__bF$buf1 ;
wire _4968__bF$buf2 ;
wire _4968__bF$buf3 ;
wire _4968__bF$buf4 ;
wire _4968__bF$buf5 ;
wire _4968__bF$buf6 ;
wire _4968__bF$buf7 ;
wire _4968__bF$buf8 ;
wire _4968__bF$buf9 ;
wire _656_ ;
wire _236_ ;
wire _6783_ ;
wire _6363_ ;
wire _7988_ ;
wire _7568_ ;
wire _7148_ ;
wire _2283_ ;
wire _3488_ ;
wire _3068_ ;
wire _5634_ ;
wire _5214_ ;
wire _6839_ ;
wire _6419_ ;
wire _1974_ ;
wire _1554_ ;
wire _1134_ ;
wire _7425__bF$buf10 ;
wire _7425__bF$buf11 ;
wire _7425__bF$buf12 ;
wire _7425__bF$buf13 ;
wire _7425__bF$buf14 ;
wire _7425__bF$buf15 ;
wire _7425__bF$buf16 ;
wire _7425__bF$buf17 ;
wire _7425__bF$buf18 ;
wire _7425__bF$buf19 ;
wire _885_ ;
wire _465_ ;
wire _2759_ ;
wire _2339_ ;
wire _3700_ ;
wire _6592_ ;
wire _6172_ ;
wire _4905_ ;
wire _7797_ ;
wire _7377_ ;
wire _2092_ ;
wire _3297_ ;
wire _9103_ ;
wire _5863_ ;
wire _5443_ ;
wire _5023_ ;
wire _6648_ ;
wire _6228_ ;
wire _1783_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _2988_ ;
wire _2568_ ;
wire _2148_ ;
wire _4714_ ;
wire _7186_ ;
wire \datapath.idinstr_16_bF$buf0  ;
wire _5919_ ;
wire _1839_ ;
wire _1419_ ;
wire _5672_ ;
wire _5252_ ;
wire _6877_ ;
wire _6457_ ;
wire _6037_ ;
wire _1592_ ;
wire _1172_ ;
wire \datapath.idinstr_22_bF$buf39  ;
wire _2797_ ;
wire _2377_ ;
wire _8603_ ;
wire _5789__bF$buf0 ;
wire _4943_ ;
wire \datapath.idinstr_20_bF$buf0  ;
wire _5789__bF$buf1 ;
wire _4523_ ;
wire _5789__bF$buf2 ;
wire _4103_ ;
wire _5789__bF$buf3 ;
wire _5789__bF$buf4 ;
wire _5728_ ;
wire _5308_ ;
wire _9141_ ;
wire _1648_ ;
wire _1228_ ;
wire _5481_ ;
wire _5061_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _6686_ ;
wire _6266_ ;
wire _2186_ ;
wire _8832_ ;
wire _8412_ ;
wire _4752_ ;
wire _4332_ ;
wire _5957_ ;
wire _5537_ ;
wire _5117_ ;
wire _31_ ;
wire _1877_ ;
wire _1457_ ;
wire _1037_ ;
wire _5290_ ;
wire _788_ ;
wire _368_ ;
wire _3603_ ;
wire _6495_ ;
wire _6075_ ;
wire _4808_ ;
wire _8641_ ;
wire _8221_ ;
wire _9006_ ;
wire _4981_ ;
wire _4561_ ;
wire _4141_ ;
wire \datapath.idinstr_19_bF$buf3  ;
wire _5766_ ;
wire _5346_ ;
wire _1686_ ;
wire _1266_ ;
wire _7912_ ;
wire _597_ ;
wire _177_ ;
wire _3832_ ;
wire _3412_ ;
wire _5722__bF$buf0 ;
wire _5722__bF$buf1 ;
wire _5722__bF$buf2 ;
wire _5722__bF$buf3 ;
wire _5722__bF$buf4 ;
wire _4617_ ;
wire [31:0] \datapath._04_  ;
wire _7089_ ;
wire _8870_ ;
wire _8450_ ;
wire _8030_ ;
wire _4790_ ;
wire _4370_ ;
wire \datapath.idinstr_23_bF$buf3  ;
wire _5995_ ;
wire _5575_ ;
wire _5155_ ;
wire _1495_ ;
wire _1075_ ;
wire _7721_ ;
wire _7301_ ;
wire _8926_ ;
wire _8506_ ;
wire _3641_ ;
wire _3221_ ;
wire _4846_ ;
wire _4426_ ;
wire _4006_ ;
wire _9044_ ;
wire _2912_ ;
wire _5384_ ;
wire _6589_ ;
wire _6169_ ;
wire _7950_ ;
wire _7530_ ;
wire _7110_ ;
wire _2089_ ;
wire _8735_ ;
wire _8315_ ;
wire _3870_ ;
wire _3450_ ;
wire _3030_ ;
wire _4655_ ;
wire _4235_ ;
wire _6801_ ;
wire _2721_ ;
wire _2301_ ;
wire _5193_ ;
wire _3926_ ;
wire _3506_ ;
wire _6398_ ;
wire _8964_ ;
wire _8544_ ;
wire _8124_ ;
wire _4884_ ;
wire _4464_ ;
wire _4044_ ;
wire _903_ ;
wire _5669_ ;
wire _5249_ ;
wire _6610_ ;
wire _9082_ ;
wire _1589_ ;
wire _1169_ ;
wire _7815_ ;
wire _2950_ ;
wire _2530_ ;
wire _2110_ ;
wire _3735_ ;
wire _3315_ ;
wire \datapath.alu.b_1_bF$buf4  ;
wire _8773_ ;
wire _8353_ ;
wire _1801_ ;
wire _9138_ ;
wire _4693_ ;
wire _4273_ ;
wire _712_ ;
wire _5898_ ;
wire _5478_ ;
wire _5058_ ;
wire [31:0] \datapath.alu.a  ;
wire _1398_ ;
wire _5052__bF$buf0 ;
wire _5052__bF$buf1 ;
wire _5052__bF$buf2 ;
wire _5052__bF$buf3 ;
wire _5052__bF$buf4 ;
wire _7624_ ;
wire _7204_ ;
wire _8829_ ;
wire _8409_ ;
wire _3964_ ;
wire _3544_ ;
wire _3124_ ;
wire _4749_ ;
wire _4329_ ;
wire _8582_ ;
wire _8162_ ;
wire _28_ ;
wire _1610_ ;
wire _4082_ ;
wire \datapath.idinstr_20_bF$buf21  ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _2815_ ;
wire \controlunit.ebreak  ;
wire _5287_ ;
wire _7853_ ;
wire _7433_ ;
wire _7013_ ;
wire _8638_ ;
wire _8218_ ;
wire _3773_ ;
wire _3353_ ;
wire \datapath.idinstr_17_bF$buf15  ;
wire _4978_ ;
wire _4558_ ;
wire \datapath.idinstr_21_bF$buf30  ;
wire _4138_ ;
wire _8391_ ;
wire _6704_ ;
wire _9176_ ;
wire _750_ ;
wire _330_ ;
wire _7909_ ;
wire _2624_ ;
wire _2204_ ;
wire _5096_ ;
wire \datapath.idinstr_15_bF$buf35  ;
wire _3829_ ;
wire _3409_ ;
wire _7662_ ;
wire _7242_ ;
wire _8867_ ;
wire _8447_ ;
wire _8027_ ;
wire _3582_ ;
wire _3162_ ;
wire _4787_ ;
wire _4367_ ;
wire _806_ ;
wire \datapath.idinstr_16_bF$buf44  ;
wire _66_ ;
wire _6933_ ;
wire _6513_ ;
wire _7718_ ;
wire _2853_ ;
wire _2433_ ;
wire _2013_ ;
wire _3638_ ;
wire _3218_ ;
wire _7891_ ;
wire _7471_ ;
wire _7051_ ;
wire _8676_ ;
wire _8256_ ;
wire _3391_ ;
wire _1704_ ;
wire _4596_ ;
wire _4176_ ;
wire _615_ ;
wire _2909_ ;
wire _5186__bF$buf0 ;
wire _5186__bF$buf1 ;
wire _5186__bF$buf2 ;
wire _5186__bF$buf3 ;
wire _5186__bF$buf4 ;
wire _6742_ ;
wire _6322_ ;
wire _7947_ ;
wire _7527_ ;
wire _7107_ ;
wire _2662_ ;
wire _2242_ ;
wire _3867_ ;
wire _3447_ ;
wire _3027_ ;
wire _7280_ ;
wire _8485_ ;
wire _8065_ ;
wire _1933_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire _2718_ ;
wire _6971_ ;
wire _6551_ ;
wire _6131_ ;
wire _7756_ ;
wire _7336_ ;
wire _2891_ ;
wire _2471_ ;
wire _2051_ ;
wire _4837__bF$buf0 ;
wire _4837__bF$buf1 ;
wire _4837__bF$buf2 ;
wire _4837__bF$buf3 ;
wire _4837__bF$buf4 ;
wire _3676_ ;
wire _3256_ ;
wire _5822_ ;
wire _5402_ ;
wire _8294_ ;
wire [31:0] \datapath.idinstr  ;
wire _6607_ ;
wire _1742_ ;
wire _1322_ ;
wire _9079_ ;
wire _653_ ;
wire _233_ ;
wire _2947_ ;
wire _2527_ ;
wire _2107_ ;
wire _6780_ ;
wire _6360_ ;
wire _7985_ ;
wire _7565_ ;
wire _7145_ ;
wire _2280_ ;
wire _4841__bF$buf0 ;
wire _4841__bF$buf1 ;
wire _4841__bF$buf2 ;
wire _4841__bF$buf3 ;
wire _4841__bF$buf4 ;
wire _3485_ ;
wire _3065_ ;
wire _5631_ ;
wire _5211_ ;
wire _709_ ;
wire _6836_ ;
wire _6416_ ;
wire _1971_ ;
wire _1551_ ;
wire _1131_ ;
wire _882_ ;
wire _462_ ;
wire _2756_ ;
wire _2336_ ;
wire _4902_ ;
wire _7794_ ;
wire _7374_ ;
wire _8999_ ;
wire _8579_ ;
wire _8159_ ;
wire _3294_ ;
wire _9100_ ;
wire _1607_ ;
wire _4499_ ;
wire _4079_ ;
wire _5860_ ;
wire _5440_ ;
wire _5020_ ;
wire \datapath.idinstr_20_bF$buf18  ;
wire _938_ ;
wire _518_ ;
wire _6645_ ;
wire _6225_ ;
wire _1780_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _2985_ ;
wire _2565_ ;
wire _2145_ ;
wire _4711_ ;
wire _7183_ ;
wire \datapath.idinstr_21_bF$buf27  ;
wire _5916_ ;
wire _8388_ ;
wire _1836_ ;
wire _1416_ ;
wire _2047__bF$buf0 ;
wire _2047__bF$buf1 ;
wire _2047__bF$buf2 ;
wire _2047__bF$buf3 ;
wire _747_ ;
wire _327_ ;
wire _6874_ ;
wire _6454_ ;
wire _6034_ ;
wire \datapath.idinstr_22_bF$buf36  ;
wire _7659_ ;
wire _7239_ ;
wire _2794_ ;
wire _2374_ ;
wire _8600_ ;
wire _3999_ ;
wire _3579_ ;
wire _3159_ ;
wire _4940_ ;
wire _4520_ ;
wire _4100_ ;
wire _5725_ ;
wire _5305_ ;
wire _8197_ ;
wire _1645_ ;
wire _1225_ ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire _6683_ ;
wire _6263_ ;
wire _7888_ ;
wire _7468_ ;
wire _7048_ ;
wire _2183_ ;
wire _3388_ ;
wire _5954_ ;
wire _5534_ ;
wire _5114_ ;
wire _6739_ ;
wire _6319_ ;
wire _1874_ ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _2659_ ;
wire _2239_ ;
wire _3600_ ;
wire _6492_ ;
wire _6072_ ;
wire _4805_ ;
wire _7697_ ;
wire _7277_ ;
wire [31:0] \datapath.regloadwb  ;
wire _3197_ ;
wire _9003_ ;
wire \datapath.idinstr_19_bF$buf0  ;
wire _5763_ ;
wire _5343_ ;
wire _6968_ ;
wire _6548_ ;
wire _6128_ ;
wire _1683_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _2888_ ;
wire _2468_ ;
wire _2048_ ;
wire _4614_ ;
wire _7086_ ;
wire _5819_ ;
wire _1739_ ;
wire _1319_ ;
wire \datapath.idinstr_23_bF$buf0  ;
wire _5992_ ;
wire _5572_ ;
wire _5152_ ;
wire _6777_ ;
wire _6357_ ;
wire _1492_ ;
wire _1072_ ;
wire _2697_ ;
wire _2277_ ;
wire _8923_ ;
wire _8503_ ;
wire _4843_ ;
wire _4423_ ;
wire _4003_ ;
wire _5628_ ;
wire _5208_ ;
wire _9041_ ;
wire _1968_ ;
wire _1548_ ;
wire _1128_ ;
wire _5381_ ;
wire _879_ ;
wire _459_ ;
wire _6586_ ;
wire _6166_ ;
wire _2086_ ;
wire _8732_ ;
wire _8312_ ;
wire _4652_ ;
wire _4232_ ;
wire _5857_ ;
wire _5437_ ;
wire _5017_ ;
wire _1777_ ;
wire _1357_ ;
wire _5190_ ;
wire _688_ ;
wire _268_ ;
wire _3923_ ;
wire _3503_ ;
wire _6395_ ;
wire _4708_ ;
wire _8961_ ;
wire _8541_ ;
wire _8121_ ;
wire _4881_ ;
wire _4461_ ;
wire _4041_ ;
wire [3:0] \datapath.alu.funsel  ;
wire _900_ ;
wire _5666_ ;
wire _5246_ ;
wire \datapath.idinstr_17_bF$buf9  ;
wire _1586_ ;
wire _1166_ ;
wire _7812_ ;
wire _497_ ;
wire _3732_ ;
wire _3312_ ;
wire \datapath.alu.b_1_bF$buf1  ;
wire _4937_ ;
wire _4517_ ;
wire \datapath._36_  ;
wire _8770_ ;
wire _8350_ ;
wire _9135_ ;
wire _4690_ ;
wire _4270_ ;
wire \datapath.idinstr_21_bF$buf9  ;
wire _4896__bF$buf0 ;
wire _5895_ ;
wire _4896__bF$buf1 ;
wire _5475_ ;
wire _4896__bF$buf2 ;
wire _5055_ ;
wire _4896__bF$buf3 ;
wire _4896__bF$buf4 ;
wire _4896__bF$buf5 ;
wire _1395_ ;
wire _7621_ ;
wire _7201_ ;
wire _8826_ ;
wire _8406_ ;
wire _3961_ ;
wire _3541_ ;
wire _3121_ ;
wire _4746_ ;
wire _4326_ ;
wire [2:0] \datapath.aluexecptions  ;
wire _25_ ;
wire _2812_ ;
wire _5284_ ;
wire _6489_ ;
wire _6069_ ;
wire _7850_ ;
wire _7430_ ;
wire _7010_ ;
wire _8635_ ;
wire _8215_ ;
wire _3770_ ;
wire _3350_ ;
wire \datapath.idinstr_17_bF$buf12  ;
wire _4975_ ;
wire _4555_ ;
wire _4135_ ;
wire _4825__bF$buf0 ;
wire _4825__bF$buf1 ;
wire _4825__bF$buf2 ;
wire _6701_ ;
wire _4825__bF$buf3 ;
wire _4825__bF$buf4 ;
wire _9173_ ;
wire _7906_ ;
wire _2621_ ;
wire _2201_ ;
wire _5093_ ;
wire \datapath.idinstr_15_bF$buf32  ;
wire _3826_ ;
wire _3406_ ;
wire _6298_ ;
wire _8864_ ;
wire _8444_ ;
wire _8024_ ;
wire \datapath.alu.b_4_bF$buf4  ;
wire _4784_ ;
wire _4364_ ;
wire _803_ ;
wire _5989_ ;
wire _5569_ ;
wire _5149_ ;
wire \datapath.idinstr_16_bF$buf41  ;
wire _63_ ;
wire _6930_ ;
wire _6510_ ;
wire _1489_ ;
wire _1069_ ;
wire _7715_ ;
wire _2850_ ;
wire _2430_ ;
wire _2010_ ;
wire _3635_ ;
wire _3215_ ;
wire _8673_ ;
wire _8253_ ;
wire _1701_ ;
wire _9038_ ;
wire _4593_ ;
wire _4173_ ;
wire _612_ ;
wire _2906_ ;
wire _5798_ ;
wire _5378_ ;
wire [1:0] bsel ;
wire _1298_ ;
wire _7944_ ;
wire _7524_ ;
wire _7104_ ;
wire [31:0] \datapath.registers.838[25]  ;
wire _8729_ ;
wire _8309_ ;
wire _3864_ ;
wire _3444_ ;
wire _3024_ ;
wire _4649_ ;
wire _4229_ ;
wire _8482_ ;
wire CLK_bF$buf80 ;
wire _8062_ ;
wire CLK_bF$buf81 ;
wire CLK_bF$buf82 ;
wire CLK_bF$buf83 ;
wire CLK_bF$buf84 ;
wire CLK_bF$buf85 ;
wire CLK_bF$buf86 ;
wire CLK_bF$buf87 ;
wire CLK_bF$buf88 ;
wire CLK_bF$buf89 ;
wire _1930_ ;
wire _1510_ ;
wire _841_ ;
wire _421_ ;
wire _2715_ ;
wire _5187_ ;
wire _7753_ ;
wire _7333_ ;
wire _8958_ ;
wire _8538_ ;
wire _8118_ ;
wire _3673_ ;
wire _3253_ ;
wire _4878_ ;
wire _4458_ ;
wire _4038_ ;
wire _8291_ ;
wire _6604_ ;
wire _9076_ ;
wire _650_ ;
wire _230_ ;
wire _7809_ ;
wire _2944_ ;
wire _2524_ ;
wire _2104_ ;
wire _3729_ ;
wire _3309_ ;
wire _7982_ ;
wire _7562_ ;
wire _7142_ ;
wire _8767_ ;
wire _8347_ ;
wire _3482_ ;
wire _3062_ ;
wire _4687_ ;
wire _4267_ ;
wire _706_ ;
wire _6833_ ;
wire _6413_ ;
wire _7618_ ;
wire _2753_ ;
wire _2333_ ;
wire _3958_ ;
wire _3538_ ;
wire _3118_ ;
wire _7791_ ;
wire _7371_ ;
wire _8996_ ;
wire _8576_ ;
wire _8156_ ;
wire \datapath.csr._20_  ;
wire _3291_ ;
wire _1604_ ;
wire _4496_ ;
wire _4076_ ;
wire \datapath.idinstr_20_bF$buf15  ;
wire _935_ ;
wire _515_ ;
wire _2809_ ;
wire _6642_ ;
wire _6222_ ;
wire _7847_ ;
wire _7427_ ;
wire _7007_ ;
wire _2982_ ;
wire _2562_ ;
wire _2142_ ;
wire _3767_ ;
wire _3347_ ;
wire _7180_ ;
wire \datapath.idinstr_21_bF$buf24  ;
wire _5913_ ;
wire _8385_ ;
wire [2:0] \controlunit.imm_sel  ;
wire _1833_ ;
wire _1413_ ;
wire _744_ ;
wire _324_ ;
wire _2618_ ;
wire _6871_ ;
wire _6451_ ;
wire _6031_ ;
wire \datapath.idinstr_15_bF$buf29  ;
wire _5118__bF$buf0 ;
wire _5118__bF$buf1 ;
wire _5118__bF$buf2 ;
wire _5118__bF$buf3 ;
wire _5118__bF$buf4 ;
wire _5118__bF$buf5 ;
wire _5118__bF$buf6 ;
wire _5118__bF$buf7 ;
wire \datapath.idinstr_22_bF$buf33  ;
wire _7656_ ;
wire _7236_ ;
wire _2791_ ;
wire _2371_ ;
wire _3996_ ;
wire _3576_ ;
wire _3156_ ;
wire _5722_ ;
wire _5302_ ;
wire _8194_ ;
wire \datapath.idinstr_16_bF$buf38  ;
wire _6927_ ;
wire _6507_ ;
wire _1642_ ;
wire _1222_ ;
wire \datapath.idinstr_20_bF$buf53  ;
wire _973_ ;
wire _553_ ;
wire _133_ ;
wire _2847_ ;
wire _2427_ ;
wire _2007_ ;
wire _6680_ ;
wire _6260_ ;
wire _2267__bF$buf0 ;
wire _2267__bF$buf1 ;
wire _2267__bF$buf2 ;
wire _2267__bF$buf3 ;
wire _7885_ ;
wire _7465_ ;
wire _7045_ ;
wire _2180_ ;
wire _3385_ ;
wire _5951_ ;
wire _5531_ ;
wire _5111_ ;
wire _609_ ;
wire _6736_ ;
wire _6316_ ;
wire _1871_ ;
wire _1451_ ;
wire _1031_ ;
wire _782_ ;
wire _362_ ;
wire _2656_ ;
wire _2236_ ;
wire _5220__bF$buf0 ;
wire _5220__bF$buf1 ;
wire _5220__bF$buf2 ;
wire _5220__bF$buf3 ;
wire _5220__bF$buf4 ;
wire _5220__bF$buf5 ;
wire _5220__bF$buf6 ;
wire _4802_ ;
wire _5220__bF$buf7 ;
wire _7694_ ;
wire _7274_ ;
wire _8899_ ;
wire _8479_ ;
wire _8059_ ;
wire _3194_ ;
wire _1824__bF$buf0 ;
wire _1824__bF$buf1 ;
wire _1824__bF$buf2 ;
wire _1824__bF$buf3 ;
wire _1824__bF$buf4 ;
wire _1824__bF$buf5 ;
wire _9000_ ;
wire _1927_ ;
wire _1507_ ;
wire _4399_ ;
wire _5760_ ;
wire _5340_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _6965_ ;
wire _6545_ ;
wire _6125_ ;
wire _1680_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _2885_ ;
wire _2465_ ;
wire _2045_ ;
wire _4611_ ;
wire _7083_ ;
wire _5816_ ;
wire _8288_ ;
wire _3136__bF$buf0 ;
wire _3136__bF$buf1 ;
wire _3136__bF$buf2 ;
wire _3136__bF$buf3 ;
wire _3136__bF$buf4 ;
wire _3136__bF$buf5 ;
wire _3136__bF$buf6 ;
wire _3136__bF$buf7 ;
wire _1736_ ;
wire _1316_ ;
wire _647_ ;
wire _227_ ;
wire _6774_ ;
wire _6354_ ;
wire _7979_ ;
wire _7559_ ;
wire _7139_ ;
wire _2694_ ;
wire _2274_ ;
wire _8920_ ;
wire _8500_ ;
wire _3899_ ;
wire _3479_ ;
wire _3059_ ;
wire _4840_ ;
wire _4420_ ;
wire _4000_ ;
wire _5625_ ;
wire _5205_ ;
wire _8097_ ;
wire _1965_ ;
wire _1545_ ;
wire _1125_ ;
wire [31:0] \datapath.wbinstr  ;
wire _876_ ;
wire _456_ ;
wire _6583_ ;
wire _6163_ ;
wire _7788_ ;
wire _7368_ ;
wire _2083_ ;
wire _3288_ ;
wire _5854_ ;
wire _5434_ ;
wire _5014_ ;
wire [1:0] \datapath.csr._37_  ;
wire _6639_ ;
wire _6219_ ;
wire _1774_ ;
wire _1354_ ;
wire _685_ ;
wire _265_ ;
wire _2979_ ;
wire _2559_ ;
wire _2139_ ;
wire _3920_ ;
wire _3500_ ;
wire _6392_ ;
wire _4705_ ;
wire _7597_ ;
wire _7177_ ;
wire _3097_ ;
wire _5663_ ;
wire _5243_ ;
wire \datapath.idinstr_17_bF$buf6  ;
wire _6868_ ;
wire _6448_ ;
wire _6028_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _2788_ ;
wire _2368_ ;
wire [31:0] \datapath.nextpc  ;
wire _4934_ ;
wire _4514_ ;
wire _7425__hier0_bF$buf0 ;
wire _7425__hier0_bF$buf1 ;
wire _7425__hier0_bF$buf2 ;
wire _7425__hier0_bF$buf3 ;
wire _7425__hier0_bF$buf4 ;
wire _7425__hier0_bF$buf5 ;
wire _5719_ ;
wire _9132_ ;
wire _1639_ ;
wire _1219_ ;
wire \datapath.idinstr_21_bF$buf6  ;
wire _5892_ ;
wire _5472_ ;
wire _5052_ ;
wire _6677_ ;
wire _6257_ ;
wire _1392_ ;
wire _2597_ ;
wire _2177_ ;
wire _8823_ ;
wire _8403_ ;
wire _4743_ ;
wire _4323_ ;
wire _5948_ ;
wire _5528_ ;
wire _5108_ ;
wire _22_ ;
wire _1868_ ;
wire _1448_ ;
wire _1028_ ;
wire _5281_ ;
wire _779_ ;
wire _359_ ;
wire _6486_ ;
wire _6066_ ;
wire _8632_ ;
wire _8212_ ;

BUFX2 BUFX2_insert1424 (
    .A(\datapath.idinstr [16]),
    .Y(\datapath.idinstr_16_hier0_bF$buf0 )
);

BUFX2 BUFX2_insert1423 (
    .A(\datapath.idinstr [16]),
    .Y(\datapath.idinstr_16_hier0_bF$buf1 )
);

BUFX2 BUFX2_insert1422 (
    .A(\datapath.idinstr [16]),
    .Y(\datapath.idinstr_16_hier0_bF$buf2 )
);

BUFX2 BUFX2_insert1421 (
    .A(\datapath.idinstr [16]),
    .Y(\datapath.idinstr_16_hier0_bF$buf3 )
);

BUFX2 BUFX2_insert1420 (
    .A(\datapath.idinstr [16]),
    .Y(\datapath.idinstr_16_hier0_bF$buf4 )
);

BUFX2 BUFX2_insert1419 (
    .A(\datapath.idinstr [16]),
    .Y(\datapath.idinstr_16_hier0_bF$buf5 )
);

BUFX2 BUFX2_insert1418 (
    .A(\datapath.idinstr [16]),
    .Y(\datapath.idinstr_16_hier0_bF$buf6 )
);

BUFX2 BUFX2_insert1417 (
    .A(\datapath.idinstr [22]),
    .Y(\datapath.idinstr_22_hier0_bF$buf0 )
);

BUFX2 BUFX2_insert1416 (
    .A(\datapath.idinstr [22]),
    .Y(\datapath.idinstr_22_hier0_bF$buf1 )
);

BUFX2 BUFX2_insert1415 (
    .A(\datapath.idinstr [22]),
    .Y(\datapath.idinstr_22_hier0_bF$buf2 )
);

BUFX2 BUFX2_insert1414 (
    .A(\datapath.idinstr [22]),
    .Y(\datapath.idinstr_22_hier0_bF$buf3 )
);

BUFX2 BUFX2_insert1413 (
    .A(\datapath.idinstr [22]),
    .Y(\datapath.idinstr_22_hier0_bF$buf4 )
);

BUFX2 BUFX2_insert1412 (
    .A(\datapath.idinstr [22]),
    .Y(\datapath.idinstr_22_hier0_bF$buf5 )
);

BUFX2 BUFX2_insert1411 (
    .A(_7425_),
    .Y(_7425__hier0_bF$buf0)
);

BUFX2 BUFX2_insert1410 (
    .A(_7425_),
    .Y(_7425__hier0_bF$buf1)
);

BUFX2 BUFX2_insert1409 (
    .A(_7425_),
    .Y(_7425__hier0_bF$buf2)
);

BUFX2 BUFX2_insert1408 (
    .A(_7425_),
    .Y(_7425__hier0_bF$buf3)
);

BUFX2 BUFX2_insert1407 (
    .A(_7425_),
    .Y(_7425__hier0_bF$buf4)
);

BUFX2 BUFX2_insert1406 (
    .A(_7425_),
    .Y(_7425__hier0_bF$buf5)
);

CLKBUF1 CLKBUF1_insert1405 (
    .A(CLK),
    .Y(CLK_hier0_bF$buf0)
);

CLKBUF1 CLKBUF1_insert1404 (
    .A(CLK),
    .Y(CLK_hier0_bF$buf1)
);

CLKBUF1 CLKBUF1_insert1403 (
    .A(CLK),
    .Y(CLK_hier0_bF$buf2)
);

CLKBUF1 CLKBUF1_insert1402 (
    .A(CLK),
    .Y(CLK_hier0_bF$buf3)
);

CLKBUF1 CLKBUF1_insert1401 (
    .A(CLK),
    .Y(CLK_hier0_bF$buf4)
);

CLKBUF1 CLKBUF1_insert1400 (
    .A(CLK),
    .Y(CLK_hier0_bF$buf5)
);

CLKBUF1 CLKBUF1_insert1399 (
    .A(CLK),
    .Y(CLK_hier0_bF$buf6)
);

CLKBUF1 CLKBUF1_insert1398 (
    .A(CLK),
    .Y(CLK_hier0_bF$buf7)
);

CLKBUF1 CLKBUF1_insert1397 (
    .A(CLK),
    .Y(CLK_hier0_bF$buf8)
);

CLKBUF1 CLKBUF1_insert1396 (
    .A(CLK),
    .Y(CLK_hier0_bF$buf9)
);

CLKBUF1 CLKBUF1_insert1395 (
    .A(CLK),
    .Y(CLK_hier0_bF$buf10)
);

CLKBUF1 CLKBUF1_insert1394 (
    .A(CLK),
    .Y(CLK_hier0_bF$buf11)
);

BUFX2 BUFX2_insert1393 (
    .A(\datapath.idinstr [20]),
    .Y(\datapath.idinstr_20_hier0_bF$buf0 )
);

BUFX2 BUFX2_insert1392 (
    .A(\datapath.idinstr [20]),
    .Y(\datapath.idinstr_20_hier0_bF$buf1 )
);

BUFX2 BUFX2_insert1391 (
    .A(\datapath.idinstr [20]),
    .Y(\datapath.idinstr_20_hier0_bF$buf2 )
);

BUFX2 BUFX2_insert1390 (
    .A(\datapath.idinstr [20]),
    .Y(\datapath.idinstr_20_hier0_bF$buf3 )
);

BUFX2 BUFX2_insert1389 (
    .A(\datapath.idinstr [20]),
    .Y(\datapath.idinstr_20_hier0_bF$buf4 )
);

BUFX2 BUFX2_insert1388 (
    .A(\datapath.idinstr [20]),
    .Y(\datapath.idinstr_20_hier0_bF$buf5 )
);

BUFX2 BUFX2_insert1387 (
    .A(\datapath.idinstr [20]),
    .Y(\datapath.idinstr_20_hier0_bF$buf6 )
);

BUFX2 BUFX2_insert1386 (
    .A(_5762_),
    .Y(_5762__hier0_bF$buf0)
);

BUFX2 BUFX2_insert1385 (
    .A(_5762_),
    .Y(_5762__hier0_bF$buf1)
);

BUFX2 BUFX2_insert1384 (
    .A(_5762_),
    .Y(_5762__hier0_bF$buf2)
);

BUFX2 BUFX2_insert1383 (
    .A(_5762_),
    .Y(_5762__hier0_bF$buf3)
);

BUFX2 BUFX2_insert1382 (
    .A(_5762_),
    .Y(_5762__hier0_bF$buf4)
);

BUFX2 BUFX2_insert1381 (
    .A(_5762_),
    .Y(_5762__hier0_bF$buf5)
);

BUFX2 BUFX2_insert1380 (
    .A(\datapath.idinstr [15]),
    .Y(\datapath.idinstr_15_hier0_bF$buf0 )
);

BUFX2 BUFX2_insert1379 (
    .A(\datapath.idinstr [15]),
    .Y(\datapath.idinstr_15_hier0_bF$buf1 )
);

BUFX2 BUFX2_insert1378 (
    .A(\datapath.idinstr [15]),
    .Y(\datapath.idinstr_15_hier0_bF$buf2 )
);

BUFX2 BUFX2_insert1377 (
    .A(\datapath.idinstr [15]),
    .Y(\datapath.idinstr_15_hier0_bF$buf3 )
);

BUFX2 BUFX2_insert1376 (
    .A(\datapath.idinstr [15]),
    .Y(\datapath.idinstr_15_hier0_bF$buf4 )
);

BUFX2 BUFX2_insert1375 (
    .A(\datapath.idinstr [15]),
    .Y(\datapath.idinstr_15_hier0_bF$buf5 )
);

BUFX2 BUFX2_insert1374 (
    .A(\datapath.idinstr [15]),
    .Y(\datapath.idinstr_15_hier0_bF$buf6 )
);

BUFX2 BUFX2_insert1373 (
    .A(\datapath.idinstr [21]),
    .Y(\datapath.idinstr_21_hier0_bF$buf0 )
);

BUFX2 BUFX2_insert1372 (
    .A(\datapath.idinstr [21]),
    .Y(\datapath.idinstr_21_hier0_bF$buf1 )
);

BUFX2 BUFX2_insert1371 (
    .A(\datapath.idinstr [21]),
    .Y(\datapath.idinstr_21_hier0_bF$buf2 )
);

BUFX2 BUFX2_insert1370 (
    .A(\datapath.idinstr [21]),
    .Y(\datapath.idinstr_21_hier0_bF$buf3 )
);

BUFX2 BUFX2_insert1369 (
    .A(\datapath.idinstr [21]),
    .Y(\datapath.idinstr_21_hier0_bF$buf4 )
);

BUFX2 BUFX2_insert1368 (
    .A(\datapath.idinstr [21]),
    .Y(\datapath.idinstr_21_hier0_bF$buf5 )
);

BUFX2 BUFX2_insert1367 (
    .A(\datapath.idinstr [21]),
    .Y(\datapath.idinstr_21_hier0_bF$buf6 )
);

BUFX2 BUFX2_insert1366 (
    .A(_2597_),
    .Y(_2597__bF$buf0)
);

BUFX2 BUFX2_insert1365 (
    .A(_2597_),
    .Y(_2597__bF$buf1)
);

BUFX2 BUFX2_insert1364 (
    .A(_2597_),
    .Y(_2597__bF$buf2)
);

BUFX2 BUFX2_insert1363 (
    .A(_2597_),
    .Y(_2597__bF$buf3)
);

BUFX2 BUFX2_insert1362 (
    .A(_2597_),
    .Y(_2597__bF$buf4)
);

BUFX2 BUFX2_insert1361 (
    .A(_2597_),
    .Y(_2597__bF$buf5)
);

BUFX2 BUFX2_insert1360 (
    .A(_5052_),
    .Y(_5052__bF$buf0)
);

BUFX2 BUFX2_insert1359 (
    .A(_5052_),
    .Y(_5052__bF$buf1)
);

BUFX2 BUFX2_insert1358 (
    .A(_5052_),
    .Y(_5052__bF$buf2)
);

BUFX2 BUFX2_insert1357 (
    .A(_5052_),
    .Y(_5052__bF$buf3)
);

BUFX2 BUFX2_insert1356 (
    .A(_5052_),
    .Y(_5052__bF$buf4)
);

BUFX2 BUFX2_insert1355 (
    .A(_4934_),
    .Y(_4934__bF$buf0)
);

BUFX2 BUFX2_insert1354 (
    .A(_4934_),
    .Y(_4934__bF$buf1)
);

BUFX2 BUFX2_insert1353 (
    .A(_4934_),
    .Y(_4934__bF$buf2)
);

BUFX2 BUFX2_insert1352 (
    .A(_4934_),
    .Y(_4934__bF$buf3)
);

BUFX2 BUFX2_insert1351 (
    .A(_4934_),
    .Y(_4934__bF$buf4)
);

BUFX2 BUFX2_insert1350 (
    .A(_4934_),
    .Y(_4934__bF$buf5)
);

BUFX2 BUFX2_insert1349 (
    .A(_4934_),
    .Y(_4934__bF$buf6)
);

BUFX2 BUFX2_insert1348 (
    .A(_4934_),
    .Y(_4934__bF$buf7)
);

BUFX2 BUFX2_insert1347 (
    .A(_4934_),
    .Y(_4934__bF$buf8)
);

BUFX2 BUFX2_insert1346 (
    .A(_4934_),
    .Y(_4934__bF$buf9)
);

BUFX2 BUFX2_insert1345 (
    .A(_5760_),
    .Y(_5760__bF$buf0)
);

BUFX2 BUFX2_insert1344 (
    .A(_5760_),
    .Y(_5760__bF$buf1)
);

BUFX2 BUFX2_insert1343 (
    .A(_5760_),
    .Y(_5760__bF$buf2)
);

BUFX2 BUFX2_insert1342 (
    .A(_5760_),
    .Y(_5760__bF$buf3)
);

BUFX2 BUFX2_insert1341 (
    .A(_5760_),
    .Y(_5760__bF$buf4)
);

BUFX2 BUFX2_insert1340 (
    .A(_5760_),
    .Y(_5760__bF$buf5)
);

BUFX2 BUFX2_insert1339 (
    .A(_5760_),
    .Y(_5760__bF$buf6)
);

BUFX2 BUFX2_insert1338 (
    .A(_5760_),
    .Y(_5760__bF$buf7)
);

BUFX2 BUFX2_insert1337 (
    .A(_5722_),
    .Y(_5722__bF$buf0)
);

BUFX2 BUFX2_insert1336 (
    .A(_5722_),
    .Y(_5722__bF$buf1)
);

BUFX2 BUFX2_insert1335 (
    .A(_5722_),
    .Y(_5722__bF$buf2)
);

BUFX2 BUFX2_insert1334 (
    .A(_5722_),
    .Y(_5722__bF$buf3)
);

BUFX2 BUFX2_insert1333 (
    .A(_5722_),
    .Y(_5722__bF$buf4)
);

BUFX2 BUFX2_insert1332 (
    .A(_1833_),
    .Y(_1833__bF$buf0)
);

BUFX2 BUFX2_insert1331 (
    .A(_1833_),
    .Y(_1833__bF$buf1)
);

BUFX2 BUFX2_insert1330 (
    .A(_1833_),
    .Y(_1833__bF$buf2)
);

BUFX2 BUFX2_insert1329 (
    .A(_1833_),
    .Y(_1833__bF$buf3)
);

BUFX2 BUFX2_insert1328 (
    .A(_1833_),
    .Y(_1833__bF$buf4)
);

BUFX2 BUFX2_insert1327 (
    .A(_1833_),
    .Y(_1833__bF$buf5)
);

BUFX2 BUFX2_insert1326 (
    .A(_1833_),
    .Y(_1833__bF$buf6)
);

BUFX2 BUFX2_insert1325 (
    .A(_1833_),
    .Y(_1833__bF$buf7)
);

BUFX2 BUFX2_insert1324 (
    .A(_5017_),
    .Y(_5017__bF$buf0)
);

BUFX2 BUFX2_insert1323 (
    .A(_5017_),
    .Y(_5017__bF$buf1)
);

BUFX2 BUFX2_insert1322 (
    .A(_5017_),
    .Y(_5017__bF$buf2)
);

BUFX2 BUFX2_insert1321 (
    .A(_5017_),
    .Y(_5017__bF$buf3)
);

BUFX2 BUFX2_insert1320 (
    .A(_5017_),
    .Y(_5017__bF$buf4)
);

BUFX2 BUFX2_insert1319 (
    .A(_5017_),
    .Y(_5017__bF$buf5)
);

BUFX2 BUFX2_insert1318 (
    .A(_5017_),
    .Y(_5017__bF$buf6)
);

BUFX2 BUFX2_insert1317 (
    .A(_5017_),
    .Y(_5017__bF$buf7)
);

BUFX2 BUFX2_insert1316 (
    .A(_4843_),
    .Y(_4843__bF$buf0)
);

BUFX2 BUFX2_insert1315 (
    .A(_4843_),
    .Y(_4843__bF$buf1)
);

BUFX2 BUFX2_insert1314 (
    .A(_4843_),
    .Y(_4843__bF$buf2)
);

BUFX2 BUFX2_insert1313 (
    .A(_4843_),
    .Y(_4843__bF$buf3)
);

BUFX2 BUFX2_insert1312 (
    .A(_4843_),
    .Y(_4843__bF$buf4)
);

BUFX2 BUFX2_insert1311 (
    .A(_5152_),
    .Y(_5152__bF$buf0)
);

BUFX2 BUFX2_insert1310 (
    .A(_5152_),
    .Y(_5152__bF$buf1)
);

BUFX2 BUFX2_insert1309 (
    .A(_5152_),
    .Y(_5152__bF$buf2)
);

BUFX2 BUFX2_insert1308 (
    .A(_5152_),
    .Y(_5152__bF$buf3)
);

BUFX2 BUFX2_insert1307 (
    .A(_5152_),
    .Y(_5152__bF$buf4)
);

BUFX2 BUFX2_insert1306 (
    .A(_5152_),
    .Y(_5152__bF$buf5)
);

BUFX2 BUFX2_insert1305 (
    .A(_5152_),
    .Y(_5152__bF$buf6)
);

BUFX2 BUFX2_insert1304 (
    .A(_5152_),
    .Y(_5152__bF$buf7)
);

BUFX2 BUFX2_insert1303 (
    .A(_4805_),
    .Y(_4805__bF$buf0)
);

BUFX2 BUFX2_insert1302 (
    .A(_4805_),
    .Y(_4805__bF$buf1)
);

BUFX2 BUFX2_insert1301 (
    .A(_4805_),
    .Y(_4805__bF$buf2)
);

BUFX2 BUFX2_insert1300 (
    .A(_4805_),
    .Y(_4805__bF$buf3)
);

BUFX2 BUFX2_insert1299 (
    .A(_4805_),
    .Y(_4805__bF$buf4)
);

BUFX2 BUFX2_insert1298 (
    .A(_5308_),
    .Y(_5308__bF$buf0)
);

BUFX2 BUFX2_insert1297 (
    .A(_5308_),
    .Y(_5308__bF$buf1)
);

BUFX2 BUFX2_insert1296 (
    .A(_5308_),
    .Y(_5308__bF$buf2)
);

BUFX2 BUFX2_insert1295 (
    .A(_5308_),
    .Y(_5308__bF$buf3)
);

BUFX2 BUFX2_insert1294 (
    .A(_5308_),
    .Y(_5308__bF$buf4)
);

BUFX2 BUFX2_insert1293 (
    .A(_5308_),
    .Y(_5308__bF$buf5)
);

BUFX2 BUFX2_insert1292 (
    .A(_5308_),
    .Y(_5308__bF$buf6)
);

BUFX2 BUFX2_insert1291 (
    .A(_5308_),
    .Y(_5308__bF$buf7)
);

BUFX2 BUFX2_insert1290 (
    .A(_1839_),
    .Y(_1839__bF$buf0)
);

BUFX2 BUFX2_insert1289 (
    .A(_1839_),
    .Y(_1839__bF$buf1)
);

BUFX2 BUFX2_insert1288 (
    .A(_1839_),
    .Y(_1839__bF$buf2)
);

BUFX2 BUFX2_insert1287 (
    .A(_1839_),
    .Y(_1839__bF$buf3)
);

BUFX2 BUFX2_insert1286 (
    .A(_1839_),
    .Y(_1839__bF$buf4)
);

BUFX2 BUFX2_insert1285 (
    .A(_1839_),
    .Y(_1839__bF$buf5)
);

BUFX2 BUFX2_insert1284 (
    .A(_1839_),
    .Y(_1839__bF$buf6)
);

BUFX2 BUFX2_insert1283 (
    .A(_4811_),
    .Y(_4811__bF$buf0)
);

BUFX2 BUFX2_insert1282 (
    .A(_4811_),
    .Y(_4811__bF$buf1)
);

BUFX2 BUFX2_insert1281 (
    .A(_4811_),
    .Y(_4811__bF$buf2)
);

BUFX2 BUFX2_insert1280 (
    .A(_4811_),
    .Y(_4811__bF$buf3)
);

BUFX2 BUFX2_insert1279 (
    .A(_4811_),
    .Y(_4811__bF$buf4)
);

BUFX2 BUFX2_insert1278 (
    .A(_2016_),
    .Y(_2016__bF$buf0)
);

BUFX2 BUFX2_insert1277 (
    .A(_2016_),
    .Y(_2016__bF$buf1)
);

BUFX2 BUFX2_insert1276 (
    .A(_2016_),
    .Y(_2016__bF$buf2)
);

BUFX2 BUFX2_insert1275 (
    .A(_2016_),
    .Y(_2016__bF$buf3)
);

BUFX2 BUFX2_insert1274 (
    .A(_4849_),
    .Y(_4849__bF$buf0)
);

BUFX2 BUFX2_insert1273 (
    .A(_4849_),
    .Y(_4849__bF$buf1)
);

BUFX2 BUFX2_insert1272 (
    .A(_4849_),
    .Y(_4849__bF$buf2)
);

BUFX2 BUFX2_insert1271 (
    .A(_4849_),
    .Y(_4849__bF$buf3)
);

BUFX2 BUFX2_insert1270 (
    .A(_4849_),
    .Y(_4849__bF$buf4)
);

BUFX2 BUFX2_insert1269 (
    .A(_5408_),
    .Y(_5408__bF$buf0)
);

BUFX2 BUFX2_insert1268 (
    .A(_5408_),
    .Y(_5408__bF$buf1)
);

BUFX2 BUFX2_insert1267 (
    .A(_5408_),
    .Y(_5408__bF$buf2)
);

BUFX2 BUFX2_insert1266 (
    .A(_5408_),
    .Y(_5408__bF$buf3)
);

BUFX2 BUFX2_insert1265 (
    .A(_5408_),
    .Y(_5408__bF$buf4)
);

BUFX2 BUFX2_insert1264 (
    .A(_5408_),
    .Y(_5408__bF$buf5)
);

BUFX2 BUFX2_insert1263 (
    .A(_5408_),
    .Y(_5408__bF$buf6)
);

BUFX2 BUFX2_insert1262 (
    .A(_5408_),
    .Y(_5408__bF$buf7)
);

BUFX2 BUFX2_insert1261 (
    .A(_5220_),
    .Y(_5220__bF$buf0)
);

BUFX2 BUFX2_insert1260 (
    .A(_5220_),
    .Y(_5220__bF$buf1)
);

BUFX2 BUFX2_insert1259 (
    .A(_5220_),
    .Y(_5220__bF$buf2)
);

BUFX2 BUFX2_insert1258 (
    .A(_5220_),
    .Y(_5220__bF$buf3)
);

BUFX2 BUFX2_insert1257 (
    .A(_5220_),
    .Y(_5220__bF$buf4)
);

BUFX2 BUFX2_insert1256 (
    .A(_5220_),
    .Y(_5220__bF$buf5)
);

BUFX2 BUFX2_insert1255 (
    .A(_5220_),
    .Y(_5220__bF$buf6)
);

BUFX2 BUFX2_insert1254 (
    .A(_5220_),
    .Y(_5220__bF$buf7)
);

BUFX2 BUFX2_insert1253 (
    .A(_2251_),
    .Y(_2251__bF$buf0)
);

BUFX2 BUFX2_insert1252 (
    .A(_2251_),
    .Y(_2251__bF$buf1)
);

BUFX2 BUFX2_insert1251 (
    .A(_2251_),
    .Y(_2251__bF$buf2)
);

BUFX2 BUFX2_insert1250 (
    .A(_2251_),
    .Y(_2251__bF$buf3)
);

BUFX2 BUFX2_insert1249 (
    .A(\datapath.idinstr_16_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_16_bF$buf0 )
);

BUFX2 BUFX2_insert1248 (
    .A(\datapath.idinstr_16_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_16_bF$buf1 )
);

BUFX2 BUFX2_insert1247 (
    .A(\datapath.idinstr_16_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_16_bF$buf2 )
);

BUFX2 BUFX2_insert1246 (
    .A(\datapath.idinstr_16_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_16_bF$buf3 )
);

BUFX2 BUFX2_insert1245 (
    .A(\datapath.idinstr_16_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_16_bF$buf4 )
);

BUFX2 BUFX2_insert1244 (
    .A(\datapath.idinstr_16_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_16_bF$buf5 )
);

BUFX2 BUFX2_insert1243 (
    .A(\datapath.idinstr_16_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_16_bF$buf6 )
);

BUFX2 BUFX2_insert1242 (
    .A(\datapath.idinstr_16_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_16_bF$buf7 )
);

BUFX2 BUFX2_insert1241 (
    .A(\datapath.idinstr_16_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_16_bF$buf8 )
);

BUFX2 BUFX2_insert1240 (
    .A(\datapath.idinstr_16_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_16_bF$buf9 )
);

BUFX2 BUFX2_insert1239 (
    .A(\datapath.idinstr_16_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_16_bF$buf10 )
);

BUFX2 BUFX2_insert1238 (
    .A(\datapath.idinstr_16_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_16_bF$buf11 )
);

BUFX2 BUFX2_insert1237 (
    .A(\datapath.idinstr_16_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_16_bF$buf12 )
);

BUFX2 BUFX2_insert1236 (
    .A(\datapath.idinstr_16_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_16_bF$buf13 )
);

BUFX2 BUFX2_insert1235 (
    .A(\datapath.idinstr_16_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_16_bF$buf14 )
);

BUFX2 BUFX2_insert1234 (
    .A(\datapath.idinstr_16_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_16_bF$buf15 )
);

BUFX2 BUFX2_insert1233 (
    .A(\datapath.idinstr_16_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_16_bF$buf16 )
);

BUFX2 BUFX2_insert1232 (
    .A(\datapath.idinstr_16_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_16_bF$buf17 )
);

BUFX2 BUFX2_insert1231 (
    .A(\datapath.idinstr_16_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_16_bF$buf18 )
);

BUFX2 BUFX2_insert1230 (
    .A(\datapath.idinstr_16_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_16_bF$buf19 )
);

BUFX2 BUFX2_insert1229 (
    .A(\datapath.idinstr_16_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_16_bF$buf20 )
);

BUFX2 BUFX2_insert1228 (
    .A(\datapath.idinstr_16_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_16_bF$buf21 )
);

BUFX2 BUFX2_insert1227 (
    .A(\datapath.idinstr_16_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_16_bF$buf22 )
);

BUFX2 BUFX2_insert1226 (
    .A(\datapath.idinstr_16_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_16_bF$buf23 )
);

BUFX2 BUFX2_insert1225 (
    .A(\datapath.idinstr_16_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_16_bF$buf24 )
);

BUFX2 BUFX2_insert1224 (
    .A(\datapath.idinstr_16_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_16_bF$buf25 )
);

BUFX2 BUFX2_insert1223 (
    .A(\datapath.idinstr_16_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_16_bF$buf26 )
);

BUFX2 BUFX2_insert1222 (
    .A(\datapath.idinstr_16_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_16_bF$buf27 )
);

BUFX2 BUFX2_insert1221 (
    .A(\datapath.idinstr_16_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_16_bF$buf28 )
);

BUFX2 BUFX2_insert1220 (
    .A(\datapath.idinstr_16_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_16_bF$buf29 )
);

BUFX2 BUFX2_insert1219 (
    .A(\datapath.idinstr_16_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_16_bF$buf30 )
);

BUFX2 BUFX2_insert1218 (
    .A(\datapath.idinstr_16_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_16_bF$buf31 )
);

BUFX2 BUFX2_insert1217 (
    .A(\datapath.idinstr_16_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_16_bF$buf32 )
);

BUFX2 BUFX2_insert1216 (
    .A(\datapath.idinstr_16_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_16_bF$buf33 )
);

BUFX2 BUFX2_insert1215 (
    .A(\datapath.idinstr_16_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_16_bF$buf34 )
);

BUFX2 BUFX2_insert1214 (
    .A(\datapath.idinstr_16_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_16_bF$buf35 )
);

BUFX2 BUFX2_insert1213 (
    .A(\datapath.idinstr_16_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_16_bF$buf36 )
);

BUFX2 BUFX2_insert1212 (
    .A(\datapath.idinstr_16_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_16_bF$buf37 )
);

BUFX2 BUFX2_insert1211 (
    .A(\datapath.idinstr_16_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_16_bF$buf38 )
);

BUFX2 BUFX2_insert1210 (
    .A(\datapath.idinstr_16_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_16_bF$buf39 )
);

BUFX2 BUFX2_insert1209 (
    .A(\datapath.idinstr_16_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_16_bF$buf40 )
);

BUFX2 BUFX2_insert1208 (
    .A(\datapath.idinstr_16_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_16_bF$buf41 )
);

BUFX2 BUFX2_insert1207 (
    .A(\datapath.idinstr_16_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_16_bF$buf42 )
);

BUFX2 BUFX2_insert1206 (
    .A(\datapath.idinstr_16_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_16_bF$buf43 )
);

BUFX2 BUFX2_insert1205 (
    .A(\datapath.idinstr_16_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_16_bF$buf44 )
);

BUFX2 BUFX2_insert1204 (
    .A(\datapath.idinstr_16_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_16_bF$buf45 )
);

BUFX2 BUFX2_insert1203 (
    .A(\datapath.idinstr_16_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_16_bF$buf46 )
);

BUFX2 BUFX2_insert1202 (
    .A(\datapath.idinstr_16_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_16_bF$buf47 )
);

BUFX2 BUFX2_insert1201 (
    .A(\datapath.idinstr_16_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_16_bF$buf48 )
);

BUFX2 BUFX2_insert1200 (
    .A(\datapath.idinstr_16_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_16_bF$buf49 )
);

BUFX2 BUFX2_insert1199 (
    .A(\datapath.idinstr_16_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_16_bF$buf50 )
);

BUFX2 BUFX2_insert1198 (
    .A(\datapath.idinstr_16_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_16_bF$buf51 )
);

BUFX2 BUFX2_insert1197 (
    .A(_9091_),
    .Y(_9091__bF$buf0)
);

BUFX2 BUFX2_insert1196 (
    .A(_9091_),
    .Y(_9091__bF$buf1)
);

BUFX2 BUFX2_insert1195 (
    .A(_9091_),
    .Y(_9091__bF$buf2)
);

BUFX2 BUFX2_insert1194 (
    .A(_9091_),
    .Y(_9091__bF$buf3)
);

BUFX2 BUFX2_insert1193 (
    .A(_9091_),
    .Y(_9091__bF$buf4)
);

BUFX2 BUFX2_insert1192 (
    .A(_4855_),
    .Y(_4855__bF$buf0)
);

BUFX2 BUFX2_insert1191 (
    .A(_4855_),
    .Y(_4855__bF$buf1)
);

BUFX2 BUFX2_insert1190 (
    .A(_4855_),
    .Y(_4855__bF$buf2)
);

BUFX2 BUFX2_insert1189 (
    .A(_4855_),
    .Y(_4855__bF$buf3)
);

BUFX2 BUFX2_insert1188 (
    .A(_4855_),
    .Y(_4855__bF$buf4)
);

BUFX2 BUFX2_insert1187 (
    .A(_4817_),
    .Y(_4817__bF$buf0)
);

BUFX2 BUFX2_insert1186 (
    .A(_4817_),
    .Y(_4817__bF$buf1)
);

BUFX2 BUFX2_insert1185 (
    .A(_4817_),
    .Y(_4817__bF$buf2)
);

BUFX2 BUFX2_insert1184 (
    .A(_4817_),
    .Y(_4817__bF$buf3)
);

BUFX2 BUFX2_insert1183 (
    .A(_4817_),
    .Y(_4817__bF$buf4)
);

BUFX2 BUFX2_insert1182 (
    .A(_0_[0]),
    .Y(_0__0_bF$buf0)
);

BUFX2 BUFX2_insert1181 (
    .A(_0_[0]),
    .Y(_0__0_bF$buf1)
);

BUFX2 BUFX2_insert1180 (
    .A(_0_[0]),
    .Y(_0__0_bF$buf2)
);

BUFX2 BUFX2_insert1179 (
    .A(_0_[0]),
    .Y(_0__0_bF$buf3)
);

BUFX2 BUFX2_insert1178 (
    .A(_0_[0]),
    .Y(_0__0_bF$buf4)
);

BUFX2 BUFX2_insert1177 (
    .A(_4799_),
    .Y(_4799__bF$buf0)
);

BUFX2 BUFX2_insert1176 (
    .A(_4799_),
    .Y(_4799__bF$buf1)
);

BUFX2 BUFX2_insert1175 (
    .A(_4799_),
    .Y(_4799__bF$buf2)
);

BUFX2 BUFX2_insert1174 (
    .A(_4799_),
    .Y(_4799__bF$buf3)
);

BUFX2 BUFX2_insert1173 (
    .A(_4799_),
    .Y(_4799__bF$buf4)
);

BUFX2 BUFX2_insert1172 (
    .A(_4799_),
    .Y(_4799__bF$buf5)
);

BUFX2 BUFX2_insert1171 (
    .A(_4799_),
    .Y(_4799__bF$buf6)
);

BUFX2 BUFX2_insert1170 (
    .A(_4799_),
    .Y(_4799__bF$buf7)
);

BUFX2 BUFX2_insert1169 (
    .A(_3136_),
    .Y(_3136__bF$buf0)
);

BUFX2 BUFX2_insert1168 (
    .A(_3136_),
    .Y(_3136__bF$buf1)
);

BUFX2 BUFX2_insert1167 (
    .A(_3136_),
    .Y(_3136__bF$buf2)
);

BUFX2 BUFX2_insert1166 (
    .A(_3136_),
    .Y(_3136__bF$buf3)
);

BUFX2 BUFX2_insert1165 (
    .A(_3136_),
    .Y(_3136__bF$buf4)
);

BUFX2 BUFX2_insert1164 (
    .A(_3136_),
    .Y(_3136__bF$buf5)
);

BUFX2 BUFX2_insert1163 (
    .A(_3136_),
    .Y(_3136__bF$buf6)
);

BUFX2 BUFX2_insert1162 (
    .A(_3136_),
    .Y(_3136__bF$buf7)
);

BUFX2 BUFX2_insert1161 (
    .A(\datapath.idinstr [19]),
    .Y(\datapath.idinstr_19_bF$buf0 )
);

BUFX2 BUFX2_insert1160 (
    .A(\datapath.idinstr [19]),
    .Y(\datapath.idinstr_19_bF$buf1 )
);

BUFX2 BUFX2_insert1159 (
    .A(\datapath.idinstr [19]),
    .Y(\datapath.idinstr_19_bF$buf2 )
);

BUFX2 BUFX2_insert1158 (
    .A(\datapath.idinstr [19]),
    .Y(\datapath.idinstr_19_bF$buf3 )
);

BUFX2 BUFX2_insert1157 (
    .A(\datapath.idinstr [19]),
    .Y(\datapath.idinstr_19_bF$buf4 )
);

BUFX2 BUFX2_insert1156 (
    .A(\datapath.idinstr [19]),
    .Y(\datapath.idinstr_19_bF$buf5 )
);

BUFX2 BUFX2_insert1155 (
    .A(_4896_),
    .Y(_4896__bF$buf0)
);

BUFX2 BUFX2_insert1154 (
    .A(_4896_),
    .Y(_4896__bF$buf1)
);

BUFX2 BUFX2_insert1153 (
    .A(_4896_),
    .Y(_4896__bF$buf2)
);

BUFX2 BUFX2_insert1152 (
    .A(_4896_),
    .Y(_4896__bF$buf3)
);

BUFX2 BUFX2_insert1151 (
    .A(_4896_),
    .Y(_4896__bF$buf4)
);

BUFX2 BUFX2_insert1150 (
    .A(_4896_),
    .Y(_4896__bF$buf5)
);

BUFX2 BUFX2_insert1149 (
    .A(_2924_),
    .Y(_2924__bF$buf0)
);

BUFX2 BUFX2_insert1148 (
    .A(_2924_),
    .Y(_2924__bF$buf1)
);

BUFX2 BUFX2_insert1147 (
    .A(_2924_),
    .Y(_2924__bF$buf2)
);

BUFX2 BUFX2_insert1146 (
    .A(_2924_),
    .Y(_2924__bF$buf3)
);

BUFX2 BUFX2_insert1145 (
    .A(_2924_),
    .Y(_2924__bF$buf4)
);

BUFX2 BUFX2_insert1144 (
    .A(_2924_),
    .Y(_2924__bF$buf5)
);

BUFX2 BUFX2_insert1143 (
    .A(_2924_),
    .Y(_2924__bF$buf6)
);

BUFX2 BUFX2_insert1142 (
    .A(_189_),
    .Y(_189__bF$buf0)
);

BUFX2 BUFX2_insert1141 (
    .A(_189_),
    .Y(_189__bF$buf1)
);

BUFX2 BUFX2_insert1140 (
    .A(_189_),
    .Y(_189__bF$buf2)
);

BUFX2 BUFX2_insert1139 (
    .A(_189_),
    .Y(_189__bF$buf3)
);

BUFX2 BUFX2_insert1138 (
    .A(_189_),
    .Y(_189__bF$buf4)
);

BUFX2 BUFX2_insert1137 (
    .A(\datapath.idinstr_22_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_22_bF$buf0 )
);

BUFX2 BUFX2_insert1136 (
    .A(\datapath.idinstr_22_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_22_bF$buf1 )
);

BUFX2 BUFX2_insert1135 (
    .A(\datapath.idinstr_22_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_22_bF$buf2 )
);

BUFX2 BUFX2_insert1134 (
    .A(\datapath.idinstr_22_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_22_bF$buf3 )
);

BUFX2 BUFX2_insert1133 (
    .A(\datapath.idinstr_22_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_22_bF$buf4 )
);

BUFX2 BUFX2_insert1132 (
    .A(\datapath.idinstr_22_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_22_bF$buf5 )
);

BUFX2 BUFX2_insert1131 (
    .A(\datapath.idinstr_22_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_22_bF$buf6 )
);

BUFX2 BUFX2_insert1130 (
    .A(\datapath.idinstr_22_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_22_bF$buf7 )
);

BUFX2 BUFX2_insert1129 (
    .A(\datapath.idinstr_22_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_22_bF$buf8 )
);

BUFX2 BUFX2_insert1128 (
    .A(\datapath.idinstr_22_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_22_bF$buf9 )
);

BUFX2 BUFX2_insert1127 (
    .A(\datapath.idinstr_22_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_22_bF$buf10 )
);

BUFX2 BUFX2_insert1126 (
    .A(\datapath.idinstr_22_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_22_bF$buf11 )
);

BUFX2 BUFX2_insert1125 (
    .A(\datapath.idinstr_22_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_22_bF$buf12 )
);

BUFX2 BUFX2_insert1124 (
    .A(\datapath.idinstr_22_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_22_bF$buf13 )
);

BUFX2 BUFX2_insert1123 (
    .A(\datapath.idinstr_22_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_22_bF$buf14 )
);

BUFX2 BUFX2_insert1122 (
    .A(\datapath.idinstr_22_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_22_bF$buf15 )
);

BUFX2 BUFX2_insert1121 (
    .A(\datapath.idinstr_22_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_22_bF$buf16 )
);

BUFX2 BUFX2_insert1120 (
    .A(\datapath.idinstr_22_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_22_bF$buf17 )
);

BUFX2 BUFX2_insert1119 (
    .A(\datapath.idinstr_22_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_22_bF$buf18 )
);

BUFX2 BUFX2_insert1118 (
    .A(\datapath.idinstr_22_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_22_bF$buf19 )
);

BUFX2 BUFX2_insert1117 (
    .A(\datapath.idinstr_22_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_22_bF$buf20 )
);

BUFX2 BUFX2_insert1116 (
    .A(\datapath.idinstr_22_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_22_bF$buf21 )
);

BUFX2 BUFX2_insert1115 (
    .A(\datapath.idinstr_22_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_22_bF$buf22 )
);

BUFX2 BUFX2_insert1114 (
    .A(\datapath.idinstr_22_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_22_bF$buf23 )
);

BUFX2 BUFX2_insert1113 (
    .A(\datapath.idinstr_22_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_22_bF$buf24 )
);

BUFX2 BUFX2_insert1112 (
    .A(\datapath.idinstr_22_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_22_bF$buf25 )
);

BUFX2 BUFX2_insert1111 (
    .A(\datapath.idinstr_22_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_22_bF$buf26 )
);

BUFX2 BUFX2_insert1110 (
    .A(\datapath.idinstr_22_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_22_bF$buf27 )
);

BUFX2 BUFX2_insert1109 (
    .A(\datapath.idinstr_22_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_22_bF$buf28 )
);

BUFX2 BUFX2_insert1108 (
    .A(\datapath.idinstr_22_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_22_bF$buf29 )
);

BUFX2 BUFX2_insert1107 (
    .A(\datapath.idinstr_22_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_22_bF$buf30 )
);

BUFX2 BUFX2_insert1106 (
    .A(\datapath.idinstr_22_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_22_bF$buf31 )
);

BUFX2 BUFX2_insert1105 (
    .A(\datapath.idinstr_22_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_22_bF$buf32 )
);

BUFX2 BUFX2_insert1104 (
    .A(\datapath.idinstr_22_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_22_bF$buf33 )
);

BUFX2 BUFX2_insert1103 (
    .A(\datapath.idinstr_22_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_22_bF$buf34 )
);

BUFX2 BUFX2_insert1102 (
    .A(\datapath.idinstr_22_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_22_bF$buf35 )
);

BUFX2 BUFX2_insert1101 (
    .A(\datapath.idinstr_22_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_22_bF$buf36 )
);

BUFX2 BUFX2_insert1100 (
    .A(\datapath.idinstr_22_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_22_bF$buf37 )
);

BUFX2 BUFX2_insert1099 (
    .A(\datapath.idinstr_22_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_22_bF$buf38 )
);

BUFX2 BUFX2_insert1098 (
    .A(\datapath.idinstr_22_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_22_bF$buf39 )
);

BUFX2 BUFX2_insert1097 (
    .A(\datapath.idinstr_22_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_22_bF$buf40 )
);

BUFX2 BUFX2_insert1096 (
    .A(\datapath.idinstr_22_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_22_bF$buf41 )
);

BUFX2 BUFX2_insert1095 (
    .A(_5264_),
    .Y(_5264__bF$buf0)
);

BUFX2 BUFX2_insert1094 (
    .A(_5264_),
    .Y(_5264__bF$buf1)
);

BUFX2 BUFX2_insert1093 (
    .A(_5264_),
    .Y(_5264__bF$buf2)
);

BUFX2 BUFX2_insert1092 (
    .A(_5264_),
    .Y(_5264__bF$buf3)
);

BUFX2 BUFX2_insert1091 (
    .A(_5264_),
    .Y(_5264__bF$buf4)
);

BUFX2 BUFX2_insert1090 (
    .A(_5264_),
    .Y(_5264__bF$buf5)
);

BUFX2 BUFX2_insert1089 (
    .A(_5264_),
    .Y(_5264__bF$buf6)
);

BUFX2 BUFX2_insert1088 (
    .A(_5264_),
    .Y(_5264__bF$buf7)
);

BUFX2 BUFX2_insert1087 (
    .A(_286_),
    .Y(_286__bF$buf0)
);

BUFX2 BUFX2_insert1086 (
    .A(_286_),
    .Y(_286__bF$buf1)
);

BUFX2 BUFX2_insert1085 (
    .A(_286_),
    .Y(_286__bF$buf2)
);

BUFX2 BUFX2_insert1084 (
    .A(_286_),
    .Y(_286__bF$buf3)
);

BUFX2 BUFX2_insert1083 (
    .A(_286_),
    .Y(_286__bF$buf4)
);

BUFX2 BUFX2_insert1082 (
    .A(_4861_),
    .Y(_4861__bF$buf0)
);

BUFX2 BUFX2_insert1081 (
    .A(_4861_),
    .Y(_4861__bF$buf1)
);

BUFX2 BUFX2_insert1080 (
    .A(_4861_),
    .Y(_4861__bF$buf2)
);

BUFX2 BUFX2_insert1079 (
    .A(_4861_),
    .Y(_4861__bF$buf3)
);

BUFX2 BUFX2_insert1078 (
    .A(_4861_),
    .Y(_4861__bF$buf4)
);

BUFX2 BUFX2_insert1077 (
    .A(_4823_),
    .Y(_4823__bF$buf0)
);

BUFX2 BUFX2_insert1076 (
    .A(_4823_),
    .Y(_4823__bF$buf1)
);

BUFX2 BUFX2_insert1075 (
    .A(_4823_),
    .Y(_4823__bF$buf2)
);

BUFX2 BUFX2_insert1074 (
    .A(_4823_),
    .Y(_4823__bF$buf3)
);

BUFX2 BUFX2_insert1073 (
    .A(_4823_),
    .Y(_4823__bF$buf4)
);

BUFX2 BUFX2_insert1072 (
    .A(_4899_),
    .Y(_4899__bF$buf0)
);

BUFX2 BUFX2_insert1071 (
    .A(_4899_),
    .Y(_4899__bF$buf1)
);

BUFX2 BUFX2_insert1070 (
    .A(_4899_),
    .Y(_4899__bF$buf2)
);

BUFX2 BUFX2_insert1069 (
    .A(_4899_),
    .Y(_4899__bF$buf3)
);

BUFX2 BUFX2_insert1068 (
    .A(_4899_),
    .Y(_4899__bF$buf4)
);

BUFX2 BUFX2_insert1067 (
    .A(_4899_),
    .Y(_4899__bF$buf5)
);

BUFX2 BUFX2_insert1066 (
    .A(_4899_),
    .Y(_4899__bF$buf6)
);

BUFX2 BUFX2_insert1065 (
    .A(_4899_),
    .Y(_4899__bF$buf7)
);

BUFX2 BUFX2_insert1064 (
    .A(_4899_),
    .Y(_4899__bF$buf8)
);

BUFX2 BUFX2_insert1063 (
    .A(_4899_),
    .Y(_4899__bF$buf9)
);

BUFX2 BUFX2_insert1062 (
    .A(_4899_),
    .Y(_4899__bF$buf10)
);

BUFX2 BUFX2_insert1061 (
    .A(_4899_),
    .Y(_4899__bF$buf11)
);

BUFX2 BUFX2_insert1060 (
    .A(_4899_),
    .Y(_4899__bF$buf12)
);

BUFX2 BUFX2_insert1059 (
    .A(_4899_),
    .Y(_4899__bF$buf13)
);

BUFX2 BUFX2_insert1058 (
    .A(_7451_),
    .Y(_7451__bF$buf0)
);

BUFX2 BUFX2_insert1057 (
    .A(_7451_),
    .Y(_7451__bF$buf1)
);

BUFX2 BUFX2_insert1056 (
    .A(_7451_),
    .Y(_7451__bF$buf2)
);

BUFX2 BUFX2_insert1055 (
    .A(_7451_),
    .Y(_7451__bF$buf3)
);

BUFX2 BUFX2_insert1054 (
    .A(_7451_),
    .Y(_7451__bF$buf4)
);

BUFX2 BUFX2_insert1053 (
    .A(_5687_),
    .Y(_5687__bF$buf0)
);

BUFX2 BUFX2_insert1052 (
    .A(_5687_),
    .Y(_5687__bF$buf1)
);

BUFX2 BUFX2_insert1051 (
    .A(_5687_),
    .Y(_5687__bF$buf2)
);

BUFX2 BUFX2_insert1050 (
    .A(_5687_),
    .Y(_5687__bF$buf3)
);

BUFX2 BUFX2_insert1049 (
    .A(_5687_),
    .Y(_5687__bF$buf4)
);

BUFX2 BUFX2_insert1048 (
    .A(_5687_),
    .Y(_5687__bF$buf5)
);

BUFX2 BUFX2_insert1047 (
    .A(_5687_),
    .Y(_5687__bF$buf6)
);

BUFX2 BUFX2_insert1046 (
    .A(_5687_),
    .Y(_5687__bF$buf7)
);

BUFX2 BUFX2_insert1045 (
    .A(_5687_),
    .Y(_5687__bF$buf8)
);

BUFX2 BUFX2_insert1044 (
    .A(_386_),
    .Y(_386__bF$buf0)
);

BUFX2 BUFX2_insert1043 (
    .A(_386_),
    .Y(_386__bF$buf1)
);

BUFX2 BUFX2_insert1042 (
    .A(_386_),
    .Y(_386__bF$buf2)
);

BUFX2 BUFX2_insert1041 (
    .A(_386_),
    .Y(_386__bF$buf3)
);

BUFX2 BUFX2_insert1040 (
    .A(_386_),
    .Y(_386__bF$buf4)
);

BUFX2 BUFX2_insert1039 (
    .A(_4829_),
    .Y(_4829__bF$buf0)
);

BUFX2 BUFX2_insert1038 (
    .A(_4829_),
    .Y(_4829__bF$buf1)
);

BUFX2 BUFX2_insert1037 (
    .A(_4829_),
    .Y(_4829__bF$buf2)
);

BUFX2 BUFX2_insert1036 (
    .A(_4829_),
    .Y(_4829__bF$buf3)
);

BUFX2 BUFX2_insert1035 (
    .A(_4829_),
    .Y(_4829__bF$buf4)
);

BUFX2 BUFX2_insert1034 (
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf0 )
);

BUFX2 BUFX2_insert1033 (
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf1 )
);

BUFX2 BUFX2_insert1032 (
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf2 )
);

BUFX2 BUFX2_insert1031 (
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf3 )
);

BUFX2 BUFX2_insert1030 (
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf4 )
);

BUFX2 BUFX2_insert1029 (
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf5 )
);

BUFX2 BUFX2_insert1028 (
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf6 )
);

BUFX2 BUFX2_insert1027 (
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf7 )
);

BUFX2 BUFX2_insert1026 (
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf8 )
);

BUFX2 BUFX2_insert1025 (
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf9 )
);

BUFX2 BUFX2_insert1024 (
    .A(_2783_),
    .Y(_2783__bF$buf0)
);

BUFX2 BUFX2_insert1023 (
    .A(_2783_),
    .Y(_2783__bF$buf1)
);

BUFX2 BUFX2_insert1022 (
    .A(_2783_),
    .Y(_2783__bF$buf2)
);

BUFX2 BUFX2_insert1021 (
    .A(_2783_),
    .Y(_2783__bF$buf3)
);

BUFX2 BUFX2_insert1020 (
    .A(_2783_),
    .Y(_2783__bF$buf4)
);

BUFX2 BUFX2_insert1019 (
    .A(_7419_),
    .Y(_7419__bF$buf0)
);

BUFX2 BUFX2_insert1018 (
    .A(_7419_),
    .Y(_7419__bF$buf1)
);

BUFX2 BUFX2_insert1017 (
    .A(_7419_),
    .Y(_7419__bF$buf2)
);

BUFX2 BUFX2_insert1016 (
    .A(_7419_),
    .Y(_7419__bF$buf3)
);

BUFX2 BUFX2_insert1015 (
    .A(_7419_),
    .Y(_7419__bF$buf4)
);

BUFX2 BUFX2_insert1014 (
    .A(_7419_),
    .Y(_7419__bF$buf5)
);

BUFX2 BUFX2_insert1013 (
    .A(_7419_),
    .Y(_7419__bF$buf6)
);

BUFX2 BUFX2_insert1012 (
    .A(_7419_),
    .Y(_7419__bF$buf7)
);

BUFX2 BUFX2_insert1011 (
    .A(_7419_),
    .Y(_7419__bF$buf8)
);

BUFX2 BUFX2_insert1010 (
    .A(_7419_),
    .Y(_7419__bF$buf9)
);

BUFX2 BUFX2_insert1009 (
    .A(_5620_),
    .Y(_5620__bF$buf0)
);

BUFX2 BUFX2_insert1008 (
    .A(_5620_),
    .Y(_5620__bF$buf1)
);

BUFX2 BUFX2_insert1007 (
    .A(_5620_),
    .Y(_5620__bF$buf2)
);

BUFX2 BUFX2_insert1006 (
    .A(_5620_),
    .Y(_5620__bF$buf3)
);

BUFX2 BUFX2_insert1005 (
    .A(_5620_),
    .Y(_5620__bF$buf4)
);

BUFX2 BUFX2_insert1004 (
    .A(\datapath.alu.b [3]),
    .Y(\datapath.alu.b_3_bF$buf0 )
);

BUFX2 BUFX2_insert1003 (
    .A(\datapath.alu.b [3]),
    .Y(\datapath.alu.b_3_bF$buf1 )
);

BUFX2 BUFX2_insert1002 (
    .A(\datapath.alu.b [3]),
    .Y(\datapath.alu.b_3_bF$buf2 )
);

BUFX2 BUFX2_insert1001 (
    .A(\datapath.alu.b [3]),
    .Y(\datapath.alu.b_3_bF$buf3 )
);

BUFX2 BUFX2_insert1000 (
    .A(\datapath.alu.b [3]),
    .Y(\datapath.alu.b_3_bF$buf4 )
);

BUFX2 BUFX2_insert999 (
    .A(\datapath.alu.b [3]),
    .Y(\datapath.alu.b_3_bF$buf5 )
);

BUFX2 BUFX2_insert998 (
    .A(\datapath.alu.b [3]),
    .Y(\datapath.alu.b_3_bF$buf6 )
);

BUFX2 BUFX2_insert997 (
    .A(\datapath.alu.b [3]),
    .Y(\datapath.alu.b_3_bF$buf7 )
);

BUFX2 BUFX2_insert996 (
    .A(_5085_),
    .Y(_5085__bF$buf0)
);

BUFX2 BUFX2_insert995 (
    .A(_5085_),
    .Y(_5085__bF$buf1)
);

BUFX2 BUFX2_insert994 (
    .A(_5085_),
    .Y(_5085__bF$buf2)
);

BUFX2 BUFX2_insert993 (
    .A(_5085_),
    .Y(_5085__bF$buf3)
);

BUFX2 BUFX2_insert992 (
    .A(_5085_),
    .Y(_5085__bF$buf4)
);

BUFX2 BUFX2_insert991 (
    .A(_5085_),
    .Y(_5085__bF$buf5)
);

BUFX2 BUFX2_insert990 (
    .A(_5085_),
    .Y(_5085__bF$buf6)
);

BUFX2 BUFX2_insert989 (
    .A(_5085_),
    .Y(_5085__bF$buf7)
);

BUFX2 BUFX2_insert988 (
    .A(_7422_),
    .Y(_7422__bF$buf0)
);

BUFX2 BUFX2_insert987 (
    .A(_7422_),
    .Y(_7422__bF$buf1)
);

BUFX2 BUFX2_insert986 (
    .A(_7422_),
    .Y(_7422__bF$buf2)
);

BUFX2 BUFX2_insert985 (
    .A(_7422_),
    .Y(_7422__bF$buf3)
);

BUFX2 BUFX2_insert984 (
    .A(_7422_),
    .Y(_7422__bF$buf4)
);

BUFX2 BUFX2_insert983 (
    .A(_4835_),
    .Y(_4835__bF$buf0)
);

BUFX2 BUFX2_insert982 (
    .A(_4835_),
    .Y(_4835__bF$buf1)
);

BUFX2 BUFX2_insert981 (
    .A(_4835_),
    .Y(_4835__bF$buf2)
);

BUFX2 BUFX2_insert980 (
    .A(_4835_),
    .Y(_4835__bF$buf3)
);

BUFX2 BUFX2_insert979 (
    .A(_4835_),
    .Y(_4835__bF$buf4)
);

BUFX2 BUFX2_insert978 (
    .A(_5755_),
    .Y(_5755__bF$buf0)
);

BUFX2 BUFX2_insert977 (
    .A(_5755_),
    .Y(_5755__bF$buf1)
);

BUFX2 BUFX2_insert976 (
    .A(_5755_),
    .Y(_5755__bF$buf2)
);

BUFX2 BUFX2_insert975 (
    .A(_5755_),
    .Y(_5755__bF$buf3)
);

BUFX2 BUFX2_insert974 (
    .A(_5755_),
    .Y(_5755__bF$buf4)
);

BUFX2 BUFX2_insert973 (
    .A(_7425__hier0_bF$buf5),
    .Y(_7425__bF$buf0)
);

BUFX2 BUFX2_insert972 (
    .A(_7425__hier0_bF$buf4),
    .Y(_7425__bF$buf1)
);

BUFX2 BUFX2_insert971 (
    .A(_7425__hier0_bF$buf3),
    .Y(_7425__bF$buf2)
);

BUFX2 BUFX2_insert970 (
    .A(_7425__hier0_bF$buf2),
    .Y(_7425__bF$buf3)
);

BUFX2 BUFX2_insert969 (
    .A(_7425__hier0_bF$buf1),
    .Y(_7425__bF$buf4)
);

BUFX2 BUFX2_insert968 (
    .A(_7425__hier0_bF$buf0),
    .Y(_7425__bF$buf5)
);

BUFX2 BUFX2_insert967 (
    .A(_7425__hier0_bF$buf5),
    .Y(_7425__bF$buf6)
);

BUFX2 BUFX2_insert966 (
    .A(_7425__hier0_bF$buf4),
    .Y(_7425__bF$buf7)
);

BUFX2 BUFX2_insert965 (
    .A(_7425__hier0_bF$buf3),
    .Y(_7425__bF$buf8)
);

BUFX2 BUFX2_insert964 (
    .A(_7425__hier0_bF$buf2),
    .Y(_7425__bF$buf9)
);

BUFX2 BUFX2_insert963 (
    .A(_7425__hier0_bF$buf1),
    .Y(_7425__bF$buf10)
);

BUFX2 BUFX2_insert962 (
    .A(_7425__hier0_bF$buf0),
    .Y(_7425__bF$buf11)
);

BUFX2 BUFX2_insert961 (
    .A(_7425__hier0_bF$buf5),
    .Y(_7425__bF$buf12)
);

BUFX2 BUFX2_insert960 (
    .A(_7425__hier0_bF$buf4),
    .Y(_7425__bF$buf13)
);

BUFX2 BUFX2_insert959 (
    .A(_7425__hier0_bF$buf3),
    .Y(_7425__bF$buf14)
);

BUFX2 BUFX2_insert958 (
    .A(_7425__hier0_bF$buf2),
    .Y(_7425__bF$buf15)
);

BUFX2 BUFX2_insert957 (
    .A(_7425__hier0_bF$buf1),
    .Y(_7425__bF$buf16)
);

BUFX2 BUFX2_insert956 (
    .A(_7425__hier0_bF$buf0),
    .Y(_7425__bF$buf17)
);

BUFX2 BUFX2_insert955 (
    .A(_7425__hier0_bF$buf5),
    .Y(_7425__bF$buf18)
);

BUFX2 BUFX2_insert954 (
    .A(_7425__hier0_bF$buf4),
    .Y(_7425__bF$buf19)
);

BUFX2 BUFX2_insert953 (
    .A(_7425__hier0_bF$buf3),
    .Y(_7425__bF$buf20)
);

BUFX2 BUFX2_insert952 (
    .A(_7425__hier0_bF$buf2),
    .Y(_7425__bF$buf21)
);

BUFX2 BUFX2_insert951 (
    .A(_7425__hier0_bF$buf1),
    .Y(_7425__bF$buf22)
);

BUFX2 BUFX2_insert950 (
    .A(_7425__hier0_bF$buf0),
    .Y(_7425__bF$buf23)
);

BUFX2 BUFX2_insert949 (
    .A(_7425__hier0_bF$buf5),
    .Y(_7425__bF$buf24)
);

BUFX2 BUFX2_insert948 (
    .A(_7425__hier0_bF$buf4),
    .Y(_7425__bF$buf25)
);

BUFX2 BUFX2_insert947 (
    .A(_7425__hier0_bF$buf3),
    .Y(_7425__bF$buf26)
);

BUFX2 BUFX2_insert946 (
    .A(_7425__hier0_bF$buf2),
    .Y(_7425__bF$buf27)
);

BUFX2 BUFX2_insert945 (
    .A(_7425__hier0_bF$buf1),
    .Y(_7425__bF$buf28)
);

BUFX2 BUFX2_insert944 (
    .A(_7425__hier0_bF$buf0),
    .Y(_7425__bF$buf29)
);

BUFX2 BUFX2_insert943 (
    .A(_7425__hier0_bF$buf5),
    .Y(_7425__bF$buf30)
);

BUFX2 BUFX2_insert942 (
    .A(_7425__hier0_bF$buf4),
    .Y(_7425__bF$buf31)
);

BUFX2 BUFX2_insert941 (
    .A(_7425__hier0_bF$buf3),
    .Y(_7425__bF$buf32)
);

BUFX2 BUFX2_insert940 (
    .A(_7425__hier0_bF$buf2),
    .Y(_7425__bF$buf33)
);

BUFX2 BUFX2_insert939 (
    .A(_7425__hier0_bF$buf1),
    .Y(_7425__bF$buf34)
);

BUFX2 BUFX2_insert938 (
    .A(_7425__hier0_bF$buf0),
    .Y(_7425__bF$buf35)
);

BUFX2 BUFX2_insert937 (
    .A(_7425__hier0_bF$buf5),
    .Y(_7425__bF$buf36)
);

BUFX2 BUFX2_insert936 (
    .A(_7425__hier0_bF$buf4),
    .Y(_7425__bF$buf37)
);

BUFX2 BUFX2_insert935 (
    .A(_7425__hier0_bF$buf3),
    .Y(_7425__bF$buf38)
);

BUFX2 BUFX2_insert934 (
    .A(_7425__hier0_bF$buf2),
    .Y(_7425__bF$buf39)
);

BUFX2 BUFX2_insert933 (
    .A(_7425__hier0_bF$buf1),
    .Y(_7425__bF$buf40)
);

BUFX2 BUFX2_insert932 (
    .A(_7425__hier0_bF$buf0),
    .Y(_7425__bF$buf41)
);

BUFX2 BUFX2_insert931 (
    .A(_7425__hier0_bF$buf5),
    .Y(_7425__bF$buf42)
);

BUFX2 BUFX2_insert930 (
    .A(_7425__hier0_bF$buf4),
    .Y(_7425__bF$buf43)
);

BUFX2 BUFX2_insert929 (
    .A(_7425__hier0_bF$buf3),
    .Y(_7425__bF$buf44)
);

BUFX2 BUFX2_insert928 (
    .A(_7425__hier0_bF$buf2),
    .Y(_7425__bF$buf45)
);

BUFX2 BUFX2_insert927 (
    .A(_7425__hier0_bF$buf1),
    .Y(_7425__bF$buf46)
);

BUFX2 BUFX2_insert926 (
    .A(_7425__hier0_bF$buf0),
    .Y(_7425__bF$buf47)
);

BUFX2 BUFX2_insert925 (
    .A(_5185_),
    .Y(_5185__bF$buf0)
);

BUFX2 BUFX2_insert924 (
    .A(_5185_),
    .Y(_5185__bF$buf1)
);

BUFX2 BUFX2_insert923 (
    .A(_5185_),
    .Y(_5185__bF$buf2)
);

BUFX2 BUFX2_insert922 (
    .A(_5185_),
    .Y(_5185__bF$buf3)
);

BUFX2 BUFX2_insert921 (
    .A(_5185_),
    .Y(_5185__bF$buf4)
);

BUFX2 BUFX2_insert920 (
    .A(_5185_),
    .Y(_5185__bF$buf5)
);

BUFX2 BUFX2_insert919 (
    .A(_4935_),
    .Y(_4935__bF$buf0)
);

BUFX2 BUFX2_insert918 (
    .A(_4935_),
    .Y(_4935__bF$buf1)
);

BUFX2 BUFX2_insert917 (
    .A(_4935_),
    .Y(_4935__bF$buf2)
);

BUFX2 BUFX2_insert916 (
    .A(_4935_),
    .Y(_4935__bF$buf3)
);

BUFX2 BUFX2_insert915 (
    .A(_4935_),
    .Y(_4935__bF$buf4)
);

BUFX2 BUFX2_insert914 (
    .A(_4935_),
    .Y(_4935__bF$buf5)
);

BUFX2 BUFX2_insert913 (
    .A(_4935_),
    .Y(_4935__bF$buf6)
);

BUFX2 BUFX2_insert912 (
    .A(_4935_),
    .Y(_4935__bF$buf7)
);

CLKBUF1 CLKBUF1_insert911 (
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf0)
);

CLKBUF1 CLKBUF1_insert910 (
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf1)
);

CLKBUF1 CLKBUF1_insert909 (
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf2)
);

CLKBUF1 CLKBUF1_insert908 (
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf3)
);

CLKBUF1 CLKBUF1_insert907 (
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf4)
);

CLKBUF1 CLKBUF1_insert906 (
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf5)
);

CLKBUF1 CLKBUF1_insert905 (
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf6)
);

CLKBUF1 CLKBUF1_insert904 (
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf7)
);

CLKBUF1 CLKBUF1_insert903 (
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf8)
);

CLKBUF1 CLKBUF1_insert902 (
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf9)
);

CLKBUF1 CLKBUF1_insert901 (
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf10)
);

CLKBUF1 CLKBUF1_insert900 (
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf11)
);

CLKBUF1 CLKBUF1_insert899 (
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf12)
);

CLKBUF1 CLKBUF1_insert898 (
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf13)
);

CLKBUF1 CLKBUF1_insert897 (
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf14)
);

CLKBUF1 CLKBUF1_insert896 (
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf15)
);

CLKBUF1 CLKBUF1_insert895 (
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf16)
);

CLKBUF1 CLKBUF1_insert894 (
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf17)
);

CLKBUF1 CLKBUF1_insert893 (
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf18)
);

CLKBUF1 CLKBUF1_insert892 (
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf19)
);

CLKBUF1 CLKBUF1_insert891 (
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf20)
);

CLKBUF1 CLKBUF1_insert890 (
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf21)
);

CLKBUF1 CLKBUF1_insert889 (
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf22)
);

CLKBUF1 CLKBUF1_insert888 (
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf23)
);

CLKBUF1 CLKBUF1_insert887 (
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf24)
);

CLKBUF1 CLKBUF1_insert886 (
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf25)
);

CLKBUF1 CLKBUF1_insert885 (
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf26)
);

CLKBUF1 CLKBUF1_insert884 (
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf27)
);

CLKBUF1 CLKBUF1_insert883 (
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf28)
);

CLKBUF1 CLKBUF1_insert882 (
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf29)
);

CLKBUF1 CLKBUF1_insert881 (
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf30)
);

CLKBUF1 CLKBUF1_insert880 (
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf31)
);

CLKBUF1 CLKBUF1_insert879 (
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf32)
);

CLKBUF1 CLKBUF1_insert878 (
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf33)
);

CLKBUF1 CLKBUF1_insert877 (
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf34)
);

CLKBUF1 CLKBUF1_insert876 (
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf35)
);

CLKBUF1 CLKBUF1_insert875 (
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf36)
);

CLKBUF1 CLKBUF1_insert874 (
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf37)
);

CLKBUF1 CLKBUF1_insert873 (
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf38)
);

CLKBUF1 CLKBUF1_insert872 (
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf39)
);

CLKBUF1 CLKBUF1_insert871 (
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf40)
);

CLKBUF1 CLKBUF1_insert870 (
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf41)
);

CLKBUF1 CLKBUF1_insert869 (
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf42)
);

CLKBUF1 CLKBUF1_insert868 (
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf43)
);

CLKBUF1 CLKBUF1_insert867 (
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf44)
);

CLKBUF1 CLKBUF1_insert866 (
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf45)
);

CLKBUF1 CLKBUF1_insert865 (
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf46)
);

CLKBUF1 CLKBUF1_insert864 (
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf47)
);

CLKBUF1 CLKBUF1_insert863 (
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf48)
);

CLKBUF1 CLKBUF1_insert862 (
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf49)
);

CLKBUF1 CLKBUF1_insert861 (
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf50)
);

CLKBUF1 CLKBUF1_insert860 (
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf51)
);

CLKBUF1 CLKBUF1_insert859 (
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf52)
);

CLKBUF1 CLKBUF1_insert858 (
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf53)
);

CLKBUF1 CLKBUF1_insert857 (
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf54)
);

CLKBUF1 CLKBUF1_insert856 (
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf55)
);

CLKBUF1 CLKBUF1_insert855 (
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf56)
);

CLKBUF1 CLKBUF1_insert854 (
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf57)
);

CLKBUF1 CLKBUF1_insert853 (
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf58)
);

CLKBUF1 CLKBUF1_insert852 (
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf59)
);

CLKBUF1 CLKBUF1_insert851 (
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf60)
);

CLKBUF1 CLKBUF1_insert850 (
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf61)
);

CLKBUF1 CLKBUF1_insert849 (
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf62)
);

CLKBUF1 CLKBUF1_insert848 (
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf63)
);

CLKBUF1 CLKBUF1_insert847 (
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf64)
);

CLKBUF1 CLKBUF1_insert846 (
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf65)
);

CLKBUF1 CLKBUF1_insert845 (
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf66)
);

CLKBUF1 CLKBUF1_insert844 (
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf67)
);

CLKBUF1 CLKBUF1_insert843 (
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf68)
);

CLKBUF1 CLKBUF1_insert842 (
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf69)
);

CLKBUF1 CLKBUF1_insert841 (
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf70)
);

CLKBUF1 CLKBUF1_insert840 (
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf71)
);

CLKBUF1 CLKBUF1_insert839 (
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf72)
);

CLKBUF1 CLKBUF1_insert838 (
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf73)
);

CLKBUF1 CLKBUF1_insert837 (
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf74)
);

CLKBUF1 CLKBUF1_insert836 (
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf75)
);

CLKBUF1 CLKBUF1_insert835 (
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf76)
);

CLKBUF1 CLKBUF1_insert834 (
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf77)
);

CLKBUF1 CLKBUF1_insert833 (
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf78)
);

CLKBUF1 CLKBUF1_insert832 (
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf79)
);

CLKBUF1 CLKBUF1_insert831 (
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf80)
);

CLKBUF1 CLKBUF1_insert830 (
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf81)
);

CLKBUF1 CLKBUF1_insert829 (
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf82)
);

CLKBUF1 CLKBUF1_insert828 (
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf83)
);

CLKBUF1 CLKBUF1_insert827 (
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf84)
);

CLKBUF1 CLKBUF1_insert826 (
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf85)
);

CLKBUF1 CLKBUF1_insert825 (
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf86)
);

CLKBUF1 CLKBUF1_insert824 (
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf87)
);

CLKBUF1 CLKBUF1_insert823 (
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf88)
);

CLKBUF1 CLKBUF1_insert822 (
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf89)
);

CLKBUF1 CLKBUF1_insert821 (
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf90)
);

CLKBUF1 CLKBUF1_insert820 (
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf91)
);

CLKBUF1 CLKBUF1_insert819 (
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf92)
);

CLKBUF1 CLKBUF1_insert818 (
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf93)
);

CLKBUF1 CLKBUF1_insert817 (
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf94)
);

CLKBUF1 CLKBUF1_insert816 (
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf95)
);

CLKBUF1 CLKBUF1_insert815 (
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf96)
);

CLKBUF1 CLKBUF1_insert814 (
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf97)
);

CLKBUF1 CLKBUF1_insert813 (
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf98)
);

CLKBUF1 CLKBUF1_insert812 (
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf99)
);

CLKBUF1 CLKBUF1_insert811 (
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf100)
);

CLKBUF1 CLKBUF1_insert810 (
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf101)
);

CLKBUF1 CLKBUF1_insert809 (
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf102)
);

CLKBUF1 CLKBUF1_insert808 (
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf103)
);

CLKBUF1 CLKBUF1_insert807 (
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf104)
);

CLKBUF1 CLKBUF1_insert806 (
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf105)
);

CLKBUF1 CLKBUF1_insert805 (
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf106)
);

CLKBUF1 CLKBUF1_insert804 (
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf107)
);

CLKBUF1 CLKBUF1_insert803 (
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf108)
);

CLKBUF1 CLKBUF1_insert802 (
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf109)
);

CLKBUF1 CLKBUF1_insert801 (
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf110)
);

CLKBUF1 CLKBUF1_insert800 (
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf111)
);

CLKBUF1 CLKBUF1_insert799 (
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf112)
);

CLKBUF1 CLKBUF1_insert798 (
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf113)
);

CLKBUF1 CLKBUF1_insert797 (
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf114)
);

CLKBUF1 CLKBUF1_insert796 (
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf115)
);

CLKBUF1 CLKBUF1_insert795 (
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf116)
);

CLKBUF1 CLKBUF1_insert794 (
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf117)
);

CLKBUF1 CLKBUF1_insert793 (
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf118)
);

CLKBUF1 CLKBUF1_insert792 (
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf119)
);

CLKBUF1 CLKBUF1_insert791 (
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf120)
);

CLKBUF1 CLKBUF1_insert790 (
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf121)
);

CLKBUF1 CLKBUF1_insert789 (
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf122)
);

CLKBUF1 CLKBUF1_insert788 (
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf123)
);

CLKBUF1 CLKBUF1_insert787 (
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf124)
);

CLKBUF1 CLKBUF1_insert786 (
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf125)
);

CLKBUF1 CLKBUF1_insert785 (
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf126)
);

CLKBUF1 CLKBUF1_insert784 (
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf127)
);

CLKBUF1 CLKBUF1_insert783 (
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf128)
);

CLKBUF1 CLKBUF1_insert782 (
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf129)
);

CLKBUF1 CLKBUF1_insert781 (
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf130)
);

CLKBUF1 CLKBUF1_insert780 (
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf131)
);

CLKBUF1 CLKBUF1_insert779 (
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf132)
);

CLKBUF1 CLKBUF1_insert778 (
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf133)
);

CLKBUF1 CLKBUF1_insert777 (
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf134)
);

CLKBUF1 CLKBUF1_insert776 (
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf135)
);

CLKBUF1 CLKBUF1_insert775 (
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf136)
);

CLKBUF1 CLKBUF1_insert774 (
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf137)
);

CLKBUF1 CLKBUF1_insert773 (
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf138)
);

CLKBUF1 CLKBUF1_insert772 (
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf139)
);

CLKBUF1 CLKBUF1_insert771 (
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf140)
);

CLKBUF1 CLKBUF1_insert770 (
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf141)
);

CLKBUF1 CLKBUF1_insert769 (
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf142)
);

CLKBUF1 CLKBUF1_insert768 (
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf143)
);

CLKBUF1 CLKBUF1_insert767 (
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf144)
);

CLKBUF1 CLKBUF1_insert766 (
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf145)
);

CLKBUF1 CLKBUF1_insert765 (
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf146)
);

CLKBUF1 CLKBUF1_insert764 (
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf147)
);

CLKBUF1 CLKBUF1_insert763 (
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf148)
);

CLKBUF1 CLKBUF1_insert762 (
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf149)
);

CLKBUF1 CLKBUF1_insert761 (
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf150)
);

CLKBUF1 CLKBUF1_insert760 (
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf151)
);

BUFX2 BUFX2_insert759 (
    .A(_4841_),
    .Y(_4841__bF$buf0)
);

BUFX2 BUFX2_insert758 (
    .A(_4841_),
    .Y(_4841__bF$buf1)
);

BUFX2 BUFX2_insert757 (
    .A(_4841_),
    .Y(_4841__bF$buf2)
);

BUFX2 BUFX2_insert756 (
    .A(_4841_),
    .Y(_4841__bF$buf3)
);

BUFX2 BUFX2_insert755 (
    .A(_4841_),
    .Y(_4841__bF$buf4)
);

BUFX2 BUFX2_insert754 (
    .A(_5341_),
    .Y(_5341__bF$buf0)
);

BUFX2 BUFX2_insert753 (
    .A(_5341_),
    .Y(_5341__bF$buf1)
);

BUFX2 BUFX2_insert752 (
    .A(_5341_),
    .Y(_5341__bF$buf2)
);

BUFX2 BUFX2_insert751 (
    .A(_5341_),
    .Y(_5341__bF$buf3)
);

BUFX2 BUFX2_insert750 (
    .A(_5341_),
    .Y(_5341__bF$buf4)
);

BUFX2 BUFX2_insert749 (
    .A(_5341_),
    .Y(_5341__bF$buf5)
);

BUFX2 BUFX2_insert748 (
    .A(_4803_),
    .Y(_4803__bF$buf0)
);

BUFX2 BUFX2_insert747 (
    .A(_4803_),
    .Y(_4803__bF$buf1)
);

BUFX2 BUFX2_insert746 (
    .A(_4803_),
    .Y(_4803__bF$buf2)
);

BUFX2 BUFX2_insert745 (
    .A(_4803_),
    .Y(_4803__bF$buf3)
);

BUFX2 BUFX2_insert744 (
    .A(_4803_),
    .Y(_4803__bF$buf4)
);

BUFX2 BUFX2_insert743 (
    .A(_4900_),
    .Y(_4900__bF$buf0)
);

BUFX2 BUFX2_insert742 (
    .A(_4900_),
    .Y(_4900__bF$buf1)
);

BUFX2 BUFX2_insert741 (
    .A(_4900_),
    .Y(_4900__bF$buf2)
);

BUFX2 BUFX2_insert740 (
    .A(_4900_),
    .Y(_4900__bF$buf3)
);

BUFX2 BUFX2_insert739 (
    .A(_4900_),
    .Y(_4900__bF$buf4)
);

BUFX2 BUFX2_insert738 (
    .A(\controlunit.csrfile_trap_wen ),
    .Y(\controlunit.csrfile_trap_wen_bF$buf0 )
);

BUFX2 BUFX2_insert737 (
    .A(\controlunit.csrfile_trap_wen ),
    .Y(\controlunit.csrfile_trap_wen_bF$buf1 )
);

BUFX2 BUFX2_insert736 (
    .A(\controlunit.csrfile_trap_wen ),
    .Y(\controlunit.csrfile_trap_wen_bF$buf2 )
);

BUFX2 BUFX2_insert735 (
    .A(\controlunit.csrfile_trap_wen ),
    .Y(\controlunit.csrfile_trap_wen_bF$buf3 )
);

BUFX2 BUFX2_insert734 (
    .A(\controlunit.csrfile_trap_wen ),
    .Y(\controlunit.csrfile_trap_wen_bF$buf4 )
);

BUFX2 BUFX2_insert733 (
    .A(\controlunit.csrfile_trap_wen ),
    .Y(\controlunit.csrfile_trap_wen_bF$buf5 )
);

BUFX2 BUFX2_insert732 (
    .A(\controlunit.csrfile_trap_wen ),
    .Y(\controlunit.csrfile_trap_wen_bF$buf6 )
);

BUFX2 BUFX2_insert731 (
    .A(\controlunit.csrfile_trap_wen ),
    .Y(\controlunit.csrfile_trap_wen_bF$buf7 )
);

BUFX2 BUFX2_insert730 (
    .A(_3410_),
    .Y(_3410__bF$buf0)
);

BUFX2 BUFX2_insert729 (
    .A(_3410_),
    .Y(_3410__bF$buf1)
);

BUFX2 BUFX2_insert728 (
    .A(_3410_),
    .Y(_3410__bF$buf2)
);

BUFX2 BUFX2_insert727 (
    .A(_3410_),
    .Y(_3410__bF$buf3)
);

BUFX2 BUFX2_insert726 (
    .A(_2014_),
    .Y(_2014__bF$buf0)
);

BUFX2 BUFX2_insert725 (
    .A(_2014_),
    .Y(_2014__bF$buf1)
);

BUFX2 BUFX2_insert724 (
    .A(_2014_),
    .Y(_2014__bF$buf2)
);

BUFX2 BUFX2_insert723 (
    .A(_2014_),
    .Y(_2014__bF$buf3)
);

BUFX2 BUFX2_insert722 (
    .A(_4847_),
    .Y(_4847__bF$buf0)
);

BUFX2 BUFX2_insert721 (
    .A(_4847_),
    .Y(_4847__bF$buf1)
);

BUFX2 BUFX2_insert720 (
    .A(_4847_),
    .Y(_4847__bF$buf2)
);

BUFX2 BUFX2_insert719 (
    .A(_4847_),
    .Y(_4847__bF$buf3)
);

BUFX2 BUFX2_insert718 (
    .A(_4847_),
    .Y(_4847__bF$buf4)
);

BUFX2 BUFX2_insert717 (
    .A(_4809_),
    .Y(_4809__bF$buf0)
);

BUFX2 BUFX2_insert716 (
    .A(_4809_),
    .Y(_4809__bF$buf1)
);

BUFX2 BUFX2_insert715 (
    .A(_4809_),
    .Y(_4809__bF$buf2)
);

BUFX2 BUFX2_insert714 (
    .A(_4809_),
    .Y(_4809__bF$buf3)
);

BUFX2 BUFX2_insert713 (
    .A(_4809_),
    .Y(_4809__bF$buf4)
);

BUFX2 BUFX2_insert712 (
    .A(_5118_),
    .Y(_5118__bF$buf0)
);

BUFX2 BUFX2_insert711 (
    .A(_5118_),
    .Y(_5118__bF$buf1)
);

BUFX2 BUFX2_insert710 (
    .A(_5118_),
    .Y(_5118__bF$buf2)
);

BUFX2 BUFX2_insert709 (
    .A(_5118_),
    .Y(_5118__bF$buf3)
);

BUFX2 BUFX2_insert708 (
    .A(_5118_),
    .Y(_5118__bF$buf4)
);

BUFX2 BUFX2_insert707 (
    .A(_5118_),
    .Y(_5118__bF$buf5)
);

BUFX2 BUFX2_insert706 (
    .A(_5118_),
    .Y(_5118__bF$buf6)
);

BUFX2 BUFX2_insert705 (
    .A(_5118_),
    .Y(_5118__bF$buf7)
);

BUFX2 BUFX2_insert704 (
    .A(_4794_),
    .Y(_4794__bF$buf0)
);

BUFX2 BUFX2_insert703 (
    .A(_4794_),
    .Y(_4794__bF$buf1)
);

BUFX2 BUFX2_insert702 (
    .A(_4794_),
    .Y(_4794__bF$buf2)
);

BUFX2 BUFX2_insert701 (
    .A(_4794_),
    .Y(_4794__bF$buf3)
);

BUFX2 BUFX2_insert700 (
    .A(_4794_),
    .Y(_4794__bF$buf4)
);

BUFX2 BUFX2_insert699 (
    .A(_4794_),
    .Y(_4794__bF$buf5)
);

BUFX2 BUFX2_insert698 (
    .A(_4794_),
    .Y(_4794__bF$buf6)
);

BUFX2 BUFX2_insert697 (
    .A(_4794_),
    .Y(_4794__bF$buf7)
);

BUFX2 BUFX2_insert696 (
    .A(_4853_),
    .Y(_4853__bF$buf0)
);

BUFX2 BUFX2_insert695 (
    .A(_4853_),
    .Y(_4853__bF$buf1)
);

BUFX2 BUFX2_insert694 (
    .A(_4853_),
    .Y(_4853__bF$buf2)
);

BUFX2 BUFX2_insert693 (
    .A(_4853_),
    .Y(_4853__bF$buf3)
);

BUFX2 BUFX2_insert692 (
    .A(_4853_),
    .Y(_4853__bF$buf4)
);

BUFX2 BUFX2_insert691 (
    .A(_184_),
    .Y(_184__bF$buf0)
);

BUFX2 BUFX2_insert690 (
    .A(_184_),
    .Y(_184__bF$buf1)
);

BUFX2 BUFX2_insert689 (
    .A(_184_),
    .Y(_184__bF$buf2)
);

BUFX2 BUFX2_insert688 (
    .A(_184_),
    .Y(_184__bF$buf3)
);

BUFX2 BUFX2_insert687 (
    .A(_184_),
    .Y(_184__bF$buf4)
);

BUFX2 BUFX2_insert686 (
    .A(_4815_),
    .Y(_4815__bF$buf0)
);

BUFX2 BUFX2_insert685 (
    .A(_4815_),
    .Y(_4815__bF$buf1)
);

BUFX2 BUFX2_insert684 (
    .A(_4815_),
    .Y(_4815__bF$buf2)
);

BUFX2 BUFX2_insert683 (
    .A(_4815_),
    .Y(_4815__bF$buf3)
);

BUFX2 BUFX2_insert682 (
    .A(_4815_),
    .Y(_4815__bF$buf4)
);

BUFX2 BUFX2_insert681 (
    .A(_3134_),
    .Y(_3134__bF$buf0)
);

BUFX2 BUFX2_insert680 (
    .A(_3134_),
    .Y(_3134__bF$buf1)
);

BUFX2 BUFX2_insert679 (
    .A(_3134_),
    .Y(_3134__bF$buf2)
);

BUFX2 BUFX2_insert678 (
    .A(_3134_),
    .Y(_3134__bF$buf3)
);

BUFX2 BUFX2_insert677 (
    .A(_3134_),
    .Y(_3134__bF$buf4)
);

BUFX2 BUFX2_insert676 (
    .A(_3134_),
    .Y(_3134__bF$buf5)
);

BUFX2 BUFX2_insert675 (
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_bF$buf0 )
);

BUFX2 BUFX2_insert674 (
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_bF$buf1 )
);

BUFX2 BUFX2_insert673 (
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_bF$buf2 )
);

BUFX2 BUFX2_insert672 (
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_bF$buf3 )
);

BUFX2 BUFX2_insert671 (
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_bF$buf4 )
);

BUFX2 BUFX2_insert670 (
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_bF$buf5 )
);

BUFX2 BUFX2_insert669 (
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_bF$buf6 )
);

BUFX2 BUFX2_insert668 (
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_bF$buf7 )
);

BUFX2 BUFX2_insert667 (
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_bF$buf8 )
);

BUFX2 BUFX2_insert666 (
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_bF$buf9 )
);

BUFX2 BUFX2_insert665 (
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_bF$buf10 )
);

BUFX2 BUFX2_insert664 (
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_bF$buf11 )
);

BUFX2 BUFX2_insert663 (
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_bF$buf12 )
);

BUFX2 BUFX2_insert662 (
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_bF$buf13 )
);

BUFX2 BUFX2_insert661 (
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_bF$buf14 )
);

BUFX2 BUFX2_insert660 (
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_bF$buf15 )
);

BUFX2 BUFX2_insert659 (
    .A(_9092_),
    .Y(_9092__bF$buf0)
);

BUFX2 BUFX2_insert658 (
    .A(_9092_),
    .Y(_9092__bF$buf1)
);

BUFX2 BUFX2_insert657 (
    .A(_9092_),
    .Y(_9092__bF$buf2)
);

BUFX2 BUFX2_insert656 (
    .A(_9092_),
    .Y(_9092__bF$buf3)
);

BUFX2 BUFX2_insert655 (
    .A(_9092_),
    .Y(_9092__bF$buf4)
);

BUFX2 BUFX2_insert654 (
    .A(_9092_),
    .Y(_9092__bF$buf5)
);

BUFX2 BUFX2_insert653 (
    .A(_9092_),
    .Y(_9092__bF$buf6)
);

BUFX2 BUFX2_insert652 (
    .A(_9092_),
    .Y(_9092__bF$buf7)
);

BUFX2 BUFX2_insert651 (
    .A(_9092_),
    .Y(_9092__bF$buf8)
);

BUFX2 BUFX2_insert650 (
    .A(_187_),
    .Y(_187__bF$buf0)
);

BUFX2 BUFX2_insert649 (
    .A(_187_),
    .Y(_187__bF$buf1)
);

BUFX2 BUFX2_insert648 (
    .A(_187_),
    .Y(_187__bF$buf2)
);

BUFX2 BUFX2_insert647 (
    .A(_187_),
    .Y(_187__bF$buf3)
);

BUFX2 BUFX2_insert646 (
    .A(_187_),
    .Y(_187__bF$buf4)
);

BUFX2 BUFX2_insert645 (
    .A(\datapath.idinstr_20_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_20_bF$buf0 )
);

BUFX2 BUFX2_insert644 (
    .A(\datapath.idinstr_20_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_20_bF$buf1 )
);

BUFX2 BUFX2_insert643 (
    .A(\datapath.idinstr_20_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_20_bF$buf2 )
);

BUFX2 BUFX2_insert642 (
    .A(\datapath.idinstr_20_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_20_bF$buf3 )
);

BUFX2 BUFX2_insert641 (
    .A(\datapath.idinstr_20_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_20_bF$buf4 )
);

BUFX2 BUFX2_insert640 (
    .A(\datapath.idinstr_20_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_20_bF$buf5 )
);

BUFX2 BUFX2_insert639 (
    .A(\datapath.idinstr_20_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_20_bF$buf6 )
);

BUFX2 BUFX2_insert638 (
    .A(\datapath.idinstr_20_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_20_bF$buf7 )
);

BUFX2 BUFX2_insert637 (
    .A(\datapath.idinstr_20_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_20_bF$buf8 )
);

BUFX2 BUFX2_insert636 (
    .A(\datapath.idinstr_20_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_20_bF$buf9 )
);

BUFX2 BUFX2_insert635 (
    .A(\datapath.idinstr_20_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_20_bF$buf10 )
);

BUFX2 BUFX2_insert634 (
    .A(\datapath.idinstr_20_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_20_bF$buf11 )
);

BUFX2 BUFX2_insert633 (
    .A(\datapath.idinstr_20_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_20_bF$buf12 )
);

BUFX2 BUFX2_insert632 (
    .A(\datapath.idinstr_20_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_20_bF$buf13 )
);

BUFX2 BUFX2_insert631 (
    .A(\datapath.idinstr_20_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_20_bF$buf14 )
);

BUFX2 BUFX2_insert630 (
    .A(\datapath.idinstr_20_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_20_bF$buf15 )
);

BUFX2 BUFX2_insert629 (
    .A(\datapath.idinstr_20_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_20_bF$buf16 )
);

BUFX2 BUFX2_insert628 (
    .A(\datapath.idinstr_20_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_20_bF$buf17 )
);

BUFX2 BUFX2_insert627 (
    .A(\datapath.idinstr_20_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_20_bF$buf18 )
);

BUFX2 BUFX2_insert626 (
    .A(\datapath.idinstr_20_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_20_bF$buf19 )
);

BUFX2 BUFX2_insert625 (
    .A(\datapath.idinstr_20_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_20_bF$buf20 )
);

BUFX2 BUFX2_insert624 (
    .A(\datapath.idinstr_20_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_20_bF$buf21 )
);

BUFX2 BUFX2_insert623 (
    .A(\datapath.idinstr_20_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_20_bF$buf22 )
);

BUFX2 BUFX2_insert622 (
    .A(\datapath.idinstr_20_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_20_bF$buf23 )
);

BUFX2 BUFX2_insert621 (
    .A(\datapath.idinstr_20_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_20_bF$buf24 )
);

BUFX2 BUFX2_insert620 (
    .A(\datapath.idinstr_20_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_20_bF$buf25 )
);

BUFX2 BUFX2_insert619 (
    .A(\datapath.idinstr_20_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_20_bF$buf26 )
);

BUFX2 BUFX2_insert618 (
    .A(\datapath.idinstr_20_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_20_bF$buf27 )
);

BUFX2 BUFX2_insert617 (
    .A(\datapath.idinstr_20_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_20_bF$buf28 )
);

BUFX2 BUFX2_insert616 (
    .A(\datapath.idinstr_20_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_20_bF$buf29 )
);

BUFX2 BUFX2_insert615 (
    .A(\datapath.idinstr_20_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_20_bF$buf30 )
);

BUFX2 BUFX2_insert614 (
    .A(\datapath.idinstr_20_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_20_bF$buf31 )
);

BUFX2 BUFX2_insert613 (
    .A(\datapath.idinstr_20_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_20_bF$buf32 )
);

BUFX2 BUFX2_insert612 (
    .A(\datapath.idinstr_20_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_20_bF$buf33 )
);

BUFX2 BUFX2_insert611 (
    .A(\datapath.idinstr_20_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_20_bF$buf34 )
);

BUFX2 BUFX2_insert610 (
    .A(\datapath.idinstr_20_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_20_bF$buf35 )
);

BUFX2 BUFX2_insert609 (
    .A(\datapath.idinstr_20_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_20_bF$buf36 )
);

BUFX2 BUFX2_insert608 (
    .A(\datapath.idinstr_20_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_20_bF$buf37 )
);

BUFX2 BUFX2_insert607 (
    .A(\datapath.idinstr_20_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_20_bF$buf38 )
);

BUFX2 BUFX2_insert606 (
    .A(\datapath.idinstr_20_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_20_bF$buf39 )
);

BUFX2 BUFX2_insert605 (
    .A(\datapath.idinstr_20_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_20_bF$buf40 )
);

BUFX2 BUFX2_insert604 (
    .A(\datapath.idinstr_20_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_20_bF$buf41 )
);

BUFX2 BUFX2_insert603 (
    .A(\datapath.idinstr_20_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_20_bF$buf42 )
);

BUFX2 BUFX2_insert602 (
    .A(\datapath.idinstr_20_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_20_bF$buf43 )
);

BUFX2 BUFX2_insert601 (
    .A(\datapath.idinstr_20_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_20_bF$buf44 )
);

BUFX2 BUFX2_insert600 (
    .A(\datapath.idinstr_20_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_20_bF$buf45 )
);

BUFX2 BUFX2_insert599 (
    .A(\datapath.idinstr_20_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_20_bF$buf46 )
);

BUFX2 BUFX2_insert598 (
    .A(\datapath.idinstr_20_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_20_bF$buf47 )
);

BUFX2 BUFX2_insert597 (
    .A(\datapath.idinstr_20_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_20_bF$buf48 )
);

BUFX2 BUFX2_insert596 (
    .A(\datapath.idinstr_20_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_20_bF$buf49 )
);

BUFX2 BUFX2_insert595 (
    .A(\datapath.idinstr_20_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_20_bF$buf50 )
);

BUFX2 BUFX2_insert594 (
    .A(\datapath.idinstr_20_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_20_bF$buf51 )
);

BUFX2 BUFX2_insert593 (
    .A(\datapath.idinstr_20_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_20_bF$buf52 )
);

BUFX2 BUFX2_insert592 (
    .A(\datapath.idinstr_20_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_20_bF$buf53 )
);

BUFX2 BUFX2_insert591 (
    .A(\datapath.idinstr_20_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_20_bF$buf54 )
);

BUFX2 BUFX2_insert590 (
    .A(\datapath.idinstr_20_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_20_bF$buf55 )
);

BUFX2 BUFX2_insert589 (
    .A(_0_[1]),
    .Y(_0__1_bF$buf0)
);

BUFX2 BUFX2_insert588 (
    .A(_0_[1]),
    .Y(_0__1_bF$buf1)
);

BUFX2 BUFX2_insert587 (
    .A(_0_[1]),
    .Y(_0__1_bF$buf2)
);

BUFX2 BUFX2_insert586 (
    .A(_0_[1]),
    .Y(_0__1_bF$buf3)
);

BUFX2 BUFX2_insert585 (
    .A(_0_[1]),
    .Y(_0__1_bF$buf4)
);

BUFX2 BUFX2_insert584 (
    .A(_0_[1]),
    .Y(_0__1_bF$buf5)
);

BUFX2 BUFX2_insert583 (
    .A(_0_[1]),
    .Y(_0__1_bF$buf6)
);

BUFX2 BUFX2_insert582 (
    .A(_0_[1]),
    .Y(_0__1_bF$buf7)
);

BUFX2 BUFX2_insert581 (
    .A(_0_[1]),
    .Y(_0__1_bF$buf8)
);

BUFX2 BUFX2_insert580 (
    .A(_0_[1]),
    .Y(_0__1_bF$buf9)
);

BUFX2 BUFX2_insert579 (
    .A(_0_[1]),
    .Y(_0__1_bF$buf10)
);

BUFX2 BUFX2_insert578 (
    .A(_4821_),
    .Y(_4821__bF$buf0)
);

BUFX2 BUFX2_insert577 (
    .A(_4821_),
    .Y(_4821__bF$buf1)
);

BUFX2 BUFX2_insert576 (
    .A(_4821_),
    .Y(_4821__bF$buf2)
);

BUFX2 BUFX2_insert575 (
    .A(_4821_),
    .Y(_4821__bF$buf3)
);

BUFX2 BUFX2_insert574 (
    .A(_4821_),
    .Y(_4821__bF$buf4)
);

BUFX2 BUFX2_insert573 (
    .A(_3557_),
    .Y(_3557__bF$buf0)
);

BUFX2 BUFX2_insert572 (
    .A(_3557_),
    .Y(_3557__bF$buf1)
);

BUFX2 BUFX2_insert571 (
    .A(_3557_),
    .Y(_3557__bF$buf2)
);

BUFX2 BUFX2_insert570 (
    .A(_3557_),
    .Y(_3557__bF$buf3)
);

BUFX2 BUFX2_insert569 (
    .A(_3557_),
    .Y(_3557__bF$buf4)
);

BUFX2 BUFX2_insert568 (
    .A(_4859_),
    .Y(_4859__bF$buf0)
);

BUFX2 BUFX2_insert567 (
    .A(_4859_),
    .Y(_4859__bF$buf1)
);

BUFX2 BUFX2_insert566 (
    .A(_4859_),
    .Y(_4859__bF$buf2)
);

BUFX2 BUFX2_insert565 (
    .A(_4859_),
    .Y(_4859__bF$buf3)
);

BUFX2 BUFX2_insert564 (
    .A(_4859_),
    .Y(_4859__bF$buf4)
);

BUFX2 BUFX2_insert563 (
    .A(\datapath.idinstr [23]),
    .Y(\datapath.idinstr_23_bF$buf0 )
);

BUFX2 BUFX2_insert562 (
    .A(\datapath.idinstr [23]),
    .Y(\datapath.idinstr_23_bF$buf1 )
);

BUFX2 BUFX2_insert561 (
    .A(\datapath.idinstr [23]),
    .Y(\datapath.idinstr_23_bF$buf2 )
);

BUFX2 BUFX2_insert560 (
    .A(\datapath.idinstr [23]),
    .Y(\datapath.idinstr_23_bF$buf3 )
);

BUFX2 BUFX2_insert559 (
    .A(\datapath.idinstr [23]),
    .Y(\datapath.idinstr_23_bF$buf4 )
);

BUFX2 BUFX2_insert558 (
    .A(\datapath.idinstr [23]),
    .Y(\datapath.idinstr_23_bF$buf5 )
);

BUFX2 BUFX2_insert557 (
    .A(\datapath.idinstr [23]),
    .Y(\datapath.idinstr_23_bF$buf6 )
);

BUFX2 BUFX2_insert556 (
    .A(_287_),
    .Y(_287__bF$buf0)
);

BUFX2 BUFX2_insert555 (
    .A(_287_),
    .Y(_287__bF$buf1)
);

BUFX2 BUFX2_insert554 (
    .A(_287_),
    .Y(_287__bF$buf2)
);

BUFX2 BUFX2_insert553 (
    .A(_287_),
    .Y(_287__bF$buf3)
);

BUFX2 BUFX2_insert552 (
    .A(_287_),
    .Y(_287__bF$buf4)
);

BUFX2 BUFX2_insert551 (
    .A(_3563_),
    .Y(_3563__bF$buf0)
);

BUFX2 BUFX2_insert550 (
    .A(_3563_),
    .Y(_3563__bF$buf1)
);

BUFX2 BUFX2_insert549 (
    .A(_3563_),
    .Y(_3563__bF$buf2)
);

BUFX2 BUFX2_insert548 (
    .A(_3563_),
    .Y(_3563__bF$buf3)
);

BUFX2 BUFX2_insert547 (
    .A(_3563_),
    .Y(_3563__bF$buf4)
);

BUFX2 BUFX2_insert546 (
    .A(_9025_),
    .Y(_9025__bF$buf0)
);

BUFX2 BUFX2_insert545 (
    .A(_9025_),
    .Y(_9025__bF$buf1)
);

BUFX2 BUFX2_insert544 (
    .A(_9025_),
    .Y(_9025__bF$buf2)
);

BUFX2 BUFX2_insert543 (
    .A(_9025_),
    .Y(_9025__bF$buf3)
);

BUFX2 BUFX2_insert542 (
    .A(_9025_),
    .Y(_9025__bF$buf4)
);

BUFX2 BUFX2_insert541 (
    .A(_4827_),
    .Y(_4827__bF$buf0)
);

BUFX2 BUFX2_insert540 (
    .A(_4827_),
    .Y(_4827__bF$buf1)
);

BUFX2 BUFX2_insert539 (
    .A(_4827_),
    .Y(_4827__bF$buf2)
);

BUFX2 BUFX2_insert538 (
    .A(_4827_),
    .Y(_4827__bF$buf3)
);

BUFX2 BUFX2_insert537 (
    .A(_4827_),
    .Y(_4827__bF$buf4)
);

BUFX2 BUFX2_insert536 (
    .A(_387_),
    .Y(_387__bF$buf0)
);

BUFX2 BUFX2_insert535 (
    .A(_387_),
    .Y(_387__bF$buf1)
);

BUFX2 BUFX2_insert534 (
    .A(_387_),
    .Y(_387__bF$buf2)
);

BUFX2 BUFX2_insert533 (
    .A(_387_),
    .Y(_387__bF$buf3)
);

BUFX2 BUFX2_insert532 (
    .A(_387_),
    .Y(_387__bF$buf4)
);

BUFX2 BUFX2_insert531 (
    .A(_5653_),
    .Y(_5653__bF$buf0)
);

BUFX2 BUFX2_insert530 (
    .A(_5653_),
    .Y(_5653__bF$buf1)
);

BUFX2 BUFX2_insert529 (
    .A(_5653_),
    .Y(_5653__bF$buf2)
);

BUFX2 BUFX2_insert528 (
    .A(_5653_),
    .Y(_5653__bF$buf3)
);

BUFX2 BUFX2_insert527 (
    .A(_5653_),
    .Y(_5653__bF$buf4)
);

BUFX2 BUFX2_insert526 (
    .A(_5653_),
    .Y(_5653__bF$buf5)
);

BUFX2 BUFX2_insert525 (
    .A(_5653_),
    .Y(_5653__bF$buf6)
);

BUFX2 BUFX2_insert524 (
    .A(_5653_),
    .Y(_5653__bF$buf7)
);

BUFX2 BUFX2_insert523 (
    .A(_2781_),
    .Y(_2781__bF$buf0)
);

BUFX2 BUFX2_insert522 (
    .A(_2781_),
    .Y(_2781__bF$buf1)
);

BUFX2 BUFX2_insert521 (
    .A(_2781_),
    .Y(_2781__bF$buf2)
);

BUFX2 BUFX2_insert520 (
    .A(_2781_),
    .Y(_2781__bF$buf3)
);

BUFX2 BUFX2_insert519 (
    .A(_2781_),
    .Y(_2781__bF$buf4)
);

BUFX2 BUFX2_insert518 (
    .A(_3014_),
    .Y(_3014__bF$buf0)
);

BUFX2 BUFX2_insert517 (
    .A(_3014_),
    .Y(_3014__bF$buf1)
);

BUFX2 BUFX2_insert516 (
    .A(_3014_),
    .Y(_3014__bF$buf2)
);

BUFX2 BUFX2_insert515 (
    .A(_3014_),
    .Y(_3014__bF$buf3)
);

BUFX2 BUFX2_insert514 (
    .A(_3014_),
    .Y(_3014__bF$buf4)
);

BUFX2 BUFX2_insert513 (
    .A(_3014_),
    .Y(_3014__bF$buf5)
);

BUFX2 BUFX2_insert512 (
    .A(_3014_),
    .Y(_3014__bF$buf6)
);

BUFX2 BUFX2_insert511 (
    .A(\datapath.alu.b [1]),
    .Y(\datapath.alu.b_1_bF$buf0 )
);

BUFX2 BUFX2_insert510 (
    .A(\datapath.alu.b [1]),
    .Y(\datapath.alu.b_1_bF$buf1 )
);

BUFX2 BUFX2_insert509 (
    .A(\datapath.alu.b [1]),
    .Y(\datapath.alu.b_1_bF$buf2 )
);

BUFX2 BUFX2_insert508 (
    .A(\datapath.alu.b [1]),
    .Y(\datapath.alu.b_1_bF$buf3 )
);

BUFX2 BUFX2_insert507 (
    .A(\datapath.alu.b [1]),
    .Y(\datapath.alu.b_1_bF$buf4 )
);

BUFX2 BUFX2_insert506 (
    .A(\datapath.alu.b [1]),
    .Y(\datapath.alu.b_1_bF$buf5 )
);

BUFX2 BUFX2_insert505 (
    .A(\datapath.alu.b [1]),
    .Y(\datapath.alu.b_1_bF$buf6 )
);

BUFX2 BUFX2_insert504 (
    .A(_7420_),
    .Y(_7420__bF$buf0)
);

BUFX2 BUFX2_insert503 (
    .A(_7420_),
    .Y(_7420__bF$buf1)
);

BUFX2 BUFX2_insert502 (
    .A(_7420_),
    .Y(_7420__bF$buf2)
);

BUFX2 BUFX2_insert501 (
    .A(_7420_),
    .Y(_7420__bF$buf3)
);

BUFX2 BUFX2_insert500 (
    .A(_7420_),
    .Y(_7420__bF$buf4)
);

BUFX2 BUFX2_insert499 (
    .A(_7420_),
    .Y(_7420__bF$buf5)
);

BUFX2 BUFX2_insert498 (
    .A(_7420_),
    .Y(_7420__bF$buf6)
);

BUFX2 BUFX2_insert497 (
    .A(_7420_),
    .Y(_7420__bF$buf7)
);

BUFX2 BUFX2_insert496 (
    .A(_7420_),
    .Y(_7420__bF$buf8)
);

BUFX2 BUFX2_insert495 (
    .A(_7420_),
    .Y(_7420__bF$buf9)
);

BUFX2 BUFX2_insert494 (
    .A(_7420_),
    .Y(_7420__bF$buf10)
);

BUFX2 BUFX2_insert493 (
    .A(_9125_),
    .Y(_9125__bF$buf0)
);

BUFX2 BUFX2_insert492 (
    .A(_9125_),
    .Y(_9125__bF$buf1)
);

BUFX2 BUFX2_insert491 (
    .A(_9125_),
    .Y(_9125__bF$buf2)
);

BUFX2 BUFX2_insert490 (
    .A(_9125_),
    .Y(_9125__bF$buf3)
);

BUFX2 BUFX2_insert489 (
    .A(_9125_),
    .Y(_9125__bF$buf4)
);

BUFX2 BUFX2_insert488 (
    .A(_4833_),
    .Y(_4833__bF$buf0)
);

BUFX2 BUFX2_insert487 (
    .A(_4833_),
    .Y(_4833__bF$buf1)
);

BUFX2 BUFX2_insert486 (
    .A(_4833_),
    .Y(_4833__bF$buf2)
);

BUFX2 BUFX2_insert485 (
    .A(_4833_),
    .Y(_4833__bF$buf3)
);

BUFX2 BUFX2_insert484 (
    .A(_4833_),
    .Y(_4833__bF$buf4)
);

BUFX2 BUFX2_insert483 (
    .A(_2267_),
    .Y(_2267__bF$buf0)
);

BUFX2 BUFX2_insert482 (
    .A(_2267_),
    .Y(_2267__bF$buf1)
);

BUFX2 BUFX2_insert481 (
    .A(_2267_),
    .Y(_2267__bF$buf2)
);

BUFX2 BUFX2_insert480 (
    .A(_2267_),
    .Y(_2267__bF$buf3)
);

BUFX2 BUFX2_insert479 (
    .A(_3017_),
    .Y(_3017__bF$buf0)
);

BUFX2 BUFX2_insert478 (
    .A(_3017_),
    .Y(_3017__bF$buf1)
);

BUFX2 BUFX2_insert477 (
    .A(_3017_),
    .Y(_3017__bF$buf2)
);

BUFX2 BUFX2_insert476 (
    .A(_3017_),
    .Y(_3017__bF$buf3)
);

BUFX2 BUFX2_insert475 (
    .A(_3017_),
    .Y(_3017__bF$buf4)
);

BUFX2 BUFX2_insert474 (
    .A(\datapath.alu.b [4]),
    .Y(\datapath.alu.b_4_bF$buf0 )
);

BUFX2 BUFX2_insert473 (
    .A(\datapath.alu.b [4]),
    .Y(\datapath.alu.b_4_bF$buf1 )
);

BUFX2 BUFX2_insert472 (
    .A(\datapath.alu.b [4]),
    .Y(\datapath.alu.b_4_bF$buf2 )
);

BUFX2 BUFX2_insert471 (
    .A(\datapath.alu.b [4]),
    .Y(\datapath.alu.b_4_bF$buf3 )
);

BUFX2 BUFX2_insert470 (
    .A(\datapath.alu.b [4]),
    .Y(\datapath.alu.b_4_bF$buf4 )
);

BUFX2 BUFX2_insert469 (
    .A(_4968_),
    .Y(_4968__bF$buf0)
);

BUFX2 BUFX2_insert468 (
    .A(_4968_),
    .Y(_4968__bF$buf1)
);

BUFX2 BUFX2_insert467 (
    .A(_4968_),
    .Y(_4968__bF$buf2)
);

BUFX2 BUFX2_insert466 (
    .A(_4968_),
    .Y(_4968__bF$buf3)
);

BUFX2 BUFX2_insert465 (
    .A(_4968_),
    .Y(_4968__bF$buf4)
);

BUFX2 BUFX2_insert464 (
    .A(_4968_),
    .Y(_4968__bF$buf5)
);

BUFX2 BUFX2_insert463 (
    .A(_4968_),
    .Y(_4968__bF$buf6)
);

BUFX2 BUFX2_insert462 (
    .A(_4968_),
    .Y(_4968__bF$buf7)
);

BUFX2 BUFX2_insert461 (
    .A(_4968_),
    .Y(_4968__bF$buf8)
);

BUFX2 BUFX2_insert460 (
    .A(_4968_),
    .Y(_4968__bF$buf9)
);

BUFX2 BUFX2_insert459 (
    .A(_7423_),
    .Y(_7423__bF$buf0)
);

BUFX2 BUFX2_insert458 (
    .A(_7423_),
    .Y(_7423__bF$buf1)
);

BUFX2 BUFX2_insert457 (
    .A(_7423_),
    .Y(_7423__bF$buf2)
);

BUFX2 BUFX2_insert456 (
    .A(_7423_),
    .Y(_7423__bF$buf3)
);

BUFX2 BUFX2_insert455 (
    .A(_7423_),
    .Y(_7423__bF$buf4)
);

BUFX2 BUFX2_insert454 (
    .A(_7423_),
    .Y(_7423__bF$buf5)
);

BUFX2 BUFX2_insert453 (
    .A(_7423_),
    .Y(_7423__bF$buf6)
);

BUFX2 BUFX2_insert452 (
    .A(_7423_),
    .Y(_7423__bF$buf7)
);

BUFX2 BUFX2_insert451 (
    .A(_5756_),
    .Y(_5756__bF$buf0)
);

BUFX2 BUFX2_insert450 (
    .A(_5756_),
    .Y(_5756__bF$buf1)
);

BUFX2 BUFX2_insert449 (
    .A(_5756_),
    .Y(_5756__bF$buf2)
);

BUFX2 BUFX2_insert448 (
    .A(_5756_),
    .Y(_5756__bF$buf3)
);

BUFX2 BUFX2_insert447 (
    .A(_5756_),
    .Y(_5756__bF$buf4)
);

BUFX2 BUFX2_insert446 (
    .A(_5756_),
    .Y(_5756__bF$buf5)
);

BUFX2 BUFX2_insert445 (
    .A(_5756_),
    .Y(_5756__bF$buf6)
);

BUFX2 BUFX2_insert444 (
    .A(_5756_),
    .Y(_5756__bF$buf7)
);

BUFX2 BUFX2_insert443 (
    .A(_5756_),
    .Y(_5756__bF$buf8)
);

BUFX2 BUFX2_insert442 (
    .A(_5756_),
    .Y(_5756__bF$buf9)
);

BUFX2 BUFX2_insert441 (
    .A(_5051_),
    .Y(_5051__bF$buf0)
);

BUFX2 BUFX2_insert440 (
    .A(_5051_),
    .Y(_5051__bF$buf1)
);

BUFX2 BUFX2_insert439 (
    .A(_5051_),
    .Y(_5051__bF$buf2)
);

BUFX2 BUFX2_insert438 (
    .A(_5051_),
    .Y(_5051__bF$buf3)
);

BUFX2 BUFX2_insert437 (
    .A(_5051_),
    .Y(_5051__bF$buf4)
);

BUFX2 BUFX2_insert436 (
    .A(_5051_),
    .Y(_5051__bF$buf5)
);

BUFX2 BUFX2_insert435 (
    .A(_4801_),
    .Y(_4801__bF$buf0)
);

BUFX2 BUFX2_insert434 (
    .A(_4801_),
    .Y(_4801__bF$buf1)
);

BUFX2 BUFX2_insert433 (
    .A(_4801_),
    .Y(_4801__bF$buf2)
);

BUFX2 BUFX2_insert432 (
    .A(_4801_),
    .Y(_4801__bF$buf3)
);

BUFX2 BUFX2_insert431 (
    .A(_4801_),
    .Y(_4801__bF$buf4)
);

BUFX2 BUFX2_insert430 (
    .A(_5186_),
    .Y(_5186__bF$buf0)
);

BUFX2 BUFX2_insert429 (
    .A(_5186_),
    .Y(_5186__bF$buf1)
);

BUFX2 BUFX2_insert428 (
    .A(_5186_),
    .Y(_5186__bF$buf2)
);

BUFX2 BUFX2_insert427 (
    .A(_5186_),
    .Y(_5186__bF$buf3)
);

BUFX2 BUFX2_insert426 (
    .A(_5186_),
    .Y(_5186__bF$buf4)
);

BUFX2 BUFX2_insert425 (
    .A(_4839_),
    .Y(_4839__bF$buf0)
);

BUFX2 BUFX2_insert424 (
    .A(_4839_),
    .Y(_4839__bF$buf1)
);

BUFX2 BUFX2_insert423 (
    .A(_4839_),
    .Y(_4839__bF$buf2)
);

BUFX2 BUFX2_insert422 (
    .A(_4839_),
    .Y(_4839__bF$buf3)
);

BUFX2 BUFX2_insert421 (
    .A(_4839_),
    .Y(_4839__bF$buf4)
);

BUFX2 BUFX2_insert420 (
    .A(_5759_),
    .Y(_5759__bF$buf0)
);

BUFX2 BUFX2_insert419 (
    .A(_5759_),
    .Y(_5759__bF$buf1)
);

BUFX2 BUFX2_insert418 (
    .A(_5759_),
    .Y(_5759__bF$buf2)
);

BUFX2 BUFX2_insert417 (
    .A(_5759_),
    .Y(_5759__bF$buf3)
);

BUFX2 BUFX2_insert416 (
    .A(_5759_),
    .Y(_5759__bF$buf4)
);

BUFX2 BUFX2_insert415 (
    .A(_2047_),
    .Y(_2047__bF$buf0)
);

BUFX2 BUFX2_insert414 (
    .A(_2047_),
    .Y(_2047__bF$buf1)
);

BUFX2 BUFX2_insert413 (
    .A(_2047_),
    .Y(_2047__bF$buf2)
);

BUFX2 BUFX2_insert412 (
    .A(_2047_),
    .Y(_2047__bF$buf3)
);

BUFX2 BUFX2_insert411 (
    .A(_5342_),
    .Y(_5342__bF$buf0)
);

BUFX2 BUFX2_insert410 (
    .A(_5342_),
    .Y(_5342__bF$buf1)
);

BUFX2 BUFX2_insert409 (
    .A(_5342_),
    .Y(_5342__bF$buf2)
);

BUFX2 BUFX2_insert408 (
    .A(_5342_),
    .Y(_5342__bF$buf3)
);

BUFX2 BUFX2_insert407 (
    .A(_5342_),
    .Y(_5342__bF$buf4)
);

BUFX2 BUFX2_insert406 (
    .A(_5762__hier0_bF$buf5),
    .Y(_5762__bF$buf0)
);

BUFX2 BUFX2_insert405 (
    .A(_5762__hier0_bF$buf4),
    .Y(_5762__bF$buf1)
);

BUFX2 BUFX2_insert404 (
    .A(_5762__hier0_bF$buf3),
    .Y(_5762__bF$buf2)
);

BUFX2 BUFX2_insert403 (
    .A(_5762__hier0_bF$buf2),
    .Y(_5762__bF$buf3)
);

BUFX2 BUFX2_insert402 (
    .A(_5762__hier0_bF$buf1),
    .Y(_5762__bF$buf4)
);

BUFX2 BUFX2_insert401 (
    .A(_5762__hier0_bF$buf0),
    .Y(_5762__bF$buf5)
);

BUFX2 BUFX2_insert400 (
    .A(_5762__hier0_bF$buf5),
    .Y(_5762__bF$buf6)
);

BUFX2 BUFX2_insert399 (
    .A(_5762__hier0_bF$buf4),
    .Y(_5762__bF$buf7)
);

BUFX2 BUFX2_insert398 (
    .A(_5762__hier0_bF$buf3),
    .Y(_5762__bF$buf8)
);

BUFX2 BUFX2_insert397 (
    .A(_5762__hier0_bF$buf2),
    .Y(_5762__bF$buf9)
);

BUFX2 BUFX2_insert396 (
    .A(_5762__hier0_bF$buf1),
    .Y(_5762__bF$buf10)
);

BUFX2 BUFX2_insert395 (
    .A(_5762__hier0_bF$buf0),
    .Y(_5762__bF$buf11)
);

BUFX2 BUFX2_insert394 (
    .A(_5762__hier0_bF$buf5),
    .Y(_5762__bF$buf12)
);

BUFX2 BUFX2_insert393 (
    .A(_5762__hier0_bF$buf4),
    .Y(_5762__bF$buf13)
);

BUFX2 BUFX2_insert392 (
    .A(_5762__hier0_bF$buf3),
    .Y(_5762__bF$buf14)
);

BUFX2 BUFX2_insert391 (
    .A(_5762__hier0_bF$buf2),
    .Y(_5762__bF$buf15)
);

BUFX2 BUFX2_insert390 (
    .A(_5762__hier0_bF$buf1),
    .Y(_5762__bF$buf16)
);

BUFX2 BUFX2_insert389 (
    .A(_5762__hier0_bF$buf0),
    .Y(_5762__bF$buf17)
);

BUFX2 BUFX2_insert388 (
    .A(_5762__hier0_bF$buf5),
    .Y(_5762__bF$buf18)
);

BUFX2 BUFX2_insert387 (
    .A(_5762__hier0_bF$buf4),
    .Y(_5762__bF$buf19)
);

BUFX2 BUFX2_insert386 (
    .A(_5762__hier0_bF$buf3),
    .Y(_5762__bF$buf20)
);

BUFX2 BUFX2_insert385 (
    .A(_5762__hier0_bF$buf2),
    .Y(_5762__bF$buf21)
);

BUFX2 BUFX2_insert384 (
    .A(_5762__hier0_bF$buf1),
    .Y(_5762__bF$buf22)
);

BUFX2 BUFX2_insert383 (
    .A(_5762__hier0_bF$buf0),
    .Y(_5762__bF$buf23)
);

BUFX2 BUFX2_insert382 (
    .A(_5762__hier0_bF$buf5),
    .Y(_5762__bF$buf24)
);

BUFX2 BUFX2_insert381 (
    .A(_5762__hier0_bF$buf4),
    .Y(_5762__bF$buf25)
);

BUFX2 BUFX2_insert380 (
    .A(_5762__hier0_bF$buf3),
    .Y(_5762__bF$buf26)
);

BUFX2 BUFX2_insert379 (
    .A(_5762__hier0_bF$buf2),
    .Y(_5762__bF$buf27)
);

BUFX2 BUFX2_insert378 (
    .A(_5762__hier0_bF$buf1),
    .Y(_5762__bF$buf28)
);

BUFX2 BUFX2_insert377 (
    .A(_5762__hier0_bF$buf0),
    .Y(_5762__bF$buf29)
);

BUFX2 BUFX2_insert376 (
    .A(_5762__hier0_bF$buf5),
    .Y(_5762__bF$buf30)
);

BUFX2 BUFX2_insert375 (
    .A(_5762__hier0_bF$buf4),
    .Y(_5762__bF$buf31)
);

BUFX2 BUFX2_insert374 (
    .A(_5762__hier0_bF$buf3),
    .Y(_5762__bF$buf32)
);

BUFX2 BUFX2_insert373 (
    .A(_5762__hier0_bF$buf2),
    .Y(_5762__bF$buf33)
);

BUFX2 BUFX2_insert372 (
    .A(_5762__hier0_bF$buf1),
    .Y(_5762__bF$buf34)
);

BUFX2 BUFX2_insert371 (
    .A(_5762__hier0_bF$buf0),
    .Y(_5762__bF$buf35)
);

BUFX2 BUFX2_insert370 (
    .A(_5762__hier0_bF$buf5),
    .Y(_5762__bF$buf36)
);

BUFX2 BUFX2_insert369 (
    .A(_5762__hier0_bF$buf4),
    .Y(_5762__bF$buf37)
);

BUFX2 BUFX2_insert368 (
    .A(_5762__hier0_bF$buf3),
    .Y(_5762__bF$buf38)
);

BUFX2 BUFX2_insert367 (
    .A(_5762__hier0_bF$buf2),
    .Y(_5762__bF$buf39)
);

BUFX2 BUFX2_insert366 (
    .A(_5762__hier0_bF$buf1),
    .Y(_5762__bF$buf40)
);

BUFX2 BUFX2_insert365 (
    .A(_5762__hier0_bF$buf0),
    .Y(_5762__bF$buf41)
);

BUFX2 BUFX2_insert364 (
    .A(_5762__hier0_bF$buf5),
    .Y(_5762__bF$buf42)
);

BUFX2 BUFX2_insert363 (
    .A(_5762__hier0_bF$buf4),
    .Y(_5762__bF$buf43)
);

BUFX2 BUFX2_insert362 (
    .A(_5762__hier0_bF$buf3),
    .Y(_5762__bF$buf44)
);

BUFX2 BUFX2_insert361 (
    .A(_5762__hier0_bF$buf2),
    .Y(_5762__bF$buf45)
);

BUFX2 BUFX2_insert360 (
    .A(_5762__hier0_bF$buf1),
    .Y(_5762__bF$buf46)
);

BUFX2 BUFX2_insert359 (
    .A(_5762__hier0_bF$buf0),
    .Y(_5762__bF$buf47)
);

BUFX2 BUFX2_insert358 (
    .A(_4786_),
    .Y(_4786__bF$buf0)
);

BUFX2 BUFX2_insert357 (
    .A(_4786_),
    .Y(_4786__bF$buf1)
);

BUFX2 BUFX2_insert356 (
    .A(_4786_),
    .Y(_4786__bF$buf2)
);

BUFX2 BUFX2_insert355 (
    .A(_4786_),
    .Y(_4786__bF$buf3)
);

BUFX2 BUFX2_insert354 (
    .A(_4786_),
    .Y(_4786__bF$buf4)
);

BUFX2 BUFX2_insert353 (
    .A(_5477_),
    .Y(_5477__bF$buf0)
);

BUFX2 BUFX2_insert352 (
    .A(_5477_),
    .Y(_5477__bF$buf1)
);

BUFX2 BUFX2_insert351 (
    .A(_5477_),
    .Y(_5477__bF$buf2)
);

BUFX2 BUFX2_insert350 (
    .A(_5477_),
    .Y(_5477__bF$buf3)
);

BUFX2 BUFX2_insert349 (
    .A(_5477_),
    .Y(_5477__bF$buf4)
);

BUFX2 BUFX2_insert348 (
    .A(_5477_),
    .Y(_5477__bF$buf5)
);

BUFX2 BUFX2_insert347 (
    .A(_5477_),
    .Y(_5477__bF$buf6)
);

BUFX2 BUFX2_insert346 (
    .A(_5477_),
    .Y(_5477__bF$buf7)
);

BUFX2 BUFX2_insert345 (
    .A(_4845_),
    .Y(_4845__bF$buf0)
);

BUFX2 BUFX2_insert344 (
    .A(_4845_),
    .Y(_4845__bF$buf1)
);

BUFX2 BUFX2_insert343 (
    .A(_4845_),
    .Y(_4845__bF$buf2)
);

BUFX2 BUFX2_insert342 (
    .A(_4845_),
    .Y(_4845__bF$buf3)
);

BUFX2 BUFX2_insert341 (
    .A(_4845_),
    .Y(_4845__bF$buf4)
);

BUFX2 BUFX2_insert340 (
    .A(_4807_),
    .Y(_4807__bF$buf0)
);

BUFX2 BUFX2_insert339 (
    .A(_4807_),
    .Y(_4807__bF$buf1)
);

BUFX2 BUFX2_insert338 (
    .A(_4807_),
    .Y(_4807__bF$buf2)
);

BUFX2 BUFX2_insert337 (
    .A(_4807_),
    .Y(_4807__bF$buf3)
);

BUFX2 BUFX2_insert336 (
    .A(_4807_),
    .Y(_4807__bF$buf4)
);

BUFX2 BUFX2_insert335 (
    .A(_5442_),
    .Y(_5442__bF$buf0)
);

BUFX2 BUFX2_insert334 (
    .A(_5442_),
    .Y(_5442__bF$buf1)
);

BUFX2 BUFX2_insert333 (
    .A(_5442_),
    .Y(_5442__bF$buf2)
);

BUFX2 BUFX2_insert332 (
    .A(_5442_),
    .Y(_5442__bF$buf3)
);

BUFX2 BUFX2_insert331 (
    .A(_5442_),
    .Y(_5442__bF$buf4)
);

BUFX2 BUFX2_insert330 (
    .A(_5442_),
    .Y(_5442__bF$buf5)
);

BUFX2 BUFX2_insert329 (
    .A(_5442_),
    .Y(_5442__bF$buf6)
);

BUFX2 BUFX2_insert328 (
    .A(_5442_),
    .Y(_5442__bF$buf7)
);

BUFX2 BUFX2_insert327 (
    .A(_1841_),
    .Y(_1841__bF$buf0)
);

BUFX2 BUFX2_insert326 (
    .A(_1841_),
    .Y(_1841__bF$buf1)
);

BUFX2 BUFX2_insert325 (
    .A(_1841_),
    .Y(_1841__bF$buf2)
);

BUFX2 BUFX2_insert324 (
    .A(_1841_),
    .Y(_1841__bF$buf3)
);

BUFX2 BUFX2_insert323 (
    .A(_1841_),
    .Y(_1841__bF$buf4)
);

BUFX2 BUFX2_insert322 (
    .A(_1841_),
    .Y(_1841__bF$buf5)
);

BUFX2 BUFX2_insert321 (
    .A(_1841_),
    .Y(_1841__bF$buf6)
);

BUFX2 BUFX2_insert320 (
    .A(_1841_),
    .Y(_1841__bF$buf7)
);

BUFX2 BUFX2_insert319 (
    .A(_4851_),
    .Y(_4851__bF$buf0)
);

BUFX2 BUFX2_insert318 (
    .A(_4851_),
    .Y(_4851__bF$buf1)
);

BUFX2 BUFX2_insert317 (
    .A(_4851_),
    .Y(_4851__bF$buf2)
);

BUFX2 BUFX2_insert316 (
    .A(_4851_),
    .Y(_4851__bF$buf3)
);

BUFX2 BUFX2_insert315 (
    .A(_4851_),
    .Y(_4851__bF$buf4)
);

BUFX2 BUFX2_insert314 (
    .A(_182_),
    .Y(_182__bF$buf0)
);

BUFX2 BUFX2_insert313 (
    .A(_182_),
    .Y(_182__bF$buf1)
);

BUFX2 BUFX2_insert312 (
    .A(_182_),
    .Y(_182__bF$buf2)
);

BUFX2 BUFX2_insert311 (
    .A(_182_),
    .Y(_182__bF$buf3)
);

BUFX2 BUFX2_insert310 (
    .A(_182_),
    .Y(_182__bF$buf4)
);

BUFX2 BUFX2_insert309 (
    .A(_4813_),
    .Y(_4813__bF$buf0)
);

BUFX2 BUFX2_insert308 (
    .A(_4813_),
    .Y(_4813__bF$buf1)
);

BUFX2 BUFX2_insert307 (
    .A(_4813_),
    .Y(_4813__bF$buf2)
);

BUFX2 BUFX2_insert306 (
    .A(_4813_),
    .Y(_4813__bF$buf3)
);

BUFX2 BUFX2_insert305 (
    .A(_4813_),
    .Y(_4813__bF$buf4)
);

BUFX2 BUFX2_insert304 (
    .A(_3132_),
    .Y(_3132__bF$buf0)
);

BUFX2 BUFX2_insert303 (
    .A(_3132_),
    .Y(_3132__bF$buf1)
);

BUFX2 BUFX2_insert302 (
    .A(_3132_),
    .Y(_3132__bF$buf2)
);

BUFX2 BUFX2_insert301 (
    .A(_3132_),
    .Y(_3132__bF$buf3)
);

BUFX2 BUFX2_insert300 (
    .A(_3132_),
    .Y(_3132__bF$buf4)
);

BUFX2 BUFX2_insert299 (
    .A(_3132_),
    .Y(_3132__bF$buf5)
);

BUFX2 BUFX2_insert298 (
    .A(\datapath.idinstr_15_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_15_bF$buf0 )
);

BUFX2 BUFX2_insert297 (
    .A(\datapath.idinstr_15_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_15_bF$buf1 )
);

BUFX2 BUFX2_insert296 (
    .A(\datapath.idinstr_15_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_15_bF$buf2 )
);

BUFX2 BUFX2_insert295 (
    .A(\datapath.idinstr_15_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_15_bF$buf3 )
);

BUFX2 BUFX2_insert294 (
    .A(\datapath.idinstr_15_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_15_bF$buf4 )
);

BUFX2 BUFX2_insert293 (
    .A(\datapath.idinstr_15_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_15_bF$buf5 )
);

BUFX2 BUFX2_insert292 (
    .A(\datapath.idinstr_15_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_15_bF$buf6 )
);

BUFX2 BUFX2_insert291 (
    .A(\datapath.idinstr_15_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_15_bF$buf7 )
);

BUFX2 BUFX2_insert290 (
    .A(\datapath.idinstr_15_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_15_bF$buf8 )
);

BUFX2 BUFX2_insert289 (
    .A(\datapath.idinstr_15_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_15_bF$buf9 )
);

BUFX2 BUFX2_insert288 (
    .A(\datapath.idinstr_15_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_15_bF$buf10 )
);

BUFX2 BUFX2_insert287 (
    .A(\datapath.idinstr_15_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_15_bF$buf11 )
);

BUFX2 BUFX2_insert286 (
    .A(\datapath.idinstr_15_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_15_bF$buf12 )
);

BUFX2 BUFX2_insert285 (
    .A(\datapath.idinstr_15_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_15_bF$buf13 )
);

BUFX2 BUFX2_insert284 (
    .A(\datapath.idinstr_15_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_15_bF$buf14 )
);

BUFX2 BUFX2_insert283 (
    .A(\datapath.idinstr_15_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_15_bF$buf15 )
);

BUFX2 BUFX2_insert282 (
    .A(\datapath.idinstr_15_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_15_bF$buf16 )
);

BUFX2 BUFX2_insert281 (
    .A(\datapath.idinstr_15_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_15_bF$buf17 )
);

BUFX2 BUFX2_insert280 (
    .A(\datapath.idinstr_15_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_15_bF$buf18 )
);

BUFX2 BUFX2_insert279 (
    .A(\datapath.idinstr_15_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_15_bF$buf19 )
);

BUFX2 BUFX2_insert278 (
    .A(\datapath.idinstr_15_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_15_bF$buf20 )
);

BUFX2 BUFX2_insert277 (
    .A(\datapath.idinstr_15_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_15_bF$buf21 )
);

BUFX2 BUFX2_insert276 (
    .A(\datapath.idinstr_15_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_15_bF$buf22 )
);

BUFX2 BUFX2_insert275 (
    .A(\datapath.idinstr_15_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_15_bF$buf23 )
);

BUFX2 BUFX2_insert274 (
    .A(\datapath.idinstr_15_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_15_bF$buf24 )
);

BUFX2 BUFX2_insert273 (
    .A(\datapath.idinstr_15_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_15_bF$buf25 )
);

BUFX2 BUFX2_insert272 (
    .A(\datapath.idinstr_15_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_15_bF$buf26 )
);

BUFX2 BUFX2_insert271 (
    .A(\datapath.idinstr_15_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_15_bF$buf27 )
);

BUFX2 BUFX2_insert270 (
    .A(\datapath.idinstr_15_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_15_bF$buf28 )
);

BUFX2 BUFX2_insert269 (
    .A(\datapath.idinstr_15_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_15_bF$buf29 )
);

BUFX2 BUFX2_insert268 (
    .A(\datapath.idinstr_15_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_15_bF$buf30 )
);

BUFX2 BUFX2_insert267 (
    .A(\datapath.idinstr_15_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_15_bF$buf31 )
);

BUFX2 BUFX2_insert266 (
    .A(\datapath.idinstr_15_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_15_bF$buf32 )
);

BUFX2 BUFX2_insert265 (
    .A(\datapath.idinstr_15_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_15_bF$buf33 )
);

BUFX2 BUFX2_insert264 (
    .A(\datapath.idinstr_15_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_15_bF$buf34 )
);

BUFX2 BUFX2_insert263 (
    .A(\datapath.idinstr_15_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_15_bF$buf35 )
);

BUFX2 BUFX2_insert262 (
    .A(\datapath.idinstr_15_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_15_bF$buf36 )
);

BUFX2 BUFX2_insert261 (
    .A(\datapath.idinstr_15_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_15_bF$buf37 )
);

BUFX2 BUFX2_insert260 (
    .A(\datapath.idinstr_15_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_15_bF$buf38 )
);

BUFX2 BUFX2_insert259 (
    .A(\datapath.idinstr_15_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_15_bF$buf39 )
);

BUFX2 BUFX2_insert258 (
    .A(\datapath.idinstr_15_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_15_bF$buf40 )
);

BUFX2 BUFX2_insert257 (
    .A(\datapath.idinstr_15_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_15_bF$buf41 )
);

BUFX2 BUFX2_insert256 (
    .A(\datapath.idinstr_15_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_15_bF$buf42 )
);

BUFX2 BUFX2_insert255 (
    .A(\datapath.idinstr_15_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_15_bF$buf43 )
);

BUFX2 BUFX2_insert254 (
    .A(\datapath.idinstr_15_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_15_bF$buf44 )
);

BUFX2 BUFX2_insert253 (
    .A(\datapath.idinstr_15_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_15_bF$buf45 )
);

BUFX2 BUFX2_insert252 (
    .A(\datapath.idinstr_15_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_15_bF$buf46 )
);

BUFX2 BUFX2_insert251 (
    .A(\datapath.idinstr_15_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_15_bF$buf47 )
);

BUFX2 BUFX2_insert250 (
    .A(\datapath.idinstr_15_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_15_bF$buf48 )
);

BUFX2 BUFX2_insert249 (
    .A(\datapath.idinstr_15_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_15_bF$buf49 )
);

BUFX2 BUFX2_insert248 (
    .A(\datapath.idinstr_15_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_15_bF$buf50 )
);

BUFX2 BUFX2_insert247 (
    .A(\datapath.idinstr_15_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_15_bF$buf51 )
);

BUFX2 BUFX2_insert246 (
    .A(\datapath.idinstr_15_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_15_bF$buf52 )
);

BUFX2 BUFX2_insert245 (
    .A(\datapath.idinstr_15_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_15_bF$buf53 )
);

BUFX2 BUFX2_insert244 (
    .A(\datapath.idinstr_15_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_15_bF$buf54 )
);

BUFX2 BUFX2_insert243 (
    .A(_2767_),
    .Y(_2767__bF$buf0)
);

BUFX2 BUFX2_insert242 (
    .A(_2767_),
    .Y(_2767__bF$buf1)
);

BUFX2 BUFX2_insert241 (
    .A(_2767_),
    .Y(_2767__bF$buf2)
);

BUFX2 BUFX2_insert240 (
    .A(_2767_),
    .Y(_2767__bF$buf3)
);

BUFX2 BUFX2_insert239 (
    .A(_2767_),
    .Y(_2767__bF$buf4)
);

BUFX2 BUFX2_insert238 (
    .A(_2118_),
    .Y(_2118__bF$buf0)
);

BUFX2 BUFX2_insert237 (
    .A(_2118_),
    .Y(_2118__bF$buf1)
);

BUFX2 BUFX2_insert236 (
    .A(_2118_),
    .Y(_2118__bF$buf2)
);

BUFX2 BUFX2_insert235 (
    .A(_2118_),
    .Y(_2118__bF$buf3)
);

BUFX2 BUFX2_insert234 (
    .A(_5510_),
    .Y(_5510__bF$buf0)
);

BUFX2 BUFX2_insert233 (
    .A(_5510_),
    .Y(_5510__bF$buf1)
);

BUFX2 BUFX2_insert232 (
    .A(_5510_),
    .Y(_5510__bF$buf2)
);

BUFX2 BUFX2_insert231 (
    .A(_5510_),
    .Y(_5510__bF$buf3)
);

BUFX2 BUFX2_insert230 (
    .A(_5510_),
    .Y(_5510__bF$buf4)
);

BUFX2 BUFX2_insert229 (
    .A(_5510_),
    .Y(_5510__bF$buf5)
);

BUFX2 BUFX2_insert228 (
    .A(_5510_),
    .Y(_5510__bF$buf6)
);

BUFX2 BUFX2_insert227 (
    .A(_5510_),
    .Y(_5510__bF$buf7)
);

BUFX2 BUFX2_insert226 (
    .A(\datapath.idinstr [18]),
    .Y(\datapath.idinstr_18_bF$buf0 )
);

BUFX2 BUFX2_insert225 (
    .A(\datapath.idinstr [18]),
    .Y(\datapath.idinstr_18_bF$buf1 )
);

BUFX2 BUFX2_insert224 (
    .A(\datapath.idinstr [18]),
    .Y(\datapath.idinstr_18_bF$buf2 )
);

BUFX2 BUFX2_insert223 (
    .A(\datapath.idinstr [18]),
    .Y(\datapath.idinstr_18_bF$buf3 )
);

BUFX2 BUFX2_insert222 (
    .A(\datapath.idinstr [18]),
    .Y(\datapath.idinstr_18_bF$buf4 )
);

BUFX2 BUFX2_insert221 (
    .A(\datapath.idinstr [18]),
    .Y(\datapath.idinstr_18_bF$buf5 )
);

BUFX2 BUFX2_insert220 (
    .A(\datapath.idinstr [18]),
    .Y(\datapath.idinstr_18_bF$buf6 )
);

BUFX2 BUFX2_insert219 (
    .A(_4857_),
    .Y(_4857__bF$buf0)
);

BUFX2 BUFX2_insert218 (
    .A(_4857_),
    .Y(_4857__bF$buf1)
);

BUFX2 BUFX2_insert217 (
    .A(_4857_),
    .Y(_4857__bF$buf2)
);

BUFX2 BUFX2_insert216 (
    .A(_4857_),
    .Y(_4857__bF$buf3)
);

BUFX2 BUFX2_insert215 (
    .A(_4857_),
    .Y(_4857__bF$buf4)
);

BUFX2 BUFX2_insert214 (
    .A(_5586_),
    .Y(_5586__bF$buf0)
);

BUFX2 BUFX2_insert213 (
    .A(_5586_),
    .Y(_5586__bF$buf1)
);

BUFX2 BUFX2_insert212 (
    .A(_5586_),
    .Y(_5586__bF$buf2)
);

BUFX2 BUFX2_insert211 (
    .A(_5586_),
    .Y(_5586__bF$buf3)
);

BUFX2 BUFX2_insert210 (
    .A(_5586_),
    .Y(_5586__bF$buf4)
);

BUFX2 BUFX2_insert209 (
    .A(_4819_),
    .Y(_4819__bF$buf0)
);

BUFX2 BUFX2_insert208 (
    .A(_4819_),
    .Y(_4819__bF$buf1)
);

BUFX2 BUFX2_insert207 (
    .A(_4819_),
    .Y(_4819__bF$buf2)
);

BUFX2 BUFX2_insert206 (
    .A(_4819_),
    .Y(_4819__bF$buf3)
);

BUFX2 BUFX2_insert205 (
    .A(_4819_),
    .Y(_4819__bF$buf4)
);

BUFX2 BUFX2_insert204 (
    .A(\datapath.idinstr_21_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_21_bF$buf0 )
);

BUFX2 BUFX2_insert203 (
    .A(\datapath.idinstr_21_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_21_bF$buf1 )
);

BUFX2 BUFX2_insert202 (
    .A(\datapath.idinstr_21_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_21_bF$buf2 )
);

BUFX2 BUFX2_insert201 (
    .A(\datapath.idinstr_21_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_21_bF$buf3 )
);

BUFX2 BUFX2_insert200 (
    .A(\datapath.idinstr_21_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_21_bF$buf4 )
);

BUFX2 BUFX2_insert199 (
    .A(\datapath.idinstr_21_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_21_bF$buf5 )
);

BUFX2 BUFX2_insert198 (
    .A(\datapath.idinstr_21_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_21_bF$buf6 )
);

BUFX2 BUFX2_insert197 (
    .A(\datapath.idinstr_21_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_21_bF$buf7 )
);

BUFX2 BUFX2_insert196 (
    .A(\datapath.idinstr_21_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_21_bF$buf8 )
);

BUFX2 BUFX2_insert195 (
    .A(\datapath.idinstr_21_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_21_bF$buf9 )
);

BUFX2 BUFX2_insert194 (
    .A(\datapath.idinstr_21_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_21_bF$buf10 )
);

BUFX2 BUFX2_insert193 (
    .A(\datapath.idinstr_21_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_21_bF$buf11 )
);

BUFX2 BUFX2_insert192 (
    .A(\datapath.idinstr_21_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_21_bF$buf12 )
);

BUFX2 BUFX2_insert191 (
    .A(\datapath.idinstr_21_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_21_bF$buf13 )
);

BUFX2 BUFX2_insert190 (
    .A(\datapath.idinstr_21_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_21_bF$buf14 )
);

BUFX2 BUFX2_insert189 (
    .A(\datapath.idinstr_21_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_21_bF$buf15 )
);

BUFX2 BUFX2_insert188 (
    .A(\datapath.idinstr_21_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_21_bF$buf16 )
);

BUFX2 BUFX2_insert187 (
    .A(\datapath.idinstr_21_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_21_bF$buf17 )
);

BUFX2 BUFX2_insert186 (
    .A(\datapath.idinstr_21_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_21_bF$buf18 )
);

BUFX2 BUFX2_insert185 (
    .A(\datapath.idinstr_21_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_21_bF$buf19 )
);

BUFX2 BUFX2_insert184 (
    .A(\datapath.idinstr_21_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_21_bF$buf20 )
);

BUFX2 BUFX2_insert183 (
    .A(\datapath.idinstr_21_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_21_bF$buf21 )
);

BUFX2 BUFX2_insert182 (
    .A(\datapath.idinstr_21_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_21_bF$buf22 )
);

BUFX2 BUFX2_insert181 (
    .A(\datapath.idinstr_21_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_21_bF$buf23 )
);

BUFX2 BUFX2_insert180 (
    .A(\datapath.idinstr_21_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_21_bF$buf24 )
);

BUFX2 BUFX2_insert179 (
    .A(\datapath.idinstr_21_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_21_bF$buf25 )
);

BUFX2 BUFX2_insert178 (
    .A(\datapath.idinstr_21_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_21_bF$buf26 )
);

BUFX2 BUFX2_insert177 (
    .A(\datapath.idinstr_21_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_21_bF$buf27 )
);

BUFX2 BUFX2_insert176 (
    .A(\datapath.idinstr_21_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_21_bF$buf28 )
);

BUFX2 BUFX2_insert175 (
    .A(\datapath.idinstr_21_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_21_bF$buf29 )
);

BUFX2 BUFX2_insert174 (
    .A(\datapath.idinstr_21_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_21_bF$buf30 )
);

BUFX2 BUFX2_insert173 (
    .A(\datapath.idinstr_21_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_21_bF$buf31 )
);

BUFX2 BUFX2_insert172 (
    .A(\datapath.idinstr_21_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_21_bF$buf32 )
);

BUFX2 BUFX2_insert171 (
    .A(\datapath.idinstr_21_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_21_bF$buf33 )
);

BUFX2 BUFX2_insert170 (
    .A(\datapath.idinstr_21_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_21_bF$buf34 )
);

BUFX2 BUFX2_insert169 (
    .A(\datapath.idinstr_21_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_21_bF$buf35 )
);

BUFX2 BUFX2_insert168 (
    .A(\datapath.idinstr_21_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_21_bF$buf36 )
);

BUFX2 BUFX2_insert167 (
    .A(\datapath.idinstr_21_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_21_bF$buf37 )
);

BUFX2 BUFX2_insert166 (
    .A(\datapath.idinstr_21_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_21_bF$buf38 )
);

BUFX2 BUFX2_insert165 (
    .A(\datapath.idinstr_21_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_21_bF$buf39 )
);

BUFX2 BUFX2_insert164 (
    .A(\datapath.idinstr_21_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_21_bF$buf40 )
);

BUFX2 BUFX2_insert163 (
    .A(\datapath.idinstr_21_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_21_bF$buf41 )
);

BUFX2 BUFX2_insert162 (
    .A(\datapath.idinstr_21_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_21_bF$buf42 )
);

BUFX2 BUFX2_insert161 (
    .A(\datapath.idinstr_21_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_21_bF$buf43 )
);

BUFX2 BUFX2_insert160 (
    .A(\datapath.idinstr_21_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_21_bF$buf44 )
);

BUFX2 BUFX2_insert159 (
    .A(\datapath.idinstr_21_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_21_bF$buf45 )
);

BUFX2 BUFX2_insert158 (
    .A(\datapath.idinstr_21_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_21_bF$buf46 )
);

BUFX2 BUFX2_insert157 (
    .A(\datapath.idinstr_21_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_21_bF$buf47 )
);

BUFX2 BUFX2_insert156 (
    .A(\datapath.idinstr_21_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_21_bF$buf48 )
);

BUFX2 BUFX2_insert155 (
    .A(\datapath.idinstr_21_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_21_bF$buf49 )
);

BUFX2 BUFX2_insert154 (
    .A(\datapath.idinstr_21_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_21_bF$buf50 )
);

BUFX2 BUFX2_insert153 (
    .A(\datapath.idinstr_21_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_21_bF$buf51 )
);

BUFX2 BUFX2_insert152 (
    .A(_5551_),
    .Y(_5551__bF$buf0)
);

BUFX2 BUFX2_insert151 (
    .A(_5551_),
    .Y(_5551__bF$buf1)
);

BUFX2 BUFX2_insert150 (
    .A(_5551_),
    .Y(_5551__bF$buf2)
);

BUFX2 BUFX2_insert149 (
    .A(_5551_),
    .Y(_5551__bF$buf3)
);

BUFX2 BUFX2_insert148 (
    .A(_5551_),
    .Y(_5551__bF$buf4)
);

BUFX2 BUFX2_insert147 (
    .A(_5551_),
    .Y(_5551__bF$buf5)
);

BUFX2 BUFX2_insert146 (
    .A(_5551_),
    .Y(_5551__bF$buf6)
);

BUFX2 BUFX2_insert145 (
    .A(_5551_),
    .Y(_5551__bF$buf7)
);

BUFX2 BUFX2_insert144 (
    .A(_2027_),
    .Y(_2027__bF$buf0)
);

BUFX2 BUFX2_insert143 (
    .A(_2027_),
    .Y(_2027__bF$buf1)
);

BUFX2 BUFX2_insert142 (
    .A(_2027_),
    .Y(_2027__bF$buf2)
);

BUFX2 BUFX2_insert141 (
    .A(_2027_),
    .Y(_2027__bF$buf3)
);

BUFX2 BUFX2_insert140 (
    .A(_3138_),
    .Y(_3138__bF$buf0)
);

BUFX2 BUFX2_insert139 (
    .A(_3138_),
    .Y(_3138__bF$buf1)
);

BUFX2 BUFX2_insert138 (
    .A(_3138_),
    .Y(_3138__bF$buf2)
);

BUFX2 BUFX2_insert137 (
    .A(_3138_),
    .Y(_3138__bF$buf3)
);

BUFX2 BUFX2_insert136 (
    .A(_3138_),
    .Y(_3138__bF$buf4)
);

BUFX2 BUFX2_insert135 (
    .A(_3138_),
    .Y(_3138__bF$buf5)
);

BUFX2 BUFX2_insert134 (
    .A(_3138_),
    .Y(_3138__bF$buf6)
);

BUFX2 BUFX2_insert133 (
    .A(_3558_),
    .Y(_3558__bF$buf0)
);

BUFX2 BUFX2_insert132 (
    .A(_3558_),
    .Y(_3558__bF$buf1)
);

BUFX2 BUFX2_insert131 (
    .A(_3558_),
    .Y(_3558__bF$buf2)
);

BUFX2 BUFX2_insert130 (
    .A(_3558_),
    .Y(_3558__bF$buf3)
);

BUFX2 BUFX2_insert129 (
    .A(_3558_),
    .Y(_3558__bF$buf4)
);

BUFX2 BUFX2_insert128 (
    .A(_9058_),
    .Y(_9058__bF$buf0)
);

BUFX2 BUFX2_insert127 (
    .A(_9058_),
    .Y(_9058__bF$buf1)
);

BUFX2 BUFX2_insert126 (
    .A(_9058_),
    .Y(_9058__bF$buf2)
);

BUFX2 BUFX2_insert125 (
    .A(_9058_),
    .Y(_9058__bF$buf3)
);

BUFX2 BUFX2_insert124 (
    .A(_9058_),
    .Y(_9058__bF$buf4)
);

BUFX2 BUFX2_insert123 (
    .A(_9058_),
    .Y(_9058__bF$buf5)
);

BUFX2 BUFX2_insert122 (
    .A(_9058_),
    .Y(_9058__bF$buf6)
);

BUFX2 BUFX2_insert121 (
    .A(_9058_),
    .Y(_9058__bF$buf7)
);

BUFX2 BUFX2_insert120 (
    .A(_2870_),
    .Y(_2870__bF$buf0)
);

BUFX2 BUFX2_insert119 (
    .A(_2870_),
    .Y(_2870__bF$buf1)
);

BUFX2 BUFX2_insert118 (
    .A(_2870_),
    .Y(_2870__bF$buf2)
);

BUFX2 BUFX2_insert117 (
    .A(_2870_),
    .Y(_2870__bF$buf3)
);

BUFX2 BUFX2_insert116 (
    .A(_2870_),
    .Y(_2870__bF$buf4)
);

BUFX2 BUFX2_insert115 (
    .A(_2870_),
    .Y(_2870__bF$buf5)
);

BUFX2 BUFX2_insert114 (
    .A(_2870_),
    .Y(_2870__bF$buf6)
);

BUFX2 BUFX2_insert113 (
    .A(_3561_),
    .Y(_3561__bF$buf0)
);

BUFX2 BUFX2_insert112 (
    .A(_3561_),
    .Y(_3561__bF$buf1)
);

BUFX2 BUFX2_insert111 (
    .A(_3561_),
    .Y(_3561__bF$buf2)
);

BUFX2 BUFX2_insert110 (
    .A(_3561_),
    .Y(_3561__bF$buf3)
);

BUFX2 BUFX2_insert109 (
    .A(_3561_),
    .Y(_3561__bF$buf4)
);

BUFX2 BUFX2_insert108 (
    .A(\datapath.idinstr [24]),
    .Y(\datapath.idinstr_24_bF$buf0 )
);

BUFX2 BUFX2_insert107 (
    .A(\datapath.idinstr [24]),
    .Y(\datapath.idinstr_24_bF$buf1 )
);

BUFX2 BUFX2_insert106 (
    .A(\datapath.idinstr [24]),
    .Y(\datapath.idinstr_24_bF$buf2 )
);

BUFX2 BUFX2_insert105 (
    .A(\datapath.idinstr [24]),
    .Y(\datapath.idinstr_24_bF$buf3 )
);

BUFX2 BUFX2_insert104 (
    .A(\datapath.idinstr [24]),
    .Y(\datapath.idinstr_24_bF$buf4 )
);

BUFX2 BUFX2_insert103 (
    .A(\datapath.idinstr [24]),
    .Y(\datapath.idinstr_24_bF$buf5 )
);

BUFX2 BUFX2_insert102 (
    .A(_288_),
    .Y(_288__bF$buf0)
);

BUFX2 BUFX2_insert101 (
    .A(_288_),
    .Y(_288__bF$buf1)
);

BUFX2 BUFX2_insert100 (
    .A(_288_),
    .Y(_288__bF$buf2)
);

BUFX2 BUFX2_insert99 (
    .A(_288_),
    .Y(_288__bF$buf3)
);

BUFX2 BUFX2_insert98 (
    .A(_288_),
    .Y(_288__bF$buf4)
);

BUFX2 BUFX2_insert97 (
    .A(_4863_),
    .Y(_4863__bF$buf0)
);

BUFX2 BUFX2_insert96 (
    .A(_4863_),
    .Y(_4863__bF$buf1)
);

BUFX2 BUFX2_insert95 (
    .A(_4863_),
    .Y(_4863__bF$buf2)
);

BUFX2 BUFX2_insert94 (
    .A(_4863_),
    .Y(_4863__bF$buf3)
);

BUFX2 BUFX2_insert93 (
    .A(_4863_),
    .Y(_4863__bF$buf4)
);

BUFX2 BUFX2_insert92 (
    .A(_4863_),
    .Y(_4863__bF$buf5)
);

BUFX2 BUFX2_insert91 (
    .A(_4863_),
    .Y(_4863__bF$buf6)
);

BUFX2 BUFX2_insert90 (
    .A(_4863_),
    .Y(_4863__bF$buf7)
);

BUFX2 BUFX2_insert89 (
    .A(_4825_),
    .Y(_4825__bF$buf0)
);

BUFX2 BUFX2_insert88 (
    .A(_4825_),
    .Y(_4825__bF$buf1)
);

BUFX2 BUFX2_insert87 (
    .A(_4825_),
    .Y(_4825__bF$buf2)
);

BUFX2 BUFX2_insert86 (
    .A(_4825_),
    .Y(_4825__bF$buf3)
);

BUFX2 BUFX2_insert85 (
    .A(_4825_),
    .Y(_4825__bF$buf4)
);

BUFX2 BUFX2_insert84 (
    .A(_9158_),
    .Y(_9158__bF$buf0)
);

BUFX2 BUFX2_insert83 (
    .A(_9158_),
    .Y(_9158__bF$buf1)
);

BUFX2 BUFX2_insert82 (
    .A(_9158_),
    .Y(_9158__bF$buf2)
);

BUFX2 BUFX2_insert81 (
    .A(_9158_),
    .Y(_9158__bF$buf3)
);

BUFX2 BUFX2_insert80 (
    .A(_9158_),
    .Y(_9158__bF$buf4)
);

BUFX2 BUFX2_insert79 (
    .A(_5689_),
    .Y(_5689__bF$buf0)
);

BUFX2 BUFX2_insert78 (
    .A(_5689_),
    .Y(_5689__bF$buf1)
);

BUFX2 BUFX2_insert77 (
    .A(_5689_),
    .Y(_5689__bF$buf2)
);

BUFX2 BUFX2_insert76 (
    .A(_5689_),
    .Y(_5689__bF$buf3)
);

BUFX2 BUFX2_insert75 (
    .A(_5689_),
    .Y(_5689__bF$buf4)
);

BUFX2 BUFX2_insert74 (
    .A(_388_),
    .Y(_388__bF$buf0)
);

BUFX2 BUFX2_insert73 (
    .A(_388_),
    .Y(_388__bF$buf1)
);

BUFX2 BUFX2_insert72 (
    .A(_388_),
    .Y(_388__bF$buf2)
);

BUFX2 BUFX2_insert71 (
    .A(_388_),
    .Y(_388__bF$buf3)
);

BUFX2 BUFX2_insert70 (
    .A(_388_),
    .Y(_388__bF$buf4)
);

BUFX2 BUFX2_insert69 (
    .A(_4831_),
    .Y(_4831__bF$buf0)
);

BUFX2 BUFX2_insert68 (
    .A(_4831_),
    .Y(_4831__bF$buf1)
);

BUFX2 BUFX2_insert67 (
    .A(_4831_),
    .Y(_4831__bF$buf2)
);

BUFX2 BUFX2_insert66 (
    .A(_4831_),
    .Y(_4831__bF$buf3)
);

BUFX2 BUFX2_insert65 (
    .A(_4831_),
    .Y(_4831__bF$buf4)
);

BUFX2 BUFX2_insert64 (
    .A(\controlunit.mret ),
    .Y(\controlunit.mret_bF$buf0 )
);

BUFX2 BUFX2_insert63 (
    .A(\controlunit.mret ),
    .Y(\controlunit.mret_bF$buf1 )
);

BUFX2 BUFX2_insert62 (
    .A(\controlunit.mret ),
    .Y(\controlunit.mret_bF$buf2 )
);

BUFX2 BUFX2_insert61 (
    .A(\controlunit.mret ),
    .Y(\controlunit.mret_bF$buf3 )
);

BUFX2 BUFX2_insert60 (
    .A(\controlunit.mret ),
    .Y(\controlunit.mret_bF$buf4 )
);

BUFX2 BUFX2_insert59 (
    .A(_1824_),
    .Y(_1824__bF$buf0)
);

BUFX2 BUFX2_insert58 (
    .A(_1824_),
    .Y(_1824__bF$buf1)
);

BUFX2 BUFX2_insert57 (
    .A(_1824_),
    .Y(_1824__bF$buf2)
);

BUFX2 BUFX2_insert56 (
    .A(_1824_),
    .Y(_1824__bF$buf3)
);

BUFX2 BUFX2_insert55 (
    .A(_1824_),
    .Y(_1824__bF$buf4)
);

BUFX2 BUFX2_insert54 (
    .A(_1824_),
    .Y(_1824__bF$buf5)
);

BUFX2 BUFX2_insert53 (
    .A(_2133_),
    .Y(_2133__bF$buf0)
);

BUFX2 BUFX2_insert52 (
    .A(_2133_),
    .Y(_2133__bF$buf1)
);

BUFX2 BUFX2_insert51 (
    .A(_2133_),
    .Y(_2133__bF$buf2)
);

BUFX2 BUFX2_insert50 (
    .A(_2133_),
    .Y(_2133__bF$buf3)
);

BUFX2 BUFX2_insert49 (
    .A(_7418_),
    .Y(_7418__bF$buf0)
);

BUFX2 BUFX2_insert48 (
    .A(_7418_),
    .Y(_7418__bF$buf1)
);

BUFX2 BUFX2_insert47 (
    .A(_7418_),
    .Y(_7418__bF$buf2)
);

BUFX2 BUFX2_insert46 (
    .A(_7418_),
    .Y(_7418__bF$buf3)
);

BUFX2 BUFX2_insert45 (
    .A(_7418_),
    .Y(_7418__bF$buf4)
);

BUFX2 BUFX2_insert44 (
    .A(_5789_),
    .Y(_5789__bF$buf0)
);

BUFX2 BUFX2_insert43 (
    .A(_5789_),
    .Y(_5789__bF$buf1)
);

BUFX2 BUFX2_insert42 (
    .A(_5789_),
    .Y(_5789__bF$buf2)
);

BUFX2 BUFX2_insert41 (
    .A(_5789_),
    .Y(_5789__bF$buf3)
);

BUFX2 BUFX2_insert40 (
    .A(_5789_),
    .Y(_5789__bF$buf4)
);

BUFX2 BUFX2_insert39 (
    .A(\datapath.alu.b [2]),
    .Y(\datapath.alu.b_2_bF$buf0 )
);

BUFX2 BUFX2_insert38 (
    .A(\datapath.alu.b [2]),
    .Y(\datapath.alu.b_2_bF$buf1 )
);

BUFX2 BUFX2_insert37 (
    .A(\datapath.alu.b [2]),
    .Y(\datapath.alu.b_2_bF$buf2 )
);

BUFX2 BUFX2_insert36 (
    .A(\datapath.alu.b [2]),
    .Y(\datapath.alu.b_2_bF$buf3 )
);

BUFX2 BUFX2_insert35 (
    .A(\datapath.alu.b [2]),
    .Y(\datapath.alu.b_2_bF$buf4 )
);

BUFX2 BUFX2_insert34 (
    .A(\datapath.alu.b [2]),
    .Y(\datapath.alu.b_2_bF$buf5 )
);

BUFX2 BUFX2_insert33 (
    .A(\datapath.alu.b [2]),
    .Y(\datapath.alu.b_2_bF$buf6 )
);

BUFX2 BUFX2_insert32 (
    .A(\datapath.alu.b [2]),
    .Y(\datapath.alu.b_2_bF$buf7 )
);

BUFX2 BUFX2_insert31 (
    .A(_4969_),
    .Y(_4969__bF$buf0)
);

BUFX2 BUFX2_insert30 (
    .A(_4969_),
    .Y(_4969__bF$buf1)
);

BUFX2 BUFX2_insert29 (
    .A(_4969_),
    .Y(_4969__bF$buf2)
);

BUFX2 BUFX2_insert28 (
    .A(_4969_),
    .Y(_4969__bF$buf3)
);

BUFX2 BUFX2_insert27 (
    .A(_4969_),
    .Y(_4969__bF$buf4)
);

BUFX2 BUFX2_insert26 (
    .A(_4969_),
    .Y(_4969__bF$buf5)
);

BUFX2 BUFX2_insert25 (
    .A(_4969_),
    .Y(_4969__bF$buf6)
);

BUFX2 BUFX2_insert24 (
    .A(_4969_),
    .Y(_4969__bF$buf7)
);

BUFX2 BUFX2_insert23 (
    .A(_5375_),
    .Y(_5375__bF$buf0)
);

BUFX2 BUFX2_insert22 (
    .A(_5375_),
    .Y(_5375__bF$buf1)
);

BUFX2 BUFX2_insert21 (
    .A(_5375_),
    .Y(_5375__bF$buf2)
);

BUFX2 BUFX2_insert20 (
    .A(_5375_),
    .Y(_5375__bF$buf3)
);

BUFX2 BUFX2_insert19 (
    .A(_5375_),
    .Y(_5375__bF$buf4)
);

BUFX2 BUFX2_insert18 (
    .A(_5375_),
    .Y(_5375__bF$buf5)
);

BUFX2 BUFX2_insert17 (
    .A(_5375_),
    .Y(_5375__bF$buf6)
);

BUFX2 BUFX2_insert16 (
    .A(_5375_),
    .Y(_5375__bF$buf7)
);

BUFX2 BUFX2_insert15 (
    .A(_4837_),
    .Y(_4837__bF$buf0)
);

BUFX2 BUFX2_insert14 (
    .A(_4837_),
    .Y(_4837__bF$buf1)
);

BUFX2 BUFX2_insert13 (
    .A(_4837_),
    .Y(_4837__bF$buf2)
);

BUFX2 BUFX2_insert12 (
    .A(_4837_),
    .Y(_4837__bF$buf3)
);

BUFX2 BUFX2_insert11 (
    .A(_4837_),
    .Y(_4837__bF$buf4)
);

BUFX2 BUFX2_insert10 (
    .A(_5757_),
    .Y(_5757__bF$buf0)
);

BUFX2 BUFX2_insert9 (
    .A(_5757_),
    .Y(_5757__bF$buf1)
);

BUFX2 BUFX2_insert8 (
    .A(_5757_),
    .Y(_5757__bF$buf2)
);

BUFX2 BUFX2_insert7 (
    .A(_5757_),
    .Y(_5757__bF$buf3)
);

BUFX2 BUFX2_insert6 (
    .A(_5757_),
    .Y(_5757__bF$buf4)
);

BUFX2 BUFX2_insert5 (
    .A(_5757_),
    .Y(_5757__bF$buf5)
);

BUFX2 BUFX2_insert4 (
    .A(_5757_),
    .Y(_5757__bF$buf6)
);

BUFX2 BUFX2_insert3 (
    .A(_5757_),
    .Y(_5757__bF$buf7)
);

BUFX2 BUFX2_insert2 (
    .A(_5757_),
    .Y(_5757__bF$buf8)
);

BUFX2 BUFX2_insert1 (
    .A(_5757_),
    .Y(_5757__bF$buf9)
);

BUFX2 BUFX2_insert0 (
    .A(_5757_),
    .Y(_5757__bF$buf10)
);

NAND2X1 _10000_ (
    .A(\datapath.registers.regb_data [31]),
    .B(_288__bF$buf4),
    .Y(_382_)
);

NAND2X1 _10001_ (
    .A(\datapath.immediatedecoder._12_ ),
    .B(_286__bF$buf4),
    .Y(_383_)
);

NAND2X1 _10002_ (
    .A(\datapath.csr.csr_data [31]),
    .B(_287__bF$buf4),
    .Y(_384_)
);

NAND3X1 _10003_ (
    .A(_383_),
    .B(_384_),
    .C(_382_),
    .Y(\datapath.muxbval [31])
);

INVX1 _10004_ (
    .A(asel[1]),
    .Y(_385_)
);

AND2X2 _10005_ (
    .A(_385_),
    .B(asel[0]),
    .Y(_386_)
);

NOR2X1 _10006_ (
    .A(asel[0]),
    .B(_385_),
    .Y(_387_)
);

NOR2X1 _10007_ (
    .A(_387__bF$buf4),
    .B(_386__bF$buf4),
    .Y(_388_)
);

NAND2X1 _10008_ (
    .A(\datapath.registers.rega_data [0]),
    .B(_388__bF$buf4),
    .Y(_389_)
);

NAND2X1 _10009_ (
    .A(\datapath.idpc [0]),
    .B(_386__bF$buf3),
    .Y(_390_)
);

NAND2X1 _10010_ (
    .A(\datapath.csr.csr_data [0]),
    .B(_387__bF$buf3),
    .Y(_391_)
);

NAND3X1 _10011_ (
    .A(_390_),
    .B(_391_),
    .C(_389_),
    .Y(\datapath.muxaval [0])
);

NAND2X1 _10012_ (
    .A(\datapath.registers.rega_data [1]),
    .B(_388__bF$buf3),
    .Y(_392_)
);

NAND2X1 _10013_ (
    .A(\datapath.idpc [1]),
    .B(_386__bF$buf2),
    .Y(_393_)
);

NAND2X1 _10014_ (
    .A(\datapath.csr.csr_data [1]),
    .B(_387__bF$buf2),
    .Y(_394_)
);

NAND3X1 _10015_ (
    .A(_393_),
    .B(_394_),
    .C(_392_),
    .Y(\datapath.muxaval [1])
);

NAND2X1 _10016_ (
    .A(\datapath.registers.rega_data [2]),
    .B(_388__bF$buf2),
    .Y(_395_)
);

NAND2X1 _10017_ (
    .A(\datapath.idpc [2]),
    .B(_386__bF$buf1),
    .Y(_396_)
);

NAND2X1 _10018_ (
    .A(\datapath.csr.csr_data [2]),
    .B(_387__bF$buf1),
    .Y(_397_)
);

NAND3X1 _10019_ (
    .A(_396_),
    .B(_397_),
    .C(_395_),
    .Y(\datapath.muxaval [2])
);

NAND2X1 _10020_ (
    .A(\datapath.registers.rega_data [3]),
    .B(_388__bF$buf1),
    .Y(_398_)
);

NAND2X1 _10021_ (
    .A(\datapath.idpc [3]),
    .B(_386__bF$buf0),
    .Y(_399_)
);

NAND2X1 _10022_ (
    .A(\datapath.csr.csr_data [3]),
    .B(_387__bF$buf0),
    .Y(_400_)
);

NAND3X1 _10023_ (
    .A(_399_),
    .B(_400_),
    .C(_398_),
    .Y(\datapath.muxaval [3])
);

NAND2X1 _10024_ (
    .A(\datapath.registers.rega_data [4]),
    .B(_388__bF$buf0),
    .Y(_401_)
);

NAND2X1 _10025_ (
    .A(\datapath.idpc [4]),
    .B(_386__bF$buf4),
    .Y(_402_)
);

NAND2X1 _10026_ (
    .A(\datapath.csr.csr_data [4]),
    .B(_387__bF$buf4),
    .Y(_403_)
);

NAND3X1 _10027_ (
    .A(_402_),
    .B(_403_),
    .C(_401_),
    .Y(\datapath.muxaval [4])
);

NAND2X1 _10028_ (
    .A(\datapath.registers.rega_data [5]),
    .B(_388__bF$buf4),
    .Y(_404_)
);

NAND2X1 _10029_ (
    .A(\datapath.idpc [5]),
    .B(_386__bF$buf3),
    .Y(_405_)
);

NAND2X1 _10030_ (
    .A(\datapath.csr.csr_data [5]),
    .B(_387__bF$buf3),
    .Y(_406_)
);

NAND3X1 _10031_ (
    .A(_405_),
    .B(_406_),
    .C(_404_),
    .Y(\datapath.muxaval [5])
);

NAND2X1 _10032_ (
    .A(\datapath.registers.rega_data [6]),
    .B(_388__bF$buf3),
    .Y(_407_)
);

NAND2X1 _10033_ (
    .A(\datapath.idpc [6]),
    .B(_386__bF$buf2),
    .Y(_408_)
);

NAND2X1 _10034_ (
    .A(\datapath.csr.csr_data [6]),
    .B(_387__bF$buf2),
    .Y(_409_)
);

NAND3X1 _10035_ (
    .A(_408_),
    .B(_409_),
    .C(_407_),
    .Y(\datapath.muxaval [6])
);

NAND2X1 _10036_ (
    .A(\datapath.registers.rega_data [7]),
    .B(_388__bF$buf2),
    .Y(_410_)
);

NAND2X1 _10037_ (
    .A(\datapath.idpc [7]),
    .B(_386__bF$buf1),
    .Y(_411_)
);

NAND2X1 _10038_ (
    .A(\datapath.csr.csr_data [7]),
    .B(_387__bF$buf1),
    .Y(_412_)
);

NAND3X1 _10039_ (
    .A(_411_),
    .B(_412_),
    .C(_410_),
    .Y(\datapath.muxaval [7])
);

NAND2X1 _10040_ (
    .A(\datapath.registers.rega_data [8]),
    .B(_388__bF$buf1),
    .Y(_413_)
);

NAND2X1 _10041_ (
    .A(\datapath.idpc [8]),
    .B(_386__bF$buf0),
    .Y(_414_)
);

NAND2X1 _10042_ (
    .A(\datapath.csr.csr_data [8]),
    .B(_387__bF$buf0),
    .Y(_415_)
);

NAND3X1 _10043_ (
    .A(_414_),
    .B(_415_),
    .C(_413_),
    .Y(\datapath.muxaval [8])
);

NAND2X1 _10044_ (
    .A(\datapath.registers.rega_data [9]),
    .B(_388__bF$buf0),
    .Y(_416_)
);

NAND2X1 _10045_ (
    .A(\datapath.idpc [9]),
    .B(_386__bF$buf4),
    .Y(_417_)
);

NAND2X1 _10046_ (
    .A(\datapath.csr.csr_data [9]),
    .B(_387__bF$buf4),
    .Y(_418_)
);

NAND3X1 _10047_ (
    .A(_417_),
    .B(_418_),
    .C(_416_),
    .Y(\datapath.muxaval [9])
);

NAND2X1 _10048_ (
    .A(\datapath.registers.rega_data [10]),
    .B(_388__bF$buf4),
    .Y(_419_)
);

NAND2X1 _10049_ (
    .A(\datapath.idpc [10]),
    .B(_386__bF$buf3),
    .Y(_420_)
);

NAND2X1 _10050_ (
    .A(\datapath.csr.csr_data [10]),
    .B(_387__bF$buf3),
    .Y(_421_)
);

NAND3X1 _10051_ (
    .A(_420_),
    .B(_421_),
    .C(_419_),
    .Y(\datapath.muxaval [10])
);

NAND2X1 _10052_ (
    .A(\datapath.registers.rega_data [11]),
    .B(_388__bF$buf3),
    .Y(_422_)
);

NAND2X1 _10053_ (
    .A(\datapath.idpc [11]),
    .B(_386__bF$buf2),
    .Y(_423_)
);

NAND2X1 _10054_ (
    .A(\datapath.csr.csr_data [11]),
    .B(_387__bF$buf2),
    .Y(_424_)
);

NAND3X1 _10055_ (
    .A(_423_),
    .B(_424_),
    .C(_422_),
    .Y(\datapath.muxaval [11])
);

NAND2X1 _10056_ (
    .A(\datapath.registers.rega_data [12]),
    .B(_388__bF$buf2),
    .Y(_425_)
);

NAND2X1 _10057_ (
    .A(\datapath.idpc [12]),
    .B(_386__bF$buf1),
    .Y(_426_)
);

NAND2X1 _10058_ (
    .A(\datapath.csr.csr_data [12]),
    .B(_387__bF$buf1),
    .Y(_427_)
);

NAND3X1 _10059_ (
    .A(_426_),
    .B(_427_),
    .C(_425_),
    .Y(\datapath.muxaval [12])
);

NAND2X1 _10060_ (
    .A(\datapath.registers.rega_data [13]),
    .B(_388__bF$buf1),
    .Y(_428_)
);

NAND2X1 _10061_ (
    .A(\datapath.idpc [13]),
    .B(_386__bF$buf0),
    .Y(_429_)
);

NAND2X1 _10062_ (
    .A(\datapath.csr.csr_data [13]),
    .B(_387__bF$buf0),
    .Y(_430_)
);

NAND3X1 _10063_ (
    .A(_429_),
    .B(_430_),
    .C(_428_),
    .Y(\datapath.muxaval [13])
);

NAND2X1 _10064_ (
    .A(\datapath.registers.rega_data [14]),
    .B(_388__bF$buf0),
    .Y(_431_)
);

NAND2X1 _10065_ (
    .A(\datapath.idpc [14]),
    .B(_386__bF$buf4),
    .Y(_432_)
);

NAND2X1 _10066_ (
    .A(\datapath.csr.csr_data [14]),
    .B(_387__bF$buf4),
    .Y(_433_)
);

NAND3X1 _10067_ (
    .A(_432_),
    .B(_433_),
    .C(_431_),
    .Y(\datapath.muxaval [14])
);

NAND2X1 _10068_ (
    .A(\datapath.registers.rega_data [15]),
    .B(_388__bF$buf4),
    .Y(_434_)
);

NAND2X1 _10069_ (
    .A(\datapath.idpc [15]),
    .B(_386__bF$buf3),
    .Y(_435_)
);

NAND2X1 _10070_ (
    .A(\datapath.csr.csr_data [15]),
    .B(_387__bF$buf3),
    .Y(_436_)
);

NAND3X1 _10071_ (
    .A(_435_),
    .B(_436_),
    .C(_434_),
    .Y(\datapath.muxaval [15])
);

NAND2X1 _10072_ (
    .A(\datapath.registers.rega_data [16]),
    .B(_388__bF$buf3),
    .Y(_437_)
);

NAND2X1 _10073_ (
    .A(\datapath.idpc [16]),
    .B(_386__bF$buf2),
    .Y(_438_)
);

NAND2X1 _10074_ (
    .A(\datapath.csr.csr_data [16]),
    .B(_387__bF$buf2),
    .Y(_439_)
);

NAND3X1 _10075_ (
    .A(_438_),
    .B(_439_),
    .C(_437_),
    .Y(\datapath.muxaval [16])
);

NAND2X1 _10076_ (
    .A(\datapath.registers.rega_data [17]),
    .B(_388__bF$buf2),
    .Y(_440_)
);

NAND2X1 _10077_ (
    .A(\datapath.idpc [17]),
    .B(_386__bF$buf1),
    .Y(_441_)
);

NAND2X1 _10078_ (
    .A(\datapath.csr.csr_data [17]),
    .B(_387__bF$buf1),
    .Y(_442_)
);

NAND3X1 _10079_ (
    .A(_441_),
    .B(_442_),
    .C(_440_),
    .Y(\datapath.muxaval [17])
);

NAND2X1 _10080_ (
    .A(\datapath.registers.rega_data [18]),
    .B(_388__bF$buf1),
    .Y(_443_)
);

NAND2X1 _10081_ (
    .A(\datapath.idpc [18]),
    .B(_386__bF$buf0),
    .Y(_444_)
);

NAND2X1 _10082_ (
    .A(\datapath.csr.csr_data [18]),
    .B(_387__bF$buf0),
    .Y(_445_)
);

NAND3X1 _10083_ (
    .A(_444_),
    .B(_445_),
    .C(_443_),
    .Y(\datapath.muxaval [18])
);

NAND2X1 _10084_ (
    .A(\datapath.registers.rega_data [19]),
    .B(_388__bF$buf0),
    .Y(_446_)
);

NAND2X1 _10085_ (
    .A(\datapath.idpc [19]),
    .B(_386__bF$buf4),
    .Y(_447_)
);

NAND2X1 _10086_ (
    .A(\datapath.csr.csr_data [19]),
    .B(_387__bF$buf4),
    .Y(_448_)
);

NAND3X1 _10087_ (
    .A(_447_),
    .B(_448_),
    .C(_446_),
    .Y(\datapath.muxaval [19])
);

NAND2X1 _10088_ (
    .A(\datapath.registers.rega_data [20]),
    .B(_388__bF$buf4),
    .Y(_449_)
);

NAND2X1 _10089_ (
    .A(\datapath.idpc [20]),
    .B(_386__bF$buf3),
    .Y(_450_)
);

NAND2X1 _10090_ (
    .A(\datapath.csr.csr_data [20]),
    .B(_387__bF$buf3),
    .Y(_451_)
);

NAND3X1 _10091_ (
    .A(_450_),
    .B(_451_),
    .C(_449_),
    .Y(\datapath.muxaval [20])
);

NAND2X1 _10092_ (
    .A(\datapath.registers.rega_data [21]),
    .B(_388__bF$buf3),
    .Y(_452_)
);

NAND2X1 _10093_ (
    .A(\datapath.idpc [21]),
    .B(_386__bF$buf2),
    .Y(_453_)
);

NAND2X1 _10094_ (
    .A(\datapath.csr.csr_data [21]),
    .B(_387__bF$buf2),
    .Y(_454_)
);

NAND3X1 _10095_ (
    .A(_453_),
    .B(_454_),
    .C(_452_),
    .Y(\datapath.muxaval [21])
);

NAND2X1 _10096_ (
    .A(\datapath.registers.rega_data [22]),
    .B(_388__bF$buf2),
    .Y(_455_)
);

NAND2X1 _10097_ (
    .A(\datapath.idpc [22]),
    .B(_386__bF$buf1),
    .Y(_456_)
);

NAND2X1 _10098_ (
    .A(\datapath.csr.csr_data [22]),
    .B(_387__bF$buf1),
    .Y(_457_)
);

NAND3X1 _10099_ (
    .A(_456_),
    .B(_457_),
    .C(_455_),
    .Y(\datapath.muxaval [22])
);

NAND2X1 _10100_ (
    .A(\datapath.registers.rega_data [23]),
    .B(_388__bF$buf1),
    .Y(_458_)
);

NAND2X1 _10101_ (
    .A(\datapath.idpc [23]),
    .B(_386__bF$buf0),
    .Y(_459_)
);

NAND2X1 _10102_ (
    .A(\datapath.csr.csr_data [23]),
    .B(_387__bF$buf0),
    .Y(_460_)
);

NAND3X1 _10103_ (
    .A(_459_),
    .B(_460_),
    .C(_458_),
    .Y(\datapath.muxaval [23])
);

NAND2X1 _10104_ (
    .A(\datapath.registers.rega_data [24]),
    .B(_388__bF$buf0),
    .Y(_461_)
);

NAND2X1 _10105_ (
    .A(\datapath.idpc [24]),
    .B(_386__bF$buf4),
    .Y(_462_)
);

NAND2X1 _10106_ (
    .A(\datapath.csr.csr_data [24]),
    .B(_387__bF$buf4),
    .Y(_463_)
);

NAND3X1 _10107_ (
    .A(_462_),
    .B(_463_),
    .C(_461_),
    .Y(\datapath.muxaval [24])
);

NAND2X1 _10108_ (
    .A(\datapath.registers.rega_data [25]),
    .B(_388__bF$buf4),
    .Y(_464_)
);

NAND2X1 _10109_ (
    .A(\datapath.idpc [25]),
    .B(_386__bF$buf3),
    .Y(_465_)
);

NAND2X1 _10110_ (
    .A(\datapath.csr.csr_data [25]),
    .B(_387__bF$buf3),
    .Y(_466_)
);

NAND3X1 _10111_ (
    .A(_465_),
    .B(_466_),
    .C(_464_),
    .Y(\datapath.muxaval [25])
);

NAND2X1 _10112_ (
    .A(\datapath.registers.rega_data [26]),
    .B(_388__bF$buf3),
    .Y(_467_)
);

NAND2X1 _10113_ (
    .A(\datapath.idpc [26]),
    .B(_386__bF$buf2),
    .Y(_468_)
);

NAND2X1 _10114_ (
    .A(\datapath.csr.csr_data [26]),
    .B(_387__bF$buf2),
    .Y(_469_)
);

NAND3X1 _10115_ (
    .A(_468_),
    .B(_469_),
    .C(_467_),
    .Y(\datapath.muxaval [26])
);

NAND2X1 _10116_ (
    .A(\datapath.registers.rega_data [27]),
    .B(_388__bF$buf2),
    .Y(_470_)
);

NAND2X1 _10117_ (
    .A(\datapath.idpc [27]),
    .B(_386__bF$buf1),
    .Y(_471_)
);

NAND2X1 _10118_ (
    .A(\datapath.csr.csr_data [27]),
    .B(_387__bF$buf1),
    .Y(_472_)
);

NAND3X1 _10119_ (
    .A(_471_),
    .B(_472_),
    .C(_470_),
    .Y(\datapath.muxaval [27])
);

NAND2X1 _10120_ (
    .A(\datapath.registers.rega_data [28]),
    .B(_388__bF$buf1),
    .Y(_473_)
);

NAND2X1 _10121_ (
    .A(\datapath.idpc [28]),
    .B(_386__bF$buf0),
    .Y(_474_)
);

NAND2X1 _10122_ (
    .A(\datapath.csr.csr_data [28]),
    .B(_387__bF$buf0),
    .Y(_475_)
);

NAND3X1 _10123_ (
    .A(_474_),
    .B(_475_),
    .C(_473_),
    .Y(\datapath.muxaval [28])
);

NAND2X1 _10124_ (
    .A(\datapath.registers.rega_data [29]),
    .B(_388__bF$buf0),
    .Y(_476_)
);

NAND2X1 _10125_ (
    .A(\datapath.idpc [29]),
    .B(_386__bF$buf4),
    .Y(_477_)
);

NAND2X1 _10126_ (
    .A(\datapath.csr.csr_data [29]),
    .B(_387__bF$buf4),
    .Y(_478_)
);

NAND3X1 _10127_ (
    .A(_477_),
    .B(_478_),
    .C(_476_),
    .Y(\datapath.muxaval [29])
);

NAND2X1 _10128_ (
    .A(\datapath.registers.rega_data [30]),
    .B(_388__bF$buf4),
    .Y(_479_)
);

NAND2X1 _10129_ (
    .A(\datapath.idpc [30]),
    .B(_386__bF$buf3),
    .Y(_480_)
);

NAND2X1 _10130_ (
    .A(\datapath.csr.csr_data [30]),
    .B(_387__bF$buf3),
    .Y(_481_)
);

NAND3X1 _10131_ (
    .A(_480_),
    .B(_481_),
    .C(_479_),
    .Y(\datapath.muxaval [30])
);

NAND2X1 _10132_ (
    .A(\datapath.registers.rega_data [31]),
    .B(_388__bF$buf3),
    .Y(_482_)
);

NAND2X1 _10133_ (
    .A(\datapath.idpc [31]),
    .B(_386__bF$buf2),
    .Y(_483_)
);

NAND2X1 _10134_ (
    .A(\datapath.csr.csr_data [31]),
    .B(_387__bF$buf2),
    .Y(_484_)
);

NAND3X1 _10135_ (
    .A(_483_),
    .B(_484_),
    .C(_482_),
    .Y(\datapath.muxaval [31])
);

INVX1 _10136_ (
    .A(\controlunit.csrfile_wen ),
    .Y(_485_)
);

INVX1 _10137_ (
    .A(\datapath.meminstr [17]),
    .Y(_486_)
);

INVX1 _10138_ (
    .A(\datapath.meminstr [16]),
    .Y(_487_)
);

NOR2X1 _10139_ (
    .A(\datapath.meminstr [18]),
    .B(\datapath.meminstr [19]),
    .Y(_488_)
);

NAND3X1 _10140_ (
    .A(_486_),
    .B(_487_),
    .C(_488_),
    .Y(_489_)
);

NOR2X1 _10141_ (
    .A(\datapath.meminstr [15]),
    .B(_489_),
    .Y(_490_)
);

AOI21X1 _10142_ (
    .A(_490_),
    .B(\datapath.meminstr [13]),
    .C(_485_),
    .Y(\datapath.allowcsrwrite )
);

NAND2X1 _10143_ (
    .A(_179_),
    .B(\datapath.csr.csr_mcause [2]),
    .Y(\controlunit.csrfile_trap_wen )
);

INVX1 _10144_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf7 ),
    .Y(_491_)
);

NOR2X1 _10145_ (
    .A(\datapath.regpcsel [0]),
    .B(\datapath.regmret ),
    .Y(_492_)
);

NAND3X1 _10146_ (
    .A(_161_),
    .B(_492_),
    .C(_491_),
    .Y(\datapath._34_ )
);

NOR2X1 _10147_ (
    .A(\datapath.regmret ),
    .B(\datapath.regpcsel [1]),
    .Y(_493_)
);

NAND2X1 _10148_ (
    .A(_493_),
    .B(_491_),
    .Y(\datapath._36_ )
);

NAND2X1 _10149_ (
    .A(\datapath.regimmalu [0]),
    .B(\datapath.alupc [0]),
    .Y(_494_)
);

NAND2X1 _10150_ (
    .A(\datapath.regimmalu [1]),
    .B(\datapath.alupc [1]),
    .Y(_495_)
);

INVX1 _10151_ (
    .A(_495_),
    .Y(_496_)
);

NOR2X1 _10152_ (
    .A(\datapath.regimmalu [1]),
    .B(\datapath.alupc [1]),
    .Y(_497_)
);

NOR2X1 _10153_ (
    .A(_497_),
    .B(_496_),
    .Y(_498_)
);

XNOR2X1 _10154_ (
    .A(_498_),
    .B(_494_),
    .Y(\datapath.jumptarget [1])
);

OAI21X1 _10155_ (
    .A(_494_),
    .B(_497_),
    .C(_495_),
    .Y(_499_)
);

AND2X2 _10156_ (
    .A(\datapath.regimmalu [2]),
    .B(\datapath.alupc [2]),
    .Y(_500_)
);

NOR2X1 _10157_ (
    .A(\datapath.regimmalu [2]),
    .B(\datapath.alupc [2]),
    .Y(_501_)
);

NOR2X1 _10158_ (
    .A(_501_),
    .B(_500_),
    .Y(_502_)
);

XOR2X1 _10159_ (
    .A(_499_),
    .B(_502_),
    .Y(\datapath.jumptarget [2])
);

AOI21X1 _10160_ (
    .A(_499_),
    .B(_502_),
    .C(_500_),
    .Y(_503_)
);

AND2X2 _10161_ (
    .A(\datapath.regimmalu [3]),
    .B(\datapath.alupc [3]),
    .Y(_504_)
);

NOR2X1 _10162_ (
    .A(\datapath.regimmalu [3]),
    .B(\datapath.alupc [3]),
    .Y(_505_)
);

NOR2X1 _10163_ (
    .A(_505_),
    .B(_504_),
    .Y(_506_)
);

XNOR2X1 _10164_ (
    .A(_503_),
    .B(_506_),
    .Y(\datapath.jumptarget [3])
);

NAND3X1 _10165_ (
    .A(_502_),
    .B(_499_),
    .C(_506_),
    .Y(_507_)
);

INVX1 _10166_ (
    .A(_505_),
    .Y(_508_)
);

AOI21X1 _10167_ (
    .A(_508_),
    .B(_500_),
    .C(_504_),
    .Y(_509_)
);

NAND2X1 _10168_ (
    .A(_509_),
    .B(_507_),
    .Y(_510_)
);

NAND2X1 _10169_ (
    .A(\datapath.regimmalu [4]),
    .B(\datapath.alupc [4]),
    .Y(_511_)
);

OR2X2 _10170_ (
    .A(\datapath.regimmalu [4]),
    .B(\datapath.alupc [4]),
    .Y(_512_)
);

NAND2X1 _10171_ (
    .A(_511_),
    .B(_512_),
    .Y(_513_)
);

XNOR2X1 _10172_ (
    .A(_510_),
    .B(_513_),
    .Y(\datapath.jumptarget [4])
);

INVX1 _10173_ (
    .A(_510_),
    .Y(_514_)
);

NOR2X1 _10174_ (
    .A(\datapath.regimmalu [4]),
    .B(\datapath.alupc [4]),
    .Y(_515_)
);

OAI21X1 _10175_ (
    .A(_515_),
    .B(_514_),
    .C(_511_),
    .Y(_516_)
);

XOR2X1 _10176_ (
    .A(\datapath.regimmalu [5]),
    .B(\datapath.alupc [5]),
    .Y(_517_)
);

XOR2X1 _10177_ (
    .A(_516_),
    .B(_517_),
    .Y(\datapath.jumptarget [5])
);

INVX1 _10178_ (
    .A(\datapath.regimmalu [5]),
    .Y(_518_)
);

INVX1 _10179_ (
    .A(\datapath.alupc [5]),
    .Y(_519_)
);

OAI21X1 _10180_ (
    .A(_518_),
    .B(_519_),
    .C(_511_),
    .Y(_520_)
);

OAI21X1 _10181_ (
    .A(\datapath.regimmalu [5]),
    .B(\datapath.alupc [5]),
    .C(_520_),
    .Y(_521_)
);

AND2X2 _10182_ (
    .A(\datapath.regimmalu [4]),
    .B(\datapath.alupc [4]),
    .Y(_522_)
);

NOR2X1 _10183_ (
    .A(_515_),
    .B(_522_),
    .Y(_523_)
);

NAND2X1 _10184_ (
    .A(_523_),
    .B(_517_),
    .Y(_524_)
);

OAI21X1 _10185_ (
    .A(_524_),
    .B(_514_),
    .C(_521_),
    .Y(_525_)
);

AND2X2 _10186_ (
    .A(\datapath.regimmalu [6]),
    .B(\datapath.alupc [6]),
    .Y(_526_)
);

NOR2X1 _10187_ (
    .A(\datapath.regimmalu [6]),
    .B(\datapath.alupc [6]),
    .Y(_527_)
);

NOR2X1 _10188_ (
    .A(_527_),
    .B(_526_),
    .Y(_528_)
);

XOR2X1 _10189_ (
    .A(_525_),
    .B(_528_),
    .Y(\datapath.jumptarget [6])
);

AOI21X1 _10190_ (
    .A(_525_),
    .B(_528_),
    .C(_526_),
    .Y(_529_)
);

AND2X2 _10191_ (
    .A(\datapath.regimmalu [7]),
    .B(\datapath.alupc [7]),
    .Y(_530_)
);

NOR2X1 _10192_ (
    .A(\datapath.regimmalu [7]),
    .B(\datapath.alupc [7]),
    .Y(_531_)
);

NOR2X1 _10193_ (
    .A(_531_),
    .B(_530_),
    .Y(_532_)
);

XNOR2X1 _10194_ (
    .A(_529_),
    .B(_532_),
    .Y(\datapath.jumptarget [7])
);

NAND2X1 _10195_ (
    .A(_528_),
    .B(_532_),
    .Y(_533_)
);

NOR2X1 _10196_ (
    .A(_524_),
    .B(_533_),
    .Y(_534_)
);

OR2X2 _10197_ (
    .A(\datapath.regimmalu [7]),
    .B(\datapath.alupc [7]),
    .Y(_535_)
);

AOI21X1 _10198_ (
    .A(_535_),
    .B(_526_),
    .C(_530_),
    .Y(_536_)
);

OAI21X1 _10199_ (
    .A(_521_),
    .B(_533_),
    .C(_536_),
    .Y(_537_)
);

AOI21X1 _10200_ (
    .A(_534_),
    .B(_510_),
    .C(_537_),
    .Y(_538_)
);

NAND2X1 _10201_ (
    .A(\datapath.regimmalu [8]),
    .B(\datapath.alupc [8]),
    .Y(_539_)
);

INVX1 _10202_ (
    .A(\datapath.regimmalu [8]),
    .Y(_540_)
);

INVX1 _10203_ (
    .A(\datapath.alupc [8]),
    .Y(_541_)
);

NAND2X1 _10204_ (
    .A(_540_),
    .B(_541_),
    .Y(_542_)
);

NAND2X1 _10205_ (
    .A(_539_),
    .B(_542_),
    .Y(_543_)
);

XOR2X1 _10206_ (
    .A(_538_),
    .B(_543_),
    .Y(\datapath.jumptarget [8])
);

OAI21X1 _10207_ (
    .A(_543_),
    .B(_538_),
    .C(_539_),
    .Y(_544_)
);

INVX1 _10208_ (
    .A(\datapath.regimmalu [9]),
    .Y(_545_)
);

NAND2X1 _10209_ (
    .A(\datapath.alupc [9]),
    .B(_545_),
    .Y(_546_)
);

INVX1 _10210_ (
    .A(\datapath.alupc [9]),
    .Y(_547_)
);

NAND2X1 _10211_ (
    .A(\datapath.regimmalu [9]),
    .B(_547_),
    .Y(_548_)
);

AND2X2 _10212_ (
    .A(_546_),
    .B(_548_),
    .Y(_549_)
);

XNOR2X1 _10213_ (
    .A(_544_),
    .B(_549_),
    .Y(\datapath.jumptarget [9])
);

OAI21X1 _10214_ (
    .A(_545_),
    .B(_547_),
    .C(_539_),
    .Y(_550_)
);

OAI21X1 _10215_ (
    .A(\datapath.regimmalu [9]),
    .B(\datapath.alupc [9]),
    .C(_550_),
    .Y(_551_)
);

NAND2X1 _10216_ (
    .A(\datapath.alupc [5]),
    .B(_518_),
    .Y(_552_)
);

NAND2X1 _10217_ (
    .A(\datapath.regimmalu [5]),
    .B(_519_),
    .Y(_553_)
);

AOI21X1 _10218_ (
    .A(_552_),
    .B(_553_),
    .C(_513_),
    .Y(_554_)
);

INVX1 _10219_ (
    .A(\datapath.alupc [6]),
    .Y(_555_)
);

OR2X2 _10220_ (
    .A(_555_),
    .B(\datapath.regimmalu [6]),
    .Y(_556_)
);

NAND2X1 _10221_ (
    .A(\datapath.regimmalu [6]),
    .B(_555_),
    .Y(_557_)
);

NAND2X1 _10222_ (
    .A(\datapath.regimmalu [7]),
    .B(\datapath.alupc [7]),
    .Y(_558_)
);

NAND2X1 _10223_ (
    .A(_558_),
    .B(_535_),
    .Y(_559_)
);

AOI21X1 _10224_ (
    .A(_556_),
    .B(_557_),
    .C(_559_),
    .Y(_560_)
);

NAND2X1 _10225_ (
    .A(_560_),
    .B(_554_),
    .Y(_561_)
);

AOI21X1 _10226_ (
    .A(_507_),
    .B(_509_),
    .C(_561_),
    .Y(_562_)
);

NAND2X1 _10227_ (
    .A(\datapath.alupc [8]),
    .B(_540_),
    .Y(_563_)
);

NAND2X1 _10228_ (
    .A(\datapath.regimmalu [8]),
    .B(_541_),
    .Y(_564_)
);

AOI22X1 _10229_ (
    .A(_563_),
    .B(_564_),
    .C(_546_),
    .D(_548_),
    .Y(_565_)
);

OAI21X1 _10230_ (
    .A(_537_),
    .B(_562_),
    .C(_565_),
    .Y(_566_)
);

NAND2X1 _10231_ (
    .A(_551_),
    .B(_566_),
    .Y(_567_)
);

AND2X2 _10232_ (
    .A(\datapath.regimmalu [10]),
    .B(\datapath.alupc [10]),
    .Y(_568_)
);

NOR2X1 _10233_ (
    .A(\datapath.regimmalu [10]),
    .B(\datapath.alupc [10]),
    .Y(_569_)
);

NOR2X1 _10234_ (
    .A(_569_),
    .B(_568_),
    .Y(_570_)
);

XOR2X1 _10235_ (
    .A(_567_),
    .B(_570_),
    .Y(\datapath.jumptarget [10])
);

AOI21X1 _10236_ (
    .A(_567_),
    .B(_570_),
    .C(_568_),
    .Y(_571_)
);

AND2X2 _10237_ (
    .A(\datapath.regimmalu [11]),
    .B(\datapath.alupc [11]),
    .Y(_572_)
);

NOR2X1 _10238_ (
    .A(\datapath.regimmalu [11]),
    .B(\datapath.alupc [11]),
    .Y(_573_)
);

NOR2X1 _10239_ (
    .A(_573_),
    .B(_572_),
    .Y(_574_)
);

XNOR2X1 _10240_ (
    .A(_571_),
    .B(_574_),
    .Y(\datapath.jumptarget [11])
);

NAND2X1 _10241_ (
    .A(_570_),
    .B(_574_),
    .Y(_575_)
);

AOI21X1 _10242_ (
    .A(_574_),
    .B(_568_),
    .C(_572_),
    .Y(_576_)
);

OAI21X1 _10243_ (
    .A(_551_),
    .B(_575_),
    .C(_576_),
    .Y(_577_)
);

NAND3X1 _10244_ (
    .A(_570_),
    .B(_574_),
    .C(_565_),
    .Y(_578_)
);

NOR2X1 _10245_ (
    .A(_578_),
    .B(_538_),
    .Y(_579_)
);

AND2X2 _10246_ (
    .A(\datapath.regimmalu [12]),
    .B(\datapath.alupc [12]),
    .Y(_580_)
);

NOR2X1 _10247_ (
    .A(\datapath.regimmalu [12]),
    .B(\datapath.alupc [12]),
    .Y(_581_)
);

NOR2X1 _10248_ (
    .A(_581_),
    .B(_580_),
    .Y(_582_)
);

OAI21X1 _10249_ (
    .A(_577_),
    .B(_579_),
    .C(_582_),
    .Y(_583_)
);

NOR2X1 _10250_ (
    .A(_577_),
    .B(_579_),
    .Y(_584_)
);

OAI21X1 _10251_ (
    .A(_580_),
    .B(_581_),
    .C(_584_),
    .Y(_585_)
);

AND2X2 _10252_ (
    .A(_585_),
    .B(_583_),
    .Y(\datapath.jumptarget [12])
);

NAND2X1 _10253_ (
    .A(\datapath.regimmalu [12]),
    .B(\datapath.alupc [12]),
    .Y(_586_)
);

OAI21X1 _10254_ (
    .A(_581_),
    .B(_584_),
    .C(_586_),
    .Y(_587_)
);

AND2X2 _10255_ (
    .A(\datapath.regimmalu [13]),
    .B(\datapath.alupc [13]),
    .Y(_588_)
);

NOR2X1 _10256_ (
    .A(\datapath.regimmalu [13]),
    .B(\datapath.alupc [13]),
    .Y(_589_)
);

NOR2X1 _10257_ (
    .A(_589_),
    .B(_588_),
    .Y(_590_)
);

XOR2X1 _10258_ (
    .A(_587_),
    .B(_590_),
    .Y(\datapath.jumptarget [13])
);

NAND2X1 _10259_ (
    .A(\datapath.regimmalu [13]),
    .B(\datapath.alupc [13]),
    .Y(_591_)
);

OAI21X1 _10260_ (
    .A(_586_),
    .B(_589_),
    .C(_591_),
    .Y(_592_)
);

NAND2X1 _10261_ (
    .A(_582_),
    .B(_590_),
    .Y(_593_)
);

NOR2X1 _10262_ (
    .A(_593_),
    .B(_584_),
    .Y(_594_)
);

NOR2X1 _10263_ (
    .A(_592_),
    .B(_594_),
    .Y(_595_)
);

AND2X2 _10264_ (
    .A(\datapath.regimmalu [14]),
    .B(\datapath.alupc [14]),
    .Y(_596_)
);

NOR2X1 _10265_ (
    .A(\datapath.regimmalu [14]),
    .B(\datapath.alupc [14]),
    .Y(_597_)
);

NOR2X1 _10266_ (
    .A(_597_),
    .B(_596_),
    .Y(_598_)
);

XNOR2X1 _10267_ (
    .A(_595_),
    .B(_598_),
    .Y(\datapath.jumptarget [14])
);

INVX1 _10268_ (
    .A(_596_),
    .Y(_599_)
);

OAI21X1 _10269_ (
    .A(_597_),
    .B(_595_),
    .C(_599_),
    .Y(_600_)
);

AND2X2 _10270_ (
    .A(\datapath.regimmalu [15]),
    .B(\datapath.alupc [15]),
    .Y(_601_)
);

NOR2X1 _10271_ (
    .A(\datapath.regimmalu [15]),
    .B(\datapath.alupc [15]),
    .Y(_602_)
);

NOR2X1 _10272_ (
    .A(_602_),
    .B(_601_),
    .Y(_603_)
);

XOR2X1 _10273_ (
    .A(_600_),
    .B(_603_),
    .Y(\datapath.jumptarget [15])
);

INVX1 _10274_ (
    .A(_575_),
    .Y(_604_)
);

NAND2X1 _10275_ (
    .A(_598_),
    .B(_603_),
    .Y(_605_)
);

NOR2X1 _10276_ (
    .A(_593_),
    .B(_605_),
    .Y(_606_)
);

NAND3X1 _10277_ (
    .A(_565_),
    .B(_604_),
    .C(_606_),
    .Y(_607_)
);

INVX1 _10278_ (
    .A(_592_),
    .Y(_608_)
);

AOI21X1 _10279_ (
    .A(_603_),
    .B(_596_),
    .C(_601_),
    .Y(_609_)
);

OAI21X1 _10280_ (
    .A(_608_),
    .B(_605_),
    .C(_609_),
    .Y(_610_)
);

AOI21X1 _10281_ (
    .A(_577_),
    .B(_606_),
    .C(_610_),
    .Y(_611_)
);

OAI21X1 _10282_ (
    .A(_607_),
    .B(_538_),
    .C(_611_),
    .Y(_612_)
);

AND2X2 _10283_ (
    .A(\datapath.regimmalu [16]),
    .B(\datapath.alupc [16]),
    .Y(_613_)
);

NOR2X1 _10284_ (
    .A(\datapath.regimmalu [16]),
    .B(\datapath.alupc [16]),
    .Y(_614_)
);

NOR2X1 _10285_ (
    .A(_614_),
    .B(_613_),
    .Y(_615_)
);

XOR2X1 _10286_ (
    .A(_612_),
    .B(_615_),
    .Y(\datapath.jumptarget [16])
);

AOI21X1 _10287_ (
    .A(_612_),
    .B(_615_),
    .C(_613_),
    .Y(_616_)
);

INVX1 _10288_ (
    .A(\datapath.regimmalu [17]),
    .Y(_617_)
);

INVX1 _10289_ (
    .A(\datapath.alupc [17]),
    .Y(_618_)
);

NOR2X1 _10290_ (
    .A(_617_),
    .B(_618_),
    .Y(_619_)
);

NOR2X1 _10291_ (
    .A(\datapath.regimmalu [17]),
    .B(\datapath.alupc [17]),
    .Y(_620_)
);

NOR2X1 _10292_ (
    .A(_620_),
    .B(_619_),
    .Y(_621_)
);

XNOR2X1 _10293_ (
    .A(_616_),
    .B(_621_),
    .Y(\datapath.jumptarget [17])
);

NOR3X1 _10294_ (
    .A(_593_),
    .B(_605_),
    .C(_578_),
    .Y(_622_)
);

OAI21X1 _10295_ (
    .A(_537_),
    .B(_562_),
    .C(_622_),
    .Y(_623_)
);

AND2X2 _10296_ (
    .A(_623_),
    .B(_611_),
    .Y(_624_)
);

INVX1 _10297_ (
    .A(_620_),
    .Y(_625_)
);

AOI21X1 _10298_ (
    .A(_625_),
    .B(_613_),
    .C(_619_),
    .Y(_626_)
);

NAND2X1 _10299_ (
    .A(_615_),
    .B(_621_),
    .Y(_627_)
);

OAI21X1 _10300_ (
    .A(_627_),
    .B(_624_),
    .C(_626_),
    .Y(_628_)
);

AND2X2 _10301_ (
    .A(\datapath.regimmalu [18]),
    .B(\datapath.alupc [18]),
    .Y(_629_)
);

NOR2X1 _10302_ (
    .A(\datapath.regimmalu [18]),
    .B(\datapath.alupc [18]),
    .Y(_630_)
);

NOR2X1 _10303_ (
    .A(_630_),
    .B(_629_),
    .Y(_631_)
);

XOR2X1 _10304_ (
    .A(_628_),
    .B(_631_),
    .Y(\datapath.jumptarget [18])
);

AOI21X1 _10305_ (
    .A(_628_),
    .B(_631_),
    .C(_629_),
    .Y(_632_)
);

AND2X2 _10306_ (
    .A(\datapath.regimmalu [19]),
    .B(\datapath.alupc [19]),
    .Y(_633_)
);

NOR2X1 _10307_ (
    .A(\datapath.regimmalu [19]),
    .B(\datapath.alupc [19]),
    .Y(_634_)
);

NOR2X1 _10308_ (
    .A(_634_),
    .B(_633_),
    .Y(_635_)
);

XNOR2X1 _10309_ (
    .A(_632_),
    .B(_635_),
    .Y(\datapath.jumptarget [19])
);

NAND2X1 _10310_ (
    .A(_631_),
    .B(_635_),
    .Y(_636_)
);

AOI21X1 _10311_ (
    .A(_635_),
    .B(_629_),
    .C(_633_),
    .Y(_637_)
);

OAI21X1 _10312_ (
    .A(_626_),
    .B(_636_),
    .C(_637_),
    .Y(_638_)
);

OR2X2 _10313_ (
    .A(_627_),
    .B(_636_),
    .Y(_639_)
);

AOI21X1 _10314_ (
    .A(_623_),
    .B(_611_),
    .C(_639_),
    .Y(_640_)
);

NOR2X1 _10315_ (
    .A(_638_),
    .B(_640_),
    .Y(_641_)
);

NAND2X1 _10316_ (
    .A(\datapath.regimmalu [20]),
    .B(\datapath.alupc [20]),
    .Y(_642_)
);

OR2X2 _10317_ (
    .A(\datapath.regimmalu [20]),
    .B(\datapath.alupc [20]),
    .Y(_643_)
);

NAND2X1 _10318_ (
    .A(_642_),
    .B(_643_),
    .Y(_644_)
);

XOR2X1 _10319_ (
    .A(_641_),
    .B(_644_),
    .Y(\datapath.jumptarget [20])
);

OAI21X1 _10320_ (
    .A(_644_),
    .B(_641_),
    .C(_642_),
    .Y(_645_)
);

NAND2X1 _10321_ (
    .A(\datapath.regimmalu [21]),
    .B(\datapath.alupc [21]),
    .Y(_646_)
);

OR2X2 _10322_ (
    .A(\datapath.regimmalu [21]),
    .B(\datapath.alupc [21]),
    .Y(_647_)
);

NAND2X1 _10323_ (
    .A(_646_),
    .B(_647_),
    .Y(_648_)
);

XNOR2X1 _10324_ (
    .A(_645_),
    .B(_648_),
    .Y(\datapath.jumptarget [21])
);

OAI21X1 _10325_ (
    .A(_642_),
    .B(_648_),
    .C(_646_),
    .Y(_649_)
);

INVX1 _10326_ (
    .A(_649_),
    .Y(_650_)
);

NOR2X1 _10327_ (
    .A(_644_),
    .B(_648_),
    .Y(_651_)
);

OAI21X1 _10328_ (
    .A(_638_),
    .B(_640_),
    .C(_651_),
    .Y(_652_)
);

NAND2X1 _10329_ (
    .A(_650_),
    .B(_652_),
    .Y(_653_)
);

NAND2X1 _10330_ (
    .A(\datapath.regimmalu [22]),
    .B(\datapath.alupc [22]),
    .Y(_654_)
);

OR2X2 _10331_ (
    .A(\datapath.regimmalu [22]),
    .B(\datapath.alupc [22]),
    .Y(_655_)
);

NAND2X1 _10332_ (
    .A(_654_),
    .B(_655_),
    .Y(_656_)
);

XNOR2X1 _10333_ (
    .A(_653_),
    .B(_656_),
    .Y(\datapath.jumptarget [22])
);

INVX1 _10334_ (
    .A(_654_),
    .Y(_657_)
);

AOI21X1 _10335_ (
    .A(_653_),
    .B(_655_),
    .C(_657_),
    .Y(_658_)
);

AND2X2 _10336_ (
    .A(\datapath.regimmalu [23]),
    .B(\datapath.alupc [23]),
    .Y(_659_)
);

NOR2X1 _10337_ (
    .A(\datapath.regimmalu [23]),
    .B(\datapath.alupc [23]),
    .Y(_660_)
);

NOR2X1 _10338_ (
    .A(_660_),
    .B(_659_),
    .Y(_661_)
);

XNOR2X1 _10339_ (
    .A(_658_),
    .B(_661_),
    .Y(\datapath.jumptarget [23])
);

OR2X2 _10340_ (
    .A(_659_),
    .B(_660_),
    .Y(_662_)
);

NOR2X1 _10341_ (
    .A(_656_),
    .B(_662_),
    .Y(_663_)
);

NAND2X1 _10342_ (
    .A(_651_),
    .B(_663_),
    .Y(_664_)
);

NOR2X1 _10343_ (
    .A(_664_),
    .B(_639_),
    .Y(_665_)
);

NAND3X1 _10344_ (
    .A(_651_),
    .B(_663_),
    .C(_638_),
    .Y(_666_)
);

NAND2X1 _10345_ (
    .A(_649_),
    .B(_663_),
    .Y(_667_)
);

AOI21X1 _10346_ (
    .A(_661_),
    .B(_657_),
    .C(_659_),
    .Y(_668_)
);

NAND3X1 _10347_ (
    .A(_667_),
    .B(_668_),
    .C(_666_),
    .Y(_669_)
);

AOI21X1 _10348_ (
    .A(_612_),
    .B(_665_),
    .C(_669_),
    .Y(_670_)
);

INVX1 _10349_ (
    .A(\datapath.regimmalu [24]),
    .Y(_671_)
);

INVX1 _10350_ (
    .A(\datapath.alupc [24]),
    .Y(_672_)
);

NOR2X1 _10351_ (
    .A(_671_),
    .B(_672_),
    .Y(_673_)
);

NOR2X1 _10352_ (
    .A(\datapath.regimmalu [24]),
    .B(\datapath.alupc [24]),
    .Y(_674_)
);

NOR2X1 _10353_ (
    .A(_674_),
    .B(_673_),
    .Y(_675_)
);

XNOR2X1 _10354_ (
    .A(_670_),
    .B(_675_),
    .Y(\datapath.jumptarget [24])
);

INVX1 _10355_ (
    .A(_673_),
    .Y(_676_)
);

OAI21X1 _10356_ (
    .A(_674_),
    .B(_670_),
    .C(_676_),
    .Y(_677_)
);

AND2X2 _10357_ (
    .A(\datapath.regimmalu [25]),
    .B(\datapath.alupc [25]),
    .Y(_678_)
);

NOR2X1 _10358_ (
    .A(\datapath.regimmalu [25]),
    .B(\datapath.alupc [25]),
    .Y(_679_)
);

NOR2X1 _10359_ (
    .A(_679_),
    .B(_678_),
    .Y(_680_)
);

XOR2X1 _10360_ (
    .A(_677_),
    .B(_680_),
    .Y(\datapath.jumptarget [25])
);

AOI21X1 _10361_ (
    .A(_680_),
    .B(_673_),
    .C(_678_),
    .Y(_681_)
);

NAND2X1 _10362_ (
    .A(_680_),
    .B(_675_),
    .Y(_682_)
);

OAI21X1 _10363_ (
    .A(_682_),
    .B(_670_),
    .C(_681_),
    .Y(_683_)
);

AND2X2 _10364_ (
    .A(\datapath.regimmalu [26]),
    .B(\datapath.alupc [26]),
    .Y(_684_)
);

NOR2X1 _10365_ (
    .A(\datapath.regimmalu [26]),
    .B(\datapath.alupc [26]),
    .Y(_685_)
);

NOR2X1 _10366_ (
    .A(_685_),
    .B(_684_),
    .Y(_686_)
);

XOR2X1 _10367_ (
    .A(_683_),
    .B(_686_),
    .Y(\datapath.jumptarget [26])
);

AOI21X1 _10368_ (
    .A(_683_),
    .B(_686_),
    .C(_684_),
    .Y(_687_)
);

XOR2X1 _10369_ (
    .A(\datapath.regimmalu [27]),
    .B(\datapath.alupc [27]),
    .Y(_688_)
);

XNOR2X1 _10370_ (
    .A(_687_),
    .B(_688_),
    .Y(\datapath.jumptarget [27])
);

NAND2X1 _10371_ (
    .A(_686_),
    .B(_688_),
    .Y(_689_)
);

NOR2X1 _10372_ (
    .A(_689_),
    .B(_682_),
    .Y(_690_)
);

INVX1 _10373_ (
    .A(_690_),
    .Y(_691_)
);

NOR2X1 _10374_ (
    .A(_689_),
    .B(_681_),
    .Y(_692_)
);

INVX1 _10375_ (
    .A(\datapath.regimmalu [27]),
    .Y(_693_)
);

INVX1 _10376_ (
    .A(\datapath.alupc [27]),
    .Y(_694_)
);

OAI21X1 _10377_ (
    .A(\datapath.regimmalu [27]),
    .B(\datapath.alupc [27]),
    .C(_684_),
    .Y(_695_)
);

OAI21X1 _10378_ (
    .A(_693_),
    .B(_694_),
    .C(_695_),
    .Y(_696_)
);

NOR2X1 _10379_ (
    .A(_696_),
    .B(_692_),
    .Y(_697_)
);

OAI21X1 _10380_ (
    .A(_691_),
    .B(_670_),
    .C(_697_),
    .Y(_698_)
);

AND2X2 _10381_ (
    .A(\datapath.regimmalu [28]),
    .B(\datapath.alupc [28]),
    .Y(_699_)
);

NOR2X1 _10382_ (
    .A(\datapath.regimmalu [28]),
    .B(\datapath.alupc [28]),
    .Y(_700_)
);

NOR2X1 _10383_ (
    .A(_700_),
    .B(_699_),
    .Y(_701_)
);

INVX1 _10384_ (
    .A(_701_),
    .Y(_702_)
);

XNOR2X1 _10385_ (
    .A(_698_),
    .B(_702_),
    .Y(\datapath.jumptarget [28])
);

AOI21X1 _10386_ (
    .A(_698_),
    .B(_701_),
    .C(_699_),
    .Y(_703_)
);

INVX1 _10387_ (
    .A(\datapath.regimmalu [29]),
    .Y(_704_)
);

INVX1 _10388_ (
    .A(\datapath.alupc [29]),
    .Y(_705_)
);

NOR2X1 _10389_ (
    .A(_704_),
    .B(_705_),
    .Y(_706_)
);

NOR2X1 _10390_ (
    .A(\datapath.regimmalu [29]),
    .B(\datapath.alupc [29]),
    .Y(_707_)
);

NOR2X1 _10391_ (
    .A(_707_),
    .B(_706_),
    .Y(_708_)
);

XNOR2X1 _10392_ (
    .A(_703_),
    .B(_708_),
    .Y(\datapath.jumptarget [29])
);

INVX1 _10393_ (
    .A(_708_),
    .Y(_709_)
);

NOR2X1 _10394_ (
    .A(_702_),
    .B(_709_),
    .Y(_710_)
);

OAI21X1 _10395_ (
    .A(\datapath.regimmalu [29]),
    .B(\datapath.alupc [29]),
    .C(_699_),
    .Y(_711_)
);

OAI21X1 _10396_ (
    .A(_704_),
    .B(_705_),
    .C(_711_),
    .Y(_712_)
);

AOI21X1 _10397_ (
    .A(_698_),
    .B(_710_),
    .C(_712_),
    .Y(_713_)
);

NAND2X1 _10398_ (
    .A(\datapath.regimmalu [30]),
    .B(\datapath.alupc [30]),
    .Y(_714_)
);

OR2X2 _10399_ (
    .A(\datapath.regimmalu [30]),
    .B(\datapath.alupc [30]),
    .Y(_715_)
);

AND2X2 _10400_ (
    .A(_715_),
    .B(_714_),
    .Y(_716_)
);

XNOR2X1 _10401_ (
    .A(_713_),
    .B(_716_),
    .Y(\datapath.jumptarget [30])
);

OR2X2 _10402_ (
    .A(_639_),
    .B(_664_),
    .Y(_717_)
);

AOI21X1 _10403_ (
    .A(_623_),
    .B(_611_),
    .C(_717_),
    .Y(_718_)
);

OAI21X1 _10404_ (
    .A(_669_),
    .B(_718_),
    .C(_690_),
    .Y(_719_)
);

INVX1 _10405_ (
    .A(_710_),
    .Y(_720_)
);

AOI21X1 _10406_ (
    .A(_719_),
    .B(_697_),
    .C(_720_),
    .Y(_721_)
);

OAI21X1 _10407_ (
    .A(_712_),
    .B(_721_),
    .C(_716_),
    .Y(_722_)
);

XNOR2X1 _10408_ (
    .A(\datapath.regimmalu [31]),
    .B(\datapath.alupc [31]),
    .Y(_723_)
);

INVX1 _10409_ (
    .A(_723_),
    .Y(_724_)
);

NAND3X1 _10410_ (
    .A(_714_),
    .B(_724_),
    .C(_722_),
    .Y(_725_)
);

INVX1 _10411_ (
    .A(_716_),
    .Y(_726_)
);

OAI21X1 _10412_ (
    .A(_726_),
    .B(_713_),
    .C(_714_),
    .Y(_727_)
);

NAND2X1 _10413_ (
    .A(_723_),
    .B(_727_),
    .Y(_728_)
);

NAND2X1 _10414_ (
    .A(_725_),
    .B(_728_),
    .Y(\datapath.jumptarget [31])
);

XOR2X1 _10415_ (
    .A(\datapath.regimmalu [0]),
    .B(\datapath.alupc [0]),
    .Y(\datapath.jumptarget [0])
);

DFFPOSX1 _10416_ (
    .CLK(CLK_bF$buf151),
    .D(\datapath.csr.csr_wdata [0]),
    .Q(\datapath.regcsrwb [0])
);

DFFPOSX1 _10417_ (
    .CLK(CLK_bF$buf150),
    .D(\datapath.csr.csr_wdata [1]),
    .Q(\datapath.regcsrwb [1])
);

DFFPOSX1 _10418_ (
    .CLK(CLK_bF$buf149),
    .D(\datapath.csr.csr_wdata [2]),
    .Q(\datapath.regcsrwb [2])
);

DFFPOSX1 _10419_ (
    .CLK(CLK_bF$buf148),
    .D(\datapath.csr.csr_wdata [3]),
    .Q(\datapath.regcsrwb [3])
);

DFFPOSX1 _10420_ (
    .CLK(CLK_bF$buf147),
    .D(\datapath.csr.csr_wdata [4]),
    .Q(\datapath.regcsrwb [4])
);

DFFPOSX1 _10421_ (
    .CLK(CLK_bF$buf146),
    .D(\datapath.csr.csr_wdata [5]),
    .Q(\datapath.regcsrwb [5])
);

DFFPOSX1 _10422_ (
    .CLK(CLK_bF$buf145),
    .D(\datapath.csr.csr_wdata [6]),
    .Q(\datapath.regcsrwb [6])
);

DFFPOSX1 _10423_ (
    .CLK(CLK_bF$buf144),
    .D(\datapath.csr.csr_wdata [7]),
    .Q(\datapath.regcsrwb [7])
);

DFFPOSX1 _10424_ (
    .CLK(CLK_bF$buf143),
    .D(\datapath.csr.csr_wdata [8]),
    .Q(\datapath.regcsrwb [8])
);

DFFPOSX1 _10425_ (
    .CLK(CLK_bF$buf142),
    .D(\datapath.csr.csr_wdata [9]),
    .Q(\datapath.regcsrwb [9])
);

DFFPOSX1 _10426_ (
    .CLK(CLK_bF$buf141),
    .D(\datapath.csr.csr_wdata [10]),
    .Q(\datapath.regcsrwb [10])
);

DFFPOSX1 _10427_ (
    .CLK(CLK_bF$buf140),
    .D(\datapath.csr.csr_wdata [11]),
    .Q(\datapath.regcsrwb [11])
);

DFFPOSX1 _10428_ (
    .CLK(CLK_bF$buf139),
    .D(\datapath.csr.csr_wdata [12]),
    .Q(\datapath.regcsrwb [12])
);

DFFPOSX1 _10429_ (
    .CLK(CLK_bF$buf138),
    .D(\datapath.csr.csr_wdata [13]),
    .Q(\datapath.regcsrwb [13])
);

DFFPOSX1 _10430_ (
    .CLK(CLK_bF$buf137),
    .D(\datapath.csr.csr_wdata [14]),
    .Q(\datapath.regcsrwb [14])
);

DFFPOSX1 _10431_ (
    .CLK(CLK_bF$buf136),
    .D(\datapath.csr.csr_wdata [15]),
    .Q(\datapath.regcsrwb [15])
);

DFFPOSX1 _10432_ (
    .CLK(CLK_bF$buf135),
    .D(\datapath.csr.csr_wdata [16]),
    .Q(\datapath.regcsrwb [16])
);

DFFPOSX1 _10433_ (
    .CLK(CLK_bF$buf134),
    .D(\datapath.csr.csr_wdata [17]),
    .Q(\datapath.regcsrwb [17])
);

DFFPOSX1 _10434_ (
    .CLK(CLK_bF$buf133),
    .D(\datapath.csr.csr_wdata [18]),
    .Q(\datapath.regcsrwb [18])
);

DFFPOSX1 _10435_ (
    .CLK(CLK_bF$buf132),
    .D(\datapath.csr.csr_wdata [19]),
    .Q(\datapath.regcsrwb [19])
);

DFFPOSX1 _10436_ (
    .CLK(CLK_bF$buf131),
    .D(\datapath.csr.csr_wdata [20]),
    .Q(\datapath.regcsrwb [20])
);

DFFPOSX1 _10437_ (
    .CLK(CLK_bF$buf130),
    .D(\datapath.csr.csr_wdata [21]),
    .Q(\datapath.regcsrwb [21])
);

DFFPOSX1 _10438_ (
    .CLK(CLK_bF$buf129),
    .D(\datapath.csr.csr_wdata [22]),
    .Q(\datapath.regcsrwb [22])
);

DFFPOSX1 _10439_ (
    .CLK(CLK_bF$buf128),
    .D(\datapath.csr.csr_wdata [23]),
    .Q(\datapath.regcsrwb [23])
);

DFFPOSX1 _10440_ (
    .CLK(CLK_bF$buf127),
    .D(\datapath.csr.csr_wdata [24]),
    .Q(\datapath.regcsrwb [24])
);

DFFPOSX1 _10441_ (
    .CLK(CLK_bF$buf126),
    .D(\datapath.csr.csr_wdata [25]),
    .Q(\datapath.regcsrwb [25])
);

DFFPOSX1 _10442_ (
    .CLK(CLK_bF$buf125),
    .D(\datapath.csr.csr_wdata [26]),
    .Q(\datapath.regcsrwb [26])
);

DFFPOSX1 _10443_ (
    .CLK(CLK_bF$buf124),
    .D(\datapath.csr.csr_wdata [27]),
    .Q(\datapath.regcsrwb [27])
);

DFFPOSX1 _10444_ (
    .CLK(CLK_bF$buf123),
    .D(\datapath.csr.csr_wdata [28]),
    .Q(\datapath.regcsrwb [28])
);

DFFPOSX1 _10445_ (
    .CLK(CLK_bF$buf122),
    .D(\datapath.csr.csr_wdata [29]),
    .Q(\datapath.regcsrwb [29])
);

DFFPOSX1 _10446_ (
    .CLK(CLK_bF$buf121),
    .D(\datapath.csr.csr_wdata [30]),
    .Q(\datapath.regcsrwb [30])
);

DFFPOSX1 _10447_ (
    .CLK(CLK_bF$buf120),
    .D(\datapath.csr.csr_wdata [31]),
    .Q(\datapath.regcsrwb [31])
);

DFFPOSX1 _10448_ (
    .CLK(CLK_bF$buf119),
    .D(\datapath.memdataload [0]),
    .Q(\datapath.regloadwb [0])
);

DFFPOSX1 _10449_ (
    .CLK(CLK_bF$buf118),
    .D(\datapath.memdataload [1]),
    .Q(\datapath.regloadwb [1])
);

DFFPOSX1 _10450_ (
    .CLK(CLK_bF$buf117),
    .D(\datapath.memdataload [2]),
    .Q(\datapath.regloadwb [2])
);

DFFPOSX1 _10451_ (
    .CLK(CLK_bF$buf116),
    .D(\datapath.memdataload [3]),
    .Q(\datapath.regloadwb [3])
);

DFFPOSX1 _10452_ (
    .CLK(CLK_bF$buf115),
    .D(\datapath.memdataload [4]),
    .Q(\datapath.regloadwb [4])
);

DFFPOSX1 _10453_ (
    .CLK(CLK_bF$buf114),
    .D(\datapath.memdataload [5]),
    .Q(\datapath.regloadwb [5])
);

DFFPOSX1 _10454_ (
    .CLK(CLK_bF$buf113),
    .D(\datapath.memdataload [6]),
    .Q(\datapath.regloadwb [6])
);

DFFPOSX1 _10455_ (
    .CLK(CLK_bF$buf112),
    .D(\datapath.memdataload [7]),
    .Q(\datapath.regloadwb [7])
);

DFFPOSX1 _10456_ (
    .CLK(CLK_bF$buf111),
    .D(\datapath.memdataload [8]),
    .Q(\datapath.regloadwb [8])
);

DFFPOSX1 _10457_ (
    .CLK(CLK_bF$buf110),
    .D(\datapath.memdataload [9]),
    .Q(\datapath.regloadwb [9])
);

DFFPOSX1 _10458_ (
    .CLK(CLK_bF$buf109),
    .D(\datapath.memdataload [10]),
    .Q(\datapath.regloadwb [10])
);

DFFPOSX1 _10459_ (
    .CLK(CLK_bF$buf108),
    .D(\datapath.memdataload [11]),
    .Q(\datapath.regloadwb [11])
);

DFFPOSX1 _10460_ (
    .CLK(CLK_bF$buf107),
    .D(\datapath.memdataload [12]),
    .Q(\datapath.regloadwb [12])
);

DFFPOSX1 _10461_ (
    .CLK(CLK_bF$buf106),
    .D(\datapath.memdataload [13]),
    .Q(\datapath.regloadwb [13])
);

DFFPOSX1 _10462_ (
    .CLK(CLK_bF$buf105),
    .D(\datapath.memdataload [14]),
    .Q(\datapath.regloadwb [14])
);

DFFPOSX1 _10463_ (
    .CLK(CLK_bF$buf104),
    .D(\datapath.memdataload [15]),
    .Q(\datapath.regloadwb [15])
);

DFFPOSX1 _10464_ (
    .CLK(CLK_bF$buf103),
    .D(\datapath.memdataload [16]),
    .Q(\datapath.regloadwb [16])
);

DFFPOSX1 _10465_ (
    .CLK(CLK_bF$buf102),
    .D(\datapath.memdataload [17]),
    .Q(\datapath.regloadwb [17])
);

DFFPOSX1 _10466_ (
    .CLK(CLK_bF$buf101),
    .D(\datapath.memdataload [18]),
    .Q(\datapath.regloadwb [18])
);

DFFPOSX1 _10467_ (
    .CLK(CLK_bF$buf100),
    .D(\datapath.memdataload [19]),
    .Q(\datapath.regloadwb [19])
);

DFFPOSX1 _10468_ (
    .CLK(CLK_bF$buf99),
    .D(\datapath.memdataload [20]),
    .Q(\datapath.regloadwb [20])
);

DFFPOSX1 _10469_ (
    .CLK(CLK_bF$buf98),
    .D(\datapath.memdataload [21]),
    .Q(\datapath.regloadwb [21])
);

DFFPOSX1 _10470_ (
    .CLK(CLK_bF$buf97),
    .D(\datapath.memdataload [22]),
    .Q(\datapath.regloadwb [22])
);

DFFPOSX1 _10471_ (
    .CLK(CLK_bF$buf96),
    .D(\datapath.memdataload [23]),
    .Q(\datapath.regloadwb [23])
);

DFFPOSX1 _10472_ (
    .CLK(CLK_bF$buf95),
    .D(\datapath.memdataload [24]),
    .Q(\datapath.regloadwb [24])
);

DFFPOSX1 _10473_ (
    .CLK(CLK_bF$buf94),
    .D(\datapath.memdataload [25]),
    .Q(\datapath.regloadwb [25])
);

DFFPOSX1 _10474_ (
    .CLK(CLK_bF$buf93),
    .D(\datapath.memdataload [26]),
    .Q(\datapath.regloadwb [26])
);

DFFPOSX1 _10475_ (
    .CLK(CLK_bF$buf92),
    .D(\datapath.memdataload [27]),
    .Q(\datapath.regloadwb [27])
);

DFFPOSX1 _10476_ (
    .CLK(CLK_bF$buf91),
    .D(\datapath.memdataload [28]),
    .Q(\datapath.regloadwb [28])
);

DFFPOSX1 _10477_ (
    .CLK(CLK_bF$buf90),
    .D(\datapath.memdataload [29]),
    .Q(\datapath.regloadwb [29])
);

DFFPOSX1 _10478_ (
    .CLK(CLK_bF$buf89),
    .D(\datapath.memdataload [30]),
    .Q(\datapath.regloadwb [30])
);

DFFPOSX1 _10479_ (
    .CLK(CLK_bF$buf88),
    .D(\datapath.memdataload [31]),
    .Q(\datapath.regloadwb [31])
);

DFFPOSX1 _10480_ (
    .CLK(CLK_bF$buf87),
    .D(_0__0_bF$buf4),
    .Q(\datapath.regcwb [0])
);

DFFPOSX1 _10481_ (
    .CLK(CLK_bF$buf86),
    .D(_0__1_bF$buf10),
    .Q(\datapath.regcwb [1])
);

DFFPOSX1 _10482_ (
    .CLK(CLK_bF$buf85),
    .D(_0_[2]),
    .Q(\datapath.regcwb [2])
);

DFFPOSX1 _10483_ (
    .CLK(CLK_bF$buf84),
    .D(_0_[3]),
    .Q(\datapath.regcwb [3])
);

DFFPOSX1 _10484_ (
    .CLK(CLK_bF$buf83),
    .D(_0_[4]),
    .Q(\datapath.regcwb [4])
);

DFFPOSX1 _10485_ (
    .CLK(CLK_bF$buf82),
    .D(_0_[5]),
    .Q(\datapath.regcwb [5])
);

DFFPOSX1 _10486_ (
    .CLK(CLK_bF$buf81),
    .D(_0_[6]),
    .Q(\datapath.regcwb [6])
);

DFFPOSX1 _10487_ (
    .CLK(CLK_bF$buf80),
    .D(_0_[7]),
    .Q(\datapath.regcwb [7])
);

DFFPOSX1 _10488_ (
    .CLK(CLK_bF$buf79),
    .D(_0_[8]),
    .Q(\datapath.regcwb [8])
);

DFFPOSX1 _10489_ (
    .CLK(CLK_bF$buf78),
    .D(_0_[9]),
    .Q(\datapath.regcwb [9])
);

DFFPOSX1 _10490_ (
    .CLK(CLK_bF$buf77),
    .D(_0_[10]),
    .Q(\datapath.regcwb [10])
);

DFFPOSX1 _10491_ (
    .CLK(CLK_bF$buf76),
    .D(_0_[11]),
    .Q(\datapath.regcwb [11])
);

DFFPOSX1 _10492_ (
    .CLK(CLK_bF$buf75),
    .D(_0_[12]),
    .Q(\datapath.regcwb [12])
);

DFFPOSX1 _10493_ (
    .CLK(CLK_bF$buf74),
    .D(_0_[13]),
    .Q(\datapath.regcwb [13])
);

DFFPOSX1 _10494_ (
    .CLK(CLK_bF$buf73),
    .D(_0_[14]),
    .Q(\datapath.regcwb [14])
);

DFFPOSX1 _10495_ (
    .CLK(CLK_bF$buf72),
    .D(_0_[15]),
    .Q(\datapath.regcwb [15])
);

DFFPOSX1 _10496_ (
    .CLK(CLK_bF$buf71),
    .D(_0_[16]),
    .Q(\datapath.regcwb [16])
);

DFFPOSX1 _10497_ (
    .CLK(CLK_bF$buf70),
    .D(_0_[17]),
    .Q(\datapath.regcwb [17])
);

DFFPOSX1 _10498_ (
    .CLK(CLK_bF$buf69),
    .D(_0_[18]),
    .Q(\datapath.regcwb [18])
);

DFFPOSX1 _10499_ (
    .CLK(CLK_bF$buf68),
    .D(_0_[19]),
    .Q(\datapath.regcwb [19])
);

DFFPOSX1 _10500_ (
    .CLK(CLK_bF$buf67),
    .D(_0_[20]),
    .Q(\datapath.regcwb [20])
);

DFFPOSX1 _10501_ (
    .CLK(CLK_bF$buf66),
    .D(_0_[21]),
    .Q(\datapath.regcwb [21])
);

DFFPOSX1 _10502_ (
    .CLK(CLK_bF$buf65),
    .D(_0_[22]),
    .Q(\datapath.regcwb [22])
);

DFFPOSX1 _10503_ (
    .CLK(CLK_bF$buf64),
    .D(_0_[23]),
    .Q(\datapath.regcwb [23])
);

DFFPOSX1 _10504_ (
    .CLK(CLK_bF$buf63),
    .D(_0_[24]),
    .Q(\datapath.regcwb [24])
);

DFFPOSX1 _10505_ (
    .CLK(CLK_bF$buf62),
    .D(_0_[25]),
    .Q(\datapath.regcwb [25])
);

DFFPOSX1 _10506_ (
    .CLK(CLK_bF$buf61),
    .D(_0_[26]),
    .Q(\datapath.regcwb [26])
);

DFFPOSX1 _10507_ (
    .CLK(CLK_bF$buf60),
    .D(_0_[27]),
    .Q(\datapath.regcwb [27])
);

DFFPOSX1 _10508_ (
    .CLK(CLK_bF$buf59),
    .D(_0_[28]),
    .Q(\datapath.regcwb [28])
);

DFFPOSX1 _10509_ (
    .CLK(CLK_bF$buf58),
    .D(_0_[29]),
    .Q(\datapath.regcwb [29])
);

DFFPOSX1 _10510_ (
    .CLK(CLK_bF$buf57),
    .D(_0_[30]),
    .Q(\datapath.regcwb [30])
);

DFFPOSX1 _10511_ (
    .CLK(CLK_bF$buf56),
    .D(_0_[31]),
    .Q(\datapath.regcwb [31])
);

DFFPOSX1 _10512_ (
    .CLK(CLK_bF$buf55),
    .D(\controlunit.csrfile_trap_wen_bF$buf6 ),
    .Q(\datapath.regwbtrap )
);

DFFPOSX1 _10513_ (
    .CLK(CLK_bF$buf54),
    .D(\controlunit.mret_bF$buf4 ),
    .Q(\datapath.regmret )
);

DFFPOSX1 _10514_ (
    .CLK(CLK_bF$buf53),
    .D(\datapath.meminstr [0]),
    .Q(\datapath.wbinstr [0])
);

DFFPOSX1 _10515_ (
    .CLK(CLK_bF$buf52),
    .D(\datapath.meminstr [1]),
    .Q(\datapath.wbinstr [1])
);

DFFPOSX1 _10516_ (
    .CLK(CLK_bF$buf51),
    .D(\datapath.meminstr [2]),
    .Q(\datapath.wbinstr [2])
);

DFFPOSX1 _10517_ (
    .CLK(CLK_bF$buf50),
    .D(\datapath.meminstr [3]),
    .Q(\datapath.wbinstr [3])
);

DFFPOSX1 _10518_ (
    .CLK(CLK_bF$buf49),
    .D(\datapath.meminstr [4]),
    .Q(\datapath.wbinstr [4])
);

DFFPOSX1 _10519_ (
    .CLK(CLK_bF$buf48),
    .D(\datapath.meminstr [5]),
    .Q(\datapath.wbinstr [5])
);

DFFPOSX1 _10520_ (
    .CLK(CLK_bF$buf47),
    .D(\datapath.meminstr [6]),
    .Q(\datapath.wbinstr [6])
);

DFFPOSX1 _10521_ (
    .CLK(CLK_bF$buf46),
    .D(\datapath.meminstr [7]),
    .Q(\datapath.wbinstr [7])
);

DFFPOSX1 _10522_ (
    .CLK(CLK_bF$buf45),
    .D(\datapath.meminstr [8]),
    .Q(\datapath.wbinstr [8])
);

DFFPOSX1 _10523_ (
    .CLK(CLK_bF$buf44),
    .D(\datapath.meminstr [9]),
    .Q(\datapath.wbinstr [9])
);

DFFPOSX1 _10524_ (
    .CLK(CLK_bF$buf43),
    .D(\datapath.meminstr [10]),
    .Q(\datapath.wbinstr [10])
);

DFFPOSX1 _10525_ (
    .CLK(CLK_bF$buf42),
    .D(\datapath.meminstr [11]),
    .Q(\datapath.wbinstr [11])
);

DFFPOSX1 _10526_ (
    .CLK(CLK_bF$buf41),
    .D(\datapath.meminstr [12]),
    .Q(\datapath.wbinstr [12])
);

DFFPOSX1 _10527_ (
    .CLK(CLK_bF$buf40),
    .D(\datapath.meminstr [13]),
    .Q(\datapath.wbinstr [13])
);

DFFPOSX1 _10528_ (
    .CLK(CLK_bF$buf39),
    .D(\datapath.meminstr [14]),
    .Q(\datapath.wbinstr [14])
);

DFFPOSX1 _10529_ (
    .CLK(CLK_bF$buf38),
    .D(\datapath.mempc_4 [0]),
    .Q(\datapath.wbpc_4 [0])
);

DFFPOSX1 _10530_ (
    .CLK(CLK_bF$buf37),
    .D(\datapath.mempc_4 [1]),
    .Q(\datapath.wbpc_4 [1])
);

DFFPOSX1 _10531_ (
    .CLK(CLK_bF$buf36),
    .D(\datapath.mempc_4 [2]),
    .Q(\datapath.wbpc_4 [2])
);

DFFPOSX1 _10532_ (
    .CLK(CLK_bF$buf35),
    .D(\datapath.mempc_4 [3]),
    .Q(\datapath.wbpc_4 [3])
);

DFFPOSX1 _10533_ (
    .CLK(CLK_bF$buf34),
    .D(\datapath.mempc_4 [4]),
    .Q(\datapath.wbpc_4 [4])
);

DFFPOSX1 _10534_ (
    .CLK(CLK_bF$buf33),
    .D(\datapath.mempc_4 [5]),
    .Q(\datapath.wbpc_4 [5])
);

DFFPOSX1 _10535_ (
    .CLK(CLK_bF$buf32),
    .D(\datapath.mempc_4 [6]),
    .Q(\datapath.wbpc_4 [6])
);

DFFPOSX1 _10536_ (
    .CLK(CLK_bF$buf31),
    .D(\datapath.mempc_4 [7]),
    .Q(\datapath.wbpc_4 [7])
);

DFFPOSX1 _10537_ (
    .CLK(CLK_bF$buf30),
    .D(\datapath.mempc_4 [8]),
    .Q(\datapath.wbpc_4 [8])
);

DFFPOSX1 _10538_ (
    .CLK(CLK_bF$buf29),
    .D(\datapath.mempc_4 [9]),
    .Q(\datapath.wbpc_4 [9])
);

DFFPOSX1 _10539_ (
    .CLK(CLK_bF$buf28),
    .D(\datapath.mempc_4 [10]),
    .Q(\datapath.wbpc_4 [10])
);

DFFPOSX1 _10540_ (
    .CLK(CLK_bF$buf27),
    .D(\datapath.mempc_4 [11]),
    .Q(\datapath.wbpc_4 [11])
);

DFFPOSX1 _10541_ (
    .CLK(CLK_bF$buf26),
    .D(\datapath.mempc_4 [12]),
    .Q(\datapath.wbpc_4 [12])
);

DFFPOSX1 _10542_ (
    .CLK(CLK_bF$buf25),
    .D(\datapath.mempc_4 [13]),
    .Q(\datapath.wbpc_4 [13])
);

DFFPOSX1 _10543_ (
    .CLK(CLK_bF$buf24),
    .D(\datapath.mempc_4 [14]),
    .Q(\datapath.wbpc_4 [14])
);

DFFPOSX1 _10544_ (
    .CLK(CLK_bF$buf23),
    .D(\datapath.mempc_4 [15]),
    .Q(\datapath.wbpc_4 [15])
);

DFFPOSX1 _10545_ (
    .CLK(CLK_bF$buf22),
    .D(\datapath.mempc_4 [16]),
    .Q(\datapath.wbpc_4 [16])
);

DFFPOSX1 _10546_ (
    .CLK(CLK_bF$buf21),
    .D(\datapath.mempc_4 [17]),
    .Q(\datapath.wbpc_4 [17])
);

DFFPOSX1 _10547_ (
    .CLK(CLK_bF$buf20),
    .D(\datapath.mempc_4 [18]),
    .Q(\datapath.wbpc_4 [18])
);

DFFPOSX1 _10548_ (
    .CLK(CLK_bF$buf19),
    .D(\datapath.mempc_4 [19]),
    .Q(\datapath.wbpc_4 [19])
);

DFFPOSX1 _10549_ (
    .CLK(CLK_bF$buf18),
    .D(\datapath.mempc_4 [20]),
    .Q(\datapath.wbpc_4 [20])
);

DFFPOSX1 _10550_ (
    .CLK(CLK_bF$buf17),
    .D(\datapath.mempc_4 [21]),
    .Q(\datapath.wbpc_4 [21])
);

DFFPOSX1 _10551_ (
    .CLK(CLK_bF$buf16),
    .D(\datapath.mempc_4 [22]),
    .Q(\datapath.wbpc_4 [22])
);

DFFPOSX1 _10552_ (
    .CLK(CLK_bF$buf15),
    .D(\datapath.mempc_4 [23]),
    .Q(\datapath.wbpc_4 [23])
);

DFFPOSX1 _10553_ (
    .CLK(CLK_bF$buf14),
    .D(\datapath.mempc_4 [24]),
    .Q(\datapath.wbpc_4 [24])
);

DFFPOSX1 _10554_ (
    .CLK(CLK_bF$buf13),
    .D(\datapath.mempc_4 [25]),
    .Q(\datapath.wbpc_4 [25])
);

DFFPOSX1 _10555_ (
    .CLK(CLK_bF$buf12),
    .D(\datapath.mempc_4 [26]),
    .Q(\datapath.wbpc_4 [26])
);

DFFPOSX1 _10556_ (
    .CLK(CLK_bF$buf11),
    .D(\datapath.mempc_4 [27]),
    .Q(\datapath.wbpc_4 [27])
);

DFFPOSX1 _10557_ (
    .CLK(CLK_bF$buf10),
    .D(\datapath.mempc_4 [28]),
    .Q(\datapath.wbpc_4 [28])
);

DFFPOSX1 _10558_ (
    .CLK(CLK_bF$buf9),
    .D(\datapath.mempc_4 [29]),
    .Q(\datapath.wbpc_4 [29])
);

DFFPOSX1 _10559_ (
    .CLK(CLK_bF$buf8),
    .D(\datapath.mempc_4 [30]),
    .Q(\datapath.wbpc_4 [30])
);

DFFPOSX1 _10560_ (
    .CLK(CLK_bF$buf7),
    .D(\datapath.mempc_4 [31]),
    .Q(\datapath.wbpc_4 [31])
);

DFFPOSX1 _10561_ (
    .CLK(CLK_bF$buf6),
    .D(\datapath.jumptarget [1]),
    .Q(\datapath.programcounter.jumps [1])
);

DFFPOSX1 _10562_ (
    .CLK(CLK_bF$buf5),
    .D(\datapath.jumptarget [2]),
    .Q(\datapath.programcounter.jumps [2])
);

DFFPOSX1 _10563_ (
    .CLK(CLK_bF$buf4),
    .D(\datapath.jumptarget [3]),
    .Q(\datapath.programcounter.jumps [3])
);

DFFPOSX1 _10564_ (
    .CLK(CLK_bF$buf3),
    .D(\datapath.jumptarget [4]),
    .Q(\datapath.programcounter.jumps [4])
);

DFFPOSX1 _10565_ (
    .CLK(CLK_bF$buf2),
    .D(\datapath.jumptarget [5]),
    .Q(\datapath.programcounter.jumps [5])
);

DFFPOSX1 _10566_ (
    .CLK(CLK_bF$buf1),
    .D(\datapath.jumptarget [6]),
    .Q(\datapath.programcounter.jumps [6])
);

DFFPOSX1 _10567_ (
    .CLK(CLK_bF$buf0),
    .D(\datapath.jumptarget [7]),
    .Q(\datapath.programcounter.jumps [7])
);

DFFPOSX1 _10568_ (
    .CLK(CLK_bF$buf151),
    .D(\datapath.jumptarget [8]),
    .Q(\datapath.programcounter.jumps [8])
);

DFFPOSX1 _10569_ (
    .CLK(CLK_bF$buf150),
    .D(\datapath.jumptarget [9]),
    .Q(\datapath.programcounter.jumps [9])
);

DFFPOSX1 _10570_ (
    .CLK(CLK_bF$buf149),
    .D(\datapath.jumptarget [10]),
    .Q(\datapath.programcounter.jumps [10])
);

DFFPOSX1 _10571_ (
    .CLK(CLK_bF$buf148),
    .D(\datapath.jumptarget [11]),
    .Q(\datapath.programcounter.jumps [11])
);

DFFPOSX1 _10572_ (
    .CLK(CLK_bF$buf147),
    .D(\datapath.jumptarget [12]),
    .Q(\datapath.programcounter.jumps [12])
);

DFFPOSX1 _10573_ (
    .CLK(CLK_bF$buf146),
    .D(\datapath.jumptarget [13]),
    .Q(\datapath.programcounter.jumps [13])
);

DFFPOSX1 _10574_ (
    .CLK(CLK_bF$buf145),
    .D(\datapath.jumptarget [14]),
    .Q(\datapath.programcounter.jumps [14])
);

DFFPOSX1 _10575_ (
    .CLK(CLK_bF$buf144),
    .D(\datapath.jumptarget [15]),
    .Q(\datapath.programcounter.jumps [15])
);

DFFPOSX1 _10576_ (
    .CLK(CLK_bF$buf143),
    .D(\datapath.jumptarget [16]),
    .Q(\datapath.programcounter.jumps [16])
);

DFFPOSX1 _10577_ (
    .CLK(CLK_bF$buf142),
    .D(\datapath.jumptarget [17]),
    .Q(\datapath.programcounter.jumps [17])
);

DFFPOSX1 _10578_ (
    .CLK(CLK_bF$buf141),
    .D(\datapath.jumptarget [18]),
    .Q(\datapath.programcounter.jumps [18])
);

DFFPOSX1 _10579_ (
    .CLK(CLK_bF$buf140),
    .D(\datapath.jumptarget [19]),
    .Q(\datapath.programcounter.jumps [19])
);

DFFPOSX1 _10580_ (
    .CLK(CLK_bF$buf139),
    .D(\datapath.jumptarget [20]),
    .Q(\datapath.programcounter.jumps [20])
);

DFFPOSX1 _10581_ (
    .CLK(CLK_bF$buf138),
    .D(\datapath.jumptarget [21]),
    .Q(\datapath.programcounter.jumps [21])
);

DFFPOSX1 _10582_ (
    .CLK(CLK_bF$buf137),
    .D(\datapath.jumptarget [22]),
    .Q(\datapath.programcounter.jumps [22])
);

DFFPOSX1 _10583_ (
    .CLK(CLK_bF$buf136),
    .D(\datapath.jumptarget [23]),
    .Q(\datapath.programcounter.jumps [23])
);

DFFPOSX1 _10584_ (
    .CLK(CLK_bF$buf135),
    .D(\datapath.jumptarget [24]),
    .Q(\datapath.programcounter.jumps [24])
);

DFFPOSX1 _10585_ (
    .CLK(CLK_bF$buf134),
    .D(\datapath.jumptarget [25]),
    .Q(\datapath.programcounter.jumps [25])
);

DFFPOSX1 _10586_ (
    .CLK(CLK_bF$buf133),
    .D(\datapath.jumptarget [26]),
    .Q(\datapath.programcounter.jumps [26])
);

DFFPOSX1 _10587_ (
    .CLK(CLK_bF$buf132),
    .D(\datapath.jumptarget [27]),
    .Q(\datapath.programcounter.jumps [27])
);

DFFPOSX1 _10588_ (
    .CLK(CLK_bF$buf131),
    .D(\datapath.jumptarget [28]),
    .Q(\datapath.programcounter.jumps [28])
);

DFFPOSX1 _10589_ (
    .CLK(CLK_bF$buf130),
    .D(\datapath.jumptarget [29]),
    .Q(\datapath.programcounter.jumps [29])
);

DFFPOSX1 _10590_ (
    .CLK(CLK_bF$buf129),
    .D(\datapath.jumptarget [30]),
    .Q(\datapath.programcounter.jumps [30])
);

DFFPOSX1 _10591_ (
    .CLK(CLK_bF$buf128),
    .D(\datapath.jumptarget [31]),
    .Q(\datapath.programcounter.jumps [31])
);

DFFPOSX1 _10592_ (
    .CLK(CLK_bF$buf127),
    .D(\datapath.regcsralu [0]),
    .Q(\datapath.csr.csr_wdata [0])
);

DFFPOSX1 _10593_ (
    .CLK(CLK_bF$buf126),
    .D(\datapath.regcsralu [1]),
    .Q(\datapath.csr.csr_wdata [1])
);

DFFPOSX1 _10594_ (
    .CLK(CLK_bF$buf125),
    .D(\datapath.regcsralu [2]),
    .Q(\datapath.csr.csr_wdata [2])
);

DFFPOSX1 _10595_ (
    .CLK(CLK_bF$buf124),
    .D(\datapath.regcsralu [3]),
    .Q(\datapath.csr.csr_wdata [3])
);

DFFPOSX1 _10596_ (
    .CLK(CLK_bF$buf123),
    .D(\datapath.regcsralu [4]),
    .Q(\datapath.csr.csr_wdata [4])
);

DFFPOSX1 _10597_ (
    .CLK(CLK_bF$buf122),
    .D(\datapath.regcsralu [5]),
    .Q(\datapath.csr.csr_wdata [5])
);

DFFPOSX1 _10598_ (
    .CLK(CLK_bF$buf121),
    .D(\datapath.regcsralu [6]),
    .Q(\datapath.csr.csr_wdata [6])
);

DFFPOSX1 _10599_ (
    .CLK(CLK_bF$buf120),
    .D(\datapath.regcsralu [7]),
    .Q(\datapath.csr.csr_wdata [7])
);

DFFPOSX1 _10600_ (
    .CLK(CLK_bF$buf119),
    .D(\datapath.regcsralu [8]),
    .Q(\datapath.csr.csr_wdata [8])
);

DFFPOSX1 _10601_ (
    .CLK(CLK_bF$buf118),
    .D(\datapath.regcsralu [9]),
    .Q(\datapath.csr.csr_wdata [9])
);

DFFPOSX1 _10602_ (
    .CLK(CLK_bF$buf117),
    .D(\datapath.regcsralu [10]),
    .Q(\datapath.csr.csr_wdata [10])
);

DFFPOSX1 _10603_ (
    .CLK(CLK_bF$buf116),
    .D(\datapath.regcsralu [11]),
    .Q(\datapath.csr.csr_wdata [11])
);

DFFPOSX1 _10604_ (
    .CLK(CLK_bF$buf115),
    .D(\datapath.regcsralu [12]),
    .Q(\datapath.csr.csr_wdata [12])
);

DFFPOSX1 _10605_ (
    .CLK(CLK_bF$buf114),
    .D(\datapath.regcsralu [13]),
    .Q(\datapath.csr.csr_wdata [13])
);

DFFPOSX1 _10606_ (
    .CLK(CLK_bF$buf113),
    .D(\datapath.regcsralu [14]),
    .Q(\datapath.csr.csr_wdata [14])
);

DFFPOSX1 _10607_ (
    .CLK(CLK_bF$buf112),
    .D(\datapath.regcsralu [15]),
    .Q(\datapath.csr.csr_wdata [15])
);

DFFPOSX1 _10608_ (
    .CLK(CLK_bF$buf111),
    .D(\datapath.regcsralu [16]),
    .Q(\datapath.csr.csr_wdata [16])
);

DFFPOSX1 _10609_ (
    .CLK(CLK_bF$buf110),
    .D(\datapath.regcsralu [17]),
    .Q(\datapath.csr.csr_wdata [17])
);

DFFPOSX1 _10610_ (
    .CLK(CLK_bF$buf109),
    .D(\datapath.regcsralu [18]),
    .Q(\datapath.csr.csr_wdata [18])
);

DFFPOSX1 _10611_ (
    .CLK(CLK_bF$buf108),
    .D(\datapath.regcsralu [19]),
    .Q(\datapath.csr.csr_wdata [19])
);

DFFPOSX1 _10612_ (
    .CLK(CLK_bF$buf107),
    .D(\datapath.regcsralu [20]),
    .Q(\datapath.csr.csr_wdata [20])
);

DFFPOSX1 _10613_ (
    .CLK(CLK_bF$buf106),
    .D(\datapath.regcsralu [21]),
    .Q(\datapath.csr.csr_wdata [21])
);

DFFPOSX1 _10614_ (
    .CLK(CLK_bF$buf105),
    .D(\datapath.regcsralu [22]),
    .Q(\datapath.csr.csr_wdata [22])
);

DFFPOSX1 _10615_ (
    .CLK(CLK_bF$buf104),
    .D(\datapath.regcsralu [23]),
    .Q(\datapath.csr.csr_wdata [23])
);

DFFPOSX1 _10616_ (
    .CLK(CLK_bF$buf103),
    .D(\datapath.regcsralu [24]),
    .Q(\datapath.csr.csr_wdata [24])
);

DFFPOSX1 _10617_ (
    .CLK(CLK_bF$buf102),
    .D(\datapath.regcsralu [25]),
    .Q(\datapath.csr.csr_wdata [25])
);

DFFPOSX1 _10618_ (
    .CLK(CLK_bF$buf101),
    .D(\datapath.regcsralu [26]),
    .Q(\datapath.csr.csr_wdata [26])
);

DFFPOSX1 _10619_ (
    .CLK(CLK_bF$buf100),
    .D(\datapath.regcsralu [27]),
    .Q(\datapath.csr.csr_wdata [27])
);

DFFPOSX1 _10620_ (
    .CLK(CLK_bF$buf99),
    .D(\datapath.regcsralu [28]),
    .Q(\datapath.csr.csr_wdata [28])
);

DFFPOSX1 _10621_ (
    .CLK(CLK_bF$buf98),
    .D(\datapath.regcsralu [29]),
    .Q(\datapath.csr.csr_wdata [29])
);

DFFPOSX1 _10622_ (
    .CLK(CLK_bF$buf97),
    .D(\datapath.regcsralu [30]),
    .Q(\datapath.csr.csr_wdata [30])
);

DFFPOSX1 _10623_ (
    .CLK(CLK_bF$buf96),
    .D(\datapath.regcsralu [31]),
    .Q(\datapath.csr.csr_wdata [31])
);

DFFPOSX1 _10624_ (
    .CLK(CLK_bF$buf95),
    .D(\datapath.regrs2alu [0]),
    .Q(\datapath.memoryinterface.data_store [0])
);

DFFPOSX1 _10625_ (
    .CLK(CLK_bF$buf94),
    .D(\datapath.regrs2alu [1]),
    .Q(\datapath.memoryinterface.data_store [1])
);

DFFPOSX1 _10626_ (
    .CLK(CLK_bF$buf93),
    .D(\datapath.regrs2alu [2]),
    .Q(\datapath.memoryinterface.data_store [2])
);

DFFPOSX1 _10627_ (
    .CLK(CLK_bF$buf92),
    .D(\datapath.regrs2alu [3]),
    .Q(\datapath.memoryinterface.data_store [3])
);

DFFPOSX1 _10628_ (
    .CLK(CLK_bF$buf91),
    .D(\datapath.regrs2alu [4]),
    .Q(\datapath.memoryinterface.data_store [4])
);

DFFPOSX1 _10629_ (
    .CLK(CLK_bF$buf90),
    .D(\datapath.regrs2alu [5]),
    .Q(\datapath.memoryinterface.data_store [5])
);

DFFPOSX1 _10630_ (
    .CLK(CLK_bF$buf89),
    .D(\datapath.regrs2alu [6]),
    .Q(\datapath.memoryinterface.data_store [6])
);

DFFPOSX1 _10631_ (
    .CLK(CLK_bF$buf88),
    .D(\datapath.regrs2alu [7]),
    .Q(\datapath.memoryinterface.data_store [7])
);

DFFPOSX1 _10632_ (
    .CLK(CLK_bF$buf87),
    .D(\datapath.regrs2alu [8]),
    .Q(\datapath.memoryinterface.data_store [8])
);

DFFPOSX1 _10633_ (
    .CLK(CLK_bF$buf86),
    .D(\datapath.regrs2alu [9]),
    .Q(\datapath.memoryinterface.data_store [9])
);

DFFPOSX1 _10634_ (
    .CLK(CLK_bF$buf85),
    .D(\datapath.regrs2alu [10]),
    .Q(\datapath.memoryinterface.data_store [10])
);

DFFPOSX1 _10635_ (
    .CLK(CLK_bF$buf84),
    .D(\datapath.regrs2alu [11]),
    .Q(\datapath.memoryinterface.data_store [11])
);

DFFPOSX1 _10636_ (
    .CLK(CLK_bF$buf83),
    .D(\datapath.regrs2alu [12]),
    .Q(\datapath.memoryinterface.data_store [12])
);

DFFPOSX1 _10637_ (
    .CLK(CLK_bF$buf82),
    .D(\datapath.regrs2alu [13]),
    .Q(\datapath.memoryinterface.data_store [13])
);

DFFPOSX1 _10638_ (
    .CLK(CLK_bF$buf81),
    .D(\datapath.regrs2alu [14]),
    .Q(\datapath.memoryinterface.data_store [14])
);

DFFPOSX1 _10639_ (
    .CLK(CLK_bF$buf80),
    .D(\datapath.regrs2alu [15]),
    .Q(\datapath.memoryinterface.data_store [15])
);

DFFPOSX1 _10640_ (
    .CLK(CLK_bF$buf79),
    .D(\datapath.regrs2alu [16]),
    .Q(\datapath.memoryinterface.data_store [16])
);

DFFPOSX1 _10641_ (
    .CLK(CLK_bF$buf78),
    .D(\datapath.regrs2alu [17]),
    .Q(\datapath.memoryinterface.data_store [17])
);

DFFPOSX1 _10642_ (
    .CLK(CLK_bF$buf77),
    .D(\datapath.regrs2alu [18]),
    .Q(\datapath.memoryinterface.data_store [18])
);

DFFPOSX1 _10643_ (
    .CLK(CLK_bF$buf76),
    .D(\datapath.regrs2alu [19]),
    .Q(\datapath.memoryinterface.data_store [19])
);

DFFPOSX1 _10644_ (
    .CLK(CLK_bF$buf75),
    .D(\datapath.regrs2alu [20]),
    .Q(\datapath.memoryinterface.data_store [20])
);

DFFPOSX1 _10645_ (
    .CLK(CLK_bF$buf74),
    .D(\datapath.regrs2alu [21]),
    .Q(\datapath.memoryinterface.data_store [21])
);

DFFPOSX1 _10646_ (
    .CLK(CLK_bF$buf73),
    .D(\datapath.regrs2alu [22]),
    .Q(\datapath.memoryinterface.data_store [22])
);

DFFPOSX1 _10647_ (
    .CLK(CLK_bF$buf72),
    .D(\datapath.regrs2alu [23]),
    .Q(\datapath.memoryinterface.data_store [23])
);

DFFPOSX1 _10648_ (
    .CLK(CLK_bF$buf71),
    .D(\datapath.regrs2alu [24]),
    .Q(\datapath.memoryinterface.data_store [24])
);

DFFPOSX1 _10649_ (
    .CLK(CLK_bF$buf70),
    .D(\datapath.regrs2alu [25]),
    .Q(\datapath.memoryinterface.data_store [25])
);

DFFPOSX1 _10650_ (
    .CLK(CLK_bF$buf69),
    .D(\datapath.regrs2alu [26]),
    .Q(\datapath.memoryinterface.data_store [26])
);

DFFPOSX1 _10651_ (
    .CLK(CLK_bF$buf68),
    .D(\datapath.regrs2alu [27]),
    .Q(\datapath.memoryinterface.data_store [27])
);

DFFPOSX1 _10652_ (
    .CLK(CLK_bF$buf67),
    .D(\datapath.regrs2alu [28]),
    .Q(\datapath.memoryinterface.data_store [28])
);

DFFPOSX1 _10653_ (
    .CLK(CLK_bF$buf66),
    .D(\datapath.regrs2alu [29]),
    .Q(\datapath.memoryinterface.data_store [29])
);

DFFPOSX1 _10654_ (
    .CLK(CLK_bF$buf65),
    .D(\datapath.regrs2alu [30]),
    .Q(\datapath.memoryinterface.data_store [30])
);

DFFPOSX1 _10655_ (
    .CLK(CLK_bF$buf64),
    .D(\datapath.regrs2alu [31]),
    .Q(\datapath.memoryinterface.data_store [31])
);

DFFPOSX1 _10656_ (
    .CLK(CLK_bF$buf63),
    .D(\datapath.alu.condtrue ),
    .Q(_0_[0])
);

DFFPOSX1 _10657_ (
    .CLK(CLK_bF$buf62),
    .D(\datapath.alu.c [1]),
    .Q(_0_[1])
);

DFFPOSX1 _10658_ (
    .CLK(CLK_bF$buf61),
    .D(\datapath.alu.c [2]),
    .Q(_0_[2])
);

DFFPOSX1 _10659_ (
    .CLK(CLK_bF$buf60),
    .D(\datapath.alu.c [3]),
    .Q(_0_[3])
);

DFFPOSX1 _10660_ (
    .CLK(CLK_bF$buf59),
    .D(\datapath.alu.c [4]),
    .Q(_0_[4])
);

DFFPOSX1 _10661_ (
    .CLK(CLK_bF$buf58),
    .D(\datapath.alu.c [5]),
    .Q(_0_[5])
);

DFFPOSX1 _10662_ (
    .CLK(CLK_bF$buf57),
    .D(\datapath.alu.c [6]),
    .Q(_0_[6])
);

DFFPOSX1 _10663_ (
    .CLK(CLK_bF$buf56),
    .D(\datapath.alu.c [7]),
    .Q(_0_[7])
);

DFFPOSX1 _10664_ (
    .CLK(CLK_bF$buf55),
    .D(\datapath.alu.c [8]),
    .Q(_0_[8])
);

DFFPOSX1 _10665_ (
    .CLK(CLK_bF$buf54),
    .D(\datapath.alu.c [9]),
    .Q(_0_[9])
);

DFFPOSX1 _10666_ (
    .CLK(CLK_bF$buf53),
    .D(\datapath.alu.c [10]),
    .Q(_0_[10])
);

DFFPOSX1 _10667_ (
    .CLK(CLK_bF$buf52),
    .D(\datapath.alu.c [11]),
    .Q(_0_[11])
);

DFFPOSX1 _10668_ (
    .CLK(CLK_bF$buf51),
    .D(\datapath.alu.c [12]),
    .Q(_0_[12])
);

DFFPOSX1 _10669_ (
    .CLK(CLK_bF$buf50),
    .D(\datapath.alu.c [13]),
    .Q(_0_[13])
);

DFFPOSX1 _10670_ (
    .CLK(CLK_bF$buf49),
    .D(\datapath.alu.c [14]),
    .Q(_0_[14])
);

DFFPOSX1 _10671_ (
    .CLK(CLK_bF$buf48),
    .D(\datapath.alu.c [15]),
    .Q(_0_[15])
);

DFFPOSX1 _10672_ (
    .CLK(CLK_bF$buf47),
    .D(\datapath.alu.c [16]),
    .Q(_0_[16])
);

DFFPOSX1 _10673_ (
    .CLK(CLK_bF$buf46),
    .D(\datapath.alu.c [17]),
    .Q(_0_[17])
);

DFFPOSX1 _10674_ (
    .CLK(CLK_bF$buf45),
    .D(\datapath.alu.c [18]),
    .Q(_0_[18])
);

DFFPOSX1 _10675_ (
    .CLK(CLK_bF$buf44),
    .D(\datapath.alu.c [19]),
    .Q(_0_[19])
);

DFFPOSX1 _10676_ (
    .CLK(CLK_bF$buf43),
    .D(\datapath.alu.c [20]),
    .Q(_0_[20])
);

DFFPOSX1 _10677_ (
    .CLK(CLK_bF$buf42),
    .D(\datapath.alu.c [21]),
    .Q(_0_[21])
);

DFFPOSX1 _10678_ (
    .CLK(CLK_bF$buf41),
    .D(\datapath.alu.c [22]),
    .Q(_0_[22])
);

DFFPOSX1 _10679_ (
    .CLK(CLK_bF$buf40),
    .D(\datapath.alu.c [23]),
    .Q(_0_[23])
);

DFFPOSX1 _10680_ (
    .CLK(CLK_bF$buf39),
    .D(\datapath.alu.c [24]),
    .Q(_0_[24])
);

DFFPOSX1 _10681_ (
    .CLK(CLK_bF$buf38),
    .D(\datapath.alu.c [25]),
    .Q(_0_[25])
);

DFFPOSX1 _10682_ (
    .CLK(CLK_bF$buf37),
    .D(\datapath.alu.c [26]),
    .Q(_0_[26])
);

DFFPOSX1 _10683_ (
    .CLK(CLK_bF$buf36),
    .D(\datapath.alu.c [27]),
    .Q(_0_[27])
);

DFFPOSX1 _10684_ (
    .CLK(CLK_bF$buf35),
    .D(\datapath.alu.c [28]),
    .Q(_0_[28])
);

DFFPOSX1 _10685_ (
    .CLK(CLK_bF$buf34),
    .D(\datapath.alu.c [29]),
    .Q(_0_[29])
);

DFFPOSX1 _10686_ (
    .CLK(CLK_bF$buf33),
    .D(\datapath.alu.c [30]),
    .Q(_0_[30])
);

DFFPOSX1 _10687_ (
    .CLK(CLK_bF$buf32),
    .D(\datapath.alu.c [31]),
    .Q(_0_[31])
);

DFFPOSX1 _10688_ (
    .CLK(CLK_bF$buf31),
    .D(\datapath.jumptarget [0]),
    .Q(\datapath.programcounter.jumps [0])
);

DFFPOSX1 _10689_ (
    .CLK(CLK_bF$buf30),
    .D(\controlunit.pc_sel [0]),
    .Q(\datapath.regpcsel [0])
);

DFFPOSX1 _10690_ (
    .CLK(CLK_bF$buf29),
    .D(\controlunit.pc_sel [1]),
    .Q(\datapath.regpcsel [1])
);

DFFPOSX1 _10691_ (
    .CLK(CLK_bF$buf28),
    .D(\datapath.alu.condtrue ),
    .Q(\datapath.regcondt )
);

DFFPOSX1 _10692_ (
    .CLK(CLK_bF$buf27),
    .D(\datapath.alu.z ),
    .Q(\datapath.regz )
);

DFFPOSX1 _10693_ (
    .CLK(CLK_bF$buf26),
    .D(\datapath.aluexecptions [0]),
    .Q(\datapath.memexecptions [0])
);

DFFPOSX1 _10694_ (
    .CLK(CLK_bF$buf25),
    .D(\datapath.aluexecptions [1]),
    .Q(\datapath.memexecptions [1])
);

DFFPOSX1 _10695_ (
    .CLK(CLK_bF$buf24),
    .D(\datapath.aluexecptions [2]),
    .Q(\datapath.memexecptions [2])
);

DFFPOSX1 _10696_ (
    .CLK(CLK_bF$buf23),
    .D(\datapath.aluinstr [0]),
    .Q(\datapath.meminstr [0])
);

DFFPOSX1 _10697_ (
    .CLK(CLK_bF$buf22),
    .D(\datapath.aluinstr [1]),
    .Q(\datapath.meminstr [1])
);

DFFPOSX1 _10698_ (
    .CLK(CLK_bF$buf21),
    .D(\datapath.aluinstr [2]),
    .Q(\datapath.meminstr [2])
);

DFFPOSX1 _10699_ (
    .CLK(CLK_bF$buf20),
    .D(\datapath.aluinstr [3]),
    .Q(\datapath.meminstr [3])
);

DFFPOSX1 _10700_ (
    .CLK(CLK_bF$buf19),
    .D(\datapath.aluinstr [4]),
    .Q(\datapath.meminstr [4])
);

DFFPOSX1 _10701_ (
    .CLK(CLK_bF$buf18),
    .D(\datapath.aluinstr [5]),
    .Q(\datapath.meminstr [5])
);

DFFPOSX1 _10702_ (
    .CLK(CLK_bF$buf17),
    .D(\datapath.aluinstr [6]),
    .Q(\datapath.meminstr [6])
);

DFFPOSX1 _10703_ (
    .CLK(CLK_bF$buf16),
    .D(\datapath.aluinstr [7]),
    .Q(\datapath.meminstr [7])
);

DFFPOSX1 _10704_ (
    .CLK(CLK_bF$buf15),
    .D(\datapath.aluinstr [8]),
    .Q(\datapath.meminstr [8])
);

DFFPOSX1 _10705_ (
    .CLK(CLK_bF$buf14),
    .D(\datapath.aluinstr [9]),
    .Q(\datapath.meminstr [9])
);

DFFPOSX1 _10706_ (
    .CLK(CLK_bF$buf13),
    .D(\datapath.aluinstr [10]),
    .Q(\datapath.meminstr [10])
);

DFFPOSX1 _10707_ (
    .CLK(CLK_bF$buf12),
    .D(\datapath.aluinstr [11]),
    .Q(\datapath.meminstr [11])
);

DFFPOSX1 _10708_ (
    .CLK(CLK_bF$buf11),
    .D(\datapath.aluinstr [12]),
    .Q(\datapath.meminstr [12])
);

DFFPOSX1 _10709_ (
    .CLK(CLK_bF$buf10),
    .D(\datapath.aluinstr [13]),
    .Q(\datapath.meminstr [13])
);

DFFPOSX1 _10710_ (
    .CLK(CLK_bF$buf9),
    .D(\datapath.aluinstr [14]),
    .Q(\datapath.meminstr [14])
);

DFFPOSX1 _10711_ (
    .CLK(CLK_bF$buf8),
    .D(\datapath.aluinstr [15]),
    .Q(\datapath.meminstr [15])
);

DFFPOSX1 _10712_ (
    .CLK(CLK_bF$buf7),
    .D(\datapath.aluinstr [16]),
    .Q(\datapath.meminstr [16])
);

DFFPOSX1 _10713_ (
    .CLK(CLK_bF$buf6),
    .D(\datapath.aluinstr [17]),
    .Q(\datapath.meminstr [17])
);

DFFPOSX1 _10714_ (
    .CLK(CLK_bF$buf5),
    .D(\datapath.aluinstr [18]),
    .Q(\datapath.meminstr [18])
);

DFFPOSX1 _10715_ (
    .CLK(CLK_bF$buf4),
    .D(\datapath.aluinstr [19]),
    .Q(\datapath.meminstr [19])
);

DFFPOSX1 _10716_ (
    .CLK(CLK_bF$buf3),
    .D(\datapath.aluinstr [20]),
    .Q(\datapath.meminstr [20])
);

DFFPOSX1 _10717_ (
    .CLK(CLK_bF$buf2),
    .D(\datapath.aluinstr [21]),
    .Q(\datapath.meminstr [21])
);

DFFPOSX1 _10718_ (
    .CLK(CLK_bF$buf1),
    .D(\datapath.aluinstr [22]),
    .Q(\datapath.meminstr [22])
);

DFFPOSX1 _10719_ (
    .CLK(CLK_bF$buf0),
    .D(\datapath.aluinstr [23]),
    .Q(\datapath.meminstr [23])
);

DFFPOSX1 _10720_ (
    .CLK(CLK_bF$buf151),
    .D(\datapath.aluinstr [24]),
    .Q(\datapath.meminstr [24])
);

DFFPOSX1 _10721_ (
    .CLK(CLK_bF$buf150),
    .D(\datapath.aluinstr [25]),
    .Q(\datapath.meminstr [25])
);

DFFPOSX1 _10722_ (
    .CLK(CLK_bF$buf149),
    .D(\datapath.aluinstr [26]),
    .Q(\datapath.meminstr [26])
);

DFFPOSX1 _10723_ (
    .CLK(CLK_bF$buf148),
    .D(\datapath.aluinstr [27]),
    .Q(\datapath.meminstr [27])
);

DFFPOSX1 _10724_ (
    .CLK(CLK_bF$buf147),
    .D(\datapath.aluinstr [28]),
    .Q(\datapath.meminstr [28])
);

DFFPOSX1 _10725_ (
    .CLK(CLK_bF$buf146),
    .D(\datapath.aluinstr [29]),
    .Q(\datapath.meminstr [29])
);

DFFPOSX1 _10726_ (
    .CLK(CLK_bF$buf145),
    .D(\datapath.aluinstr [30]),
    .Q(\datapath.meminstr [30])
);

DFFPOSX1 _10727_ (
    .CLK(CLK_bF$buf144),
    .D(\datapath.aluinstr [31]),
    .Q(\datapath.meminstr [31])
);

DFFPOSX1 _10728_ (
    .CLK(CLK_bF$buf143),
    .D(\datapath.alupc_4 [0]),
    .Q(\datapath.mempc_4 [0])
);

DFFPOSX1 _10729_ (
    .CLK(CLK_bF$buf142),
    .D(\datapath.alupc_4 [1]),
    .Q(\datapath.mempc_4 [1])
);

DFFPOSX1 _10730_ (
    .CLK(CLK_bF$buf141),
    .D(\datapath.alupc_4 [2]),
    .Q(\datapath.mempc_4 [2])
);

DFFPOSX1 _10731_ (
    .CLK(CLK_bF$buf140),
    .D(\datapath.alupc_4 [3]),
    .Q(\datapath.mempc_4 [3])
);

DFFPOSX1 _10732_ (
    .CLK(CLK_bF$buf139),
    .D(\datapath.alupc_4 [4]),
    .Q(\datapath.mempc_4 [4])
);

DFFPOSX1 _10733_ (
    .CLK(CLK_bF$buf138),
    .D(\datapath.alupc_4 [5]),
    .Q(\datapath.mempc_4 [5])
);

DFFPOSX1 _10734_ (
    .CLK(CLK_bF$buf137),
    .D(\datapath.alupc_4 [6]),
    .Q(\datapath.mempc_4 [6])
);

DFFPOSX1 _10735_ (
    .CLK(CLK_bF$buf136),
    .D(\datapath.alupc_4 [7]),
    .Q(\datapath.mempc_4 [7])
);

DFFPOSX1 _10736_ (
    .CLK(CLK_bF$buf135),
    .D(\datapath.alupc_4 [8]),
    .Q(\datapath.mempc_4 [8])
);

DFFPOSX1 _10737_ (
    .CLK(CLK_bF$buf134),
    .D(\datapath.alupc_4 [9]),
    .Q(\datapath.mempc_4 [9])
);

DFFPOSX1 _10738_ (
    .CLK(CLK_bF$buf133),
    .D(\datapath.alupc_4 [10]),
    .Q(\datapath.mempc_4 [10])
);

DFFPOSX1 _10739_ (
    .CLK(CLK_bF$buf132),
    .D(\datapath.alupc_4 [11]),
    .Q(\datapath.mempc_4 [11])
);

DFFPOSX1 _10740_ (
    .CLK(CLK_bF$buf131),
    .D(\datapath.alupc_4 [12]),
    .Q(\datapath.mempc_4 [12])
);

DFFPOSX1 _10741_ (
    .CLK(CLK_bF$buf130),
    .D(\datapath.alupc_4 [13]),
    .Q(\datapath.mempc_4 [13])
);

DFFPOSX1 _10742_ (
    .CLK(CLK_bF$buf129),
    .D(\datapath.alupc_4 [14]),
    .Q(\datapath.mempc_4 [14])
);

DFFPOSX1 _10743_ (
    .CLK(CLK_bF$buf128),
    .D(\datapath.alupc_4 [15]),
    .Q(\datapath.mempc_4 [15])
);

DFFPOSX1 _10744_ (
    .CLK(CLK_bF$buf127),
    .D(\datapath.alupc_4 [16]),
    .Q(\datapath.mempc_4 [16])
);

DFFPOSX1 _10745_ (
    .CLK(CLK_bF$buf126),
    .D(\datapath.alupc_4 [17]),
    .Q(\datapath.mempc_4 [17])
);

DFFPOSX1 _10746_ (
    .CLK(CLK_bF$buf125),
    .D(\datapath.alupc_4 [18]),
    .Q(\datapath.mempc_4 [18])
);

DFFPOSX1 _10747_ (
    .CLK(CLK_bF$buf124),
    .D(\datapath.alupc_4 [19]),
    .Q(\datapath.mempc_4 [19])
);

DFFPOSX1 _10748_ (
    .CLK(CLK_bF$buf123),
    .D(\datapath.alupc_4 [20]),
    .Q(\datapath.mempc_4 [20])
);

DFFPOSX1 _10749_ (
    .CLK(CLK_bF$buf122),
    .D(\datapath.alupc_4 [21]),
    .Q(\datapath.mempc_4 [21])
);

DFFPOSX1 _10750_ (
    .CLK(CLK_bF$buf121),
    .D(\datapath.alupc_4 [22]),
    .Q(\datapath.mempc_4 [22])
);

DFFPOSX1 _10751_ (
    .CLK(CLK_bF$buf120),
    .D(\datapath.alupc_4 [23]),
    .Q(\datapath.mempc_4 [23])
);

DFFPOSX1 _10752_ (
    .CLK(CLK_bF$buf119),
    .D(\datapath.alupc_4 [24]),
    .Q(\datapath.mempc_4 [24])
);

DFFPOSX1 _10753_ (
    .CLK(CLK_bF$buf118),
    .D(\datapath.alupc_4 [25]),
    .Q(\datapath.mempc_4 [25])
);

DFFPOSX1 _10754_ (
    .CLK(CLK_bF$buf117),
    .D(\datapath.alupc_4 [26]),
    .Q(\datapath.mempc_4 [26])
);

DFFPOSX1 _10755_ (
    .CLK(CLK_bF$buf116),
    .D(\datapath.alupc_4 [27]),
    .Q(\datapath.mempc_4 [27])
);

DFFPOSX1 _10756_ (
    .CLK(CLK_bF$buf115),
    .D(\datapath.alupc_4 [28]),
    .Q(\datapath.mempc_4 [28])
);

DFFPOSX1 _10757_ (
    .CLK(CLK_bF$buf114),
    .D(\datapath.alupc_4 [29]),
    .Q(\datapath.mempc_4 [29])
);

DFFPOSX1 _10758_ (
    .CLK(CLK_bF$buf113),
    .D(\datapath.alupc_4 [30]),
    .Q(\datapath.mempc_4 [30])
);

DFFPOSX1 _10759_ (
    .CLK(CLK_bF$buf112),
    .D(\datapath.alupc_4 [31]),
    .Q(\datapath.mempc_4 [31])
);

DFFPOSX1 _10760_ (
    .CLK(CLK_bF$buf111),
    .D(\datapath.alupc [2]),
    .Q(\datapath.csr.csr_mepc [2])
);

DFFPOSX1 _10761_ (
    .CLK(CLK_bF$buf110),
    .D(\datapath.alupc [3]),
    .Q(\datapath.csr.csr_mepc [3])
);

DFFPOSX1 _10762_ (
    .CLK(CLK_bF$buf109),
    .D(\datapath.alupc [4]),
    .Q(\datapath.csr.csr_mepc [4])
);

DFFPOSX1 _10763_ (
    .CLK(CLK_bF$buf108),
    .D(\datapath.alupc [5]),
    .Q(\datapath.csr.csr_mepc [5])
);

DFFPOSX1 _10764_ (
    .CLK(CLK_bF$buf107),
    .D(\datapath.alupc [6]),
    .Q(\datapath.csr.csr_mepc [6])
);

DFFPOSX1 _10765_ (
    .CLK(CLK_bF$buf106),
    .D(\datapath.alupc [7]),
    .Q(\datapath.csr.csr_mepc [7])
);

DFFPOSX1 _10766_ (
    .CLK(CLK_bF$buf105),
    .D(\datapath.alupc [8]),
    .Q(\datapath.csr.csr_mepc [8])
);

DFFPOSX1 _10767_ (
    .CLK(CLK_bF$buf104),
    .D(\datapath.alupc [9]),
    .Q(\datapath.csr.csr_mepc [9])
);

DFFPOSX1 _10768_ (
    .CLK(CLK_bF$buf103),
    .D(\datapath.alupc [10]),
    .Q(\datapath.csr.csr_mepc [10])
);

DFFPOSX1 _10769_ (
    .CLK(CLK_bF$buf102),
    .D(\datapath.alupc [11]),
    .Q(\datapath.csr.csr_mepc [11])
);

DFFPOSX1 _10770_ (
    .CLK(CLK_bF$buf101),
    .D(\datapath.alupc [12]),
    .Q(\datapath.csr.csr_mepc [12])
);

DFFPOSX1 _10771_ (
    .CLK(CLK_bF$buf100),
    .D(\datapath.alupc [13]),
    .Q(\datapath.csr.csr_mepc [13])
);

DFFPOSX1 _10772_ (
    .CLK(CLK_bF$buf99),
    .D(\datapath.alupc [14]),
    .Q(\datapath.csr.csr_mepc [14])
);

DFFPOSX1 _10773_ (
    .CLK(CLK_bF$buf98),
    .D(\datapath.alupc [15]),
    .Q(\datapath.csr.csr_mepc [15])
);

DFFPOSX1 _10774_ (
    .CLK(CLK_bF$buf97),
    .D(\datapath.alupc [16]),
    .Q(\datapath.csr.csr_mepc [16])
);

DFFPOSX1 _10775_ (
    .CLK(CLK_bF$buf96),
    .D(\datapath.alupc [17]),
    .Q(\datapath.csr.csr_mepc [17])
);

DFFPOSX1 _10776_ (
    .CLK(CLK_bF$buf95),
    .D(\datapath.alupc [18]),
    .Q(\datapath.csr.csr_mepc [18])
);

DFFPOSX1 _10777_ (
    .CLK(CLK_bF$buf94),
    .D(\datapath.alupc [19]),
    .Q(\datapath.csr.csr_mepc [19])
);

DFFPOSX1 _10778_ (
    .CLK(CLK_bF$buf93),
    .D(\datapath.alupc [20]),
    .Q(\datapath.csr.csr_mepc [20])
);

DFFPOSX1 _10779_ (
    .CLK(CLK_bF$buf92),
    .D(\datapath.alupc [21]),
    .Q(\datapath.csr.csr_mepc [21])
);

DFFPOSX1 _10780_ (
    .CLK(CLK_bF$buf91),
    .D(\datapath.alupc [22]),
    .Q(\datapath.csr.csr_mepc [22])
);

DFFPOSX1 _10781_ (
    .CLK(CLK_bF$buf90),
    .D(\datapath.alupc [23]),
    .Q(\datapath.csr.csr_mepc [23])
);

DFFPOSX1 _10782_ (
    .CLK(CLK_bF$buf89),
    .D(\datapath.alupc [24]),
    .Q(\datapath.csr.csr_mepc [24])
);

DFFPOSX1 _10783_ (
    .CLK(CLK_bF$buf88),
    .D(\datapath.alupc [25]),
    .Q(\datapath.csr.csr_mepc [25])
);

DFFPOSX1 _10784_ (
    .CLK(CLK_bF$buf87),
    .D(\datapath.alupc [26]),
    .Q(\datapath.csr.csr_mepc [26])
);

DFFPOSX1 _10785_ (
    .CLK(CLK_bF$buf86),
    .D(\datapath.alupc [27]),
    .Q(\datapath.csr.csr_mepc [27])
);

DFFPOSX1 _10786_ (
    .CLK(CLK_bF$buf85),
    .D(\datapath.alupc [28]),
    .Q(\datapath.csr.csr_mepc [28])
);

DFFPOSX1 _10787_ (
    .CLK(CLK_bF$buf84),
    .D(\datapath.alupc [29]),
    .Q(\datapath.csr.csr_mepc [29])
);

DFFPOSX1 _10788_ (
    .CLK(CLK_bF$buf83),
    .D(\datapath.alupc [30]),
    .Q(\datapath.csr.csr_mepc [30])
);

DFFPOSX1 _10789_ (
    .CLK(CLK_bF$buf82),
    .D(\datapath.alupc [31]),
    .Q(\datapath.csr.csr_mepc [31])
);

DFFPOSX1 _10790_ (
    .CLK(CLK_bF$buf81),
    .D(\datapath.immediatedecoder._06_ ),
    .Q(\datapath.regimmalu [0])
);

DFFPOSX1 _10791_ (
    .CLK(CLK_bF$buf80),
    .D(\datapath.imm [1]),
    .Q(\datapath.regimmalu [1])
);

DFFPOSX1 _10792_ (
    .CLK(CLK_bF$buf79),
    .D(\datapath.imm [2]),
    .Q(\datapath.regimmalu [2])
);

DFFPOSX1 _10793_ (
    .CLK(CLK_bF$buf78),
    .D(\datapath.imm [3]),
    .Q(\datapath.regimmalu [3])
);

DFFPOSX1 _10794_ (
    .CLK(CLK_bF$buf77),
    .D(\datapath.imm [4]),
    .Q(\datapath.regimmalu [4])
);

DFFPOSX1 _10795_ (
    .CLK(CLK_bF$buf76),
    .D(\datapath.imm [5]),
    .Q(\datapath.regimmalu [5])
);

DFFPOSX1 _10796_ (
    .CLK(CLK_bF$buf75),
    .D(\datapath.imm [6]),
    .Q(\datapath.regimmalu [6])
);

DFFPOSX1 _10797_ (
    .CLK(CLK_bF$buf74),
    .D(\datapath.imm [7]),
    .Q(\datapath.regimmalu [7])
);

DFFPOSX1 _10798_ (
    .CLK(CLK_bF$buf73),
    .D(\datapath.imm [8]),
    .Q(\datapath.regimmalu [8])
);

DFFPOSX1 _10799_ (
    .CLK(CLK_bF$buf72),
    .D(\datapath.imm [9]),
    .Q(\datapath.regimmalu [9])
);

DFFPOSX1 _10800_ (
    .CLK(CLK_bF$buf71),
    .D(\datapath.imm [10]),
    .Q(\datapath.regimmalu [10])
);

DFFPOSX1 _10801_ (
    .CLK(CLK_bF$buf70),
    .D(\datapath.immediatedecoder._09_ ),
    .Q(\datapath.regimmalu [11])
);

DFFPOSX1 _10802_ (
    .CLK(CLK_bF$buf69),
    .D(\datapath.imm [12]),
    .Q(\datapath.regimmalu [12])
);

DFFPOSX1 _10803_ (
    .CLK(CLK_bF$buf68),
    .D(\datapath.imm [13]),
    .Q(\datapath.regimmalu [13])
);

DFFPOSX1 _10804_ (
    .CLK(CLK_bF$buf67),
    .D(\datapath.imm [14]),
    .Q(\datapath.regimmalu [14])
);

DFFPOSX1 _10805_ (
    .CLK(CLK_bF$buf66),
    .D(\datapath.imm [15]),
    .Q(\datapath.regimmalu [15])
);

DFFPOSX1 _10806_ (
    .CLK(CLK_bF$buf65),
    .D(\datapath.imm [16]),
    .Q(\datapath.regimmalu [16])
);

DFFPOSX1 _10807_ (
    .CLK(CLK_bF$buf64),
    .D(\datapath.imm [17]),
    .Q(\datapath.regimmalu [17])
);

DFFPOSX1 _10808_ (
    .CLK(CLK_bF$buf63),
    .D(\datapath.imm [18]),
    .Q(\datapath.regimmalu [18])
);

DFFPOSX1 _10809_ (
    .CLK(CLK_bF$buf62),
    .D(\datapath.imm [19]),
    .Q(\datapath.regimmalu [19])
);

DFFPOSX1 _10810_ (
    .CLK(CLK_bF$buf61),
    .D(\datapath.imm [20]),
    .Q(\datapath.regimmalu [20])
);

DFFPOSX1 _10811_ (
    .CLK(CLK_bF$buf60),
    .D(\datapath.imm [21]),
    .Q(\datapath.regimmalu [21])
);

DFFPOSX1 _10812_ (
    .CLK(CLK_bF$buf59),
    .D(\datapath.imm [22]),
    .Q(\datapath.regimmalu [22])
);

DFFPOSX1 _10813_ (
    .CLK(CLK_bF$buf58),
    .D(\datapath.imm [23]),
    .Q(\datapath.regimmalu [23])
);

DFFPOSX1 _10814_ (
    .CLK(CLK_bF$buf57),
    .D(\datapath.imm [24]),
    .Q(\datapath.regimmalu [24])
);

DFFPOSX1 _10815_ (
    .CLK(CLK_bF$buf56),
    .D(\datapath.imm [25]),
    .Q(\datapath.regimmalu [25])
);

DFFPOSX1 _10816_ (
    .CLK(CLK_bF$buf55),
    .D(\datapath.imm [26]),
    .Q(\datapath.regimmalu [26])
);

DFFPOSX1 _10817_ (
    .CLK(CLK_bF$buf54),
    .D(\datapath.imm [27]),
    .Q(\datapath.regimmalu [27])
);

DFFPOSX1 _10818_ (
    .CLK(CLK_bF$buf53),
    .D(\datapath.imm [28]),
    .Q(\datapath.regimmalu [28])
);

DFFPOSX1 _10819_ (
    .CLK(CLK_bF$buf52),
    .D(\datapath.imm [29]),
    .Q(\datapath.regimmalu [29])
);

DFFPOSX1 _10820_ (
    .CLK(CLK_bF$buf51),
    .D(\datapath.imm [30]),
    .Q(\datapath.regimmalu [30])
);

DFFPOSX1 _10821_ (
    .CLK(CLK_bF$buf50),
    .D(\datapath.immediatedecoder._12_ ),
    .Q(\datapath.regimmalu [31])
);

DFFPOSX1 _10822_ (
    .CLK(CLK_bF$buf49),
    .D(\datapath.csr.csr_data [0]),
    .Q(\datapath.regcsralu [0])
);

DFFPOSX1 _10823_ (
    .CLK(CLK_bF$buf48),
    .D(\datapath.csr.csr_data [1]),
    .Q(\datapath.regcsralu [1])
);

DFFPOSX1 _10824_ (
    .CLK(CLK_bF$buf47),
    .D(\datapath.csr.csr_data [2]),
    .Q(\datapath.regcsralu [2])
);

DFFPOSX1 _10825_ (
    .CLK(CLK_bF$buf46),
    .D(\datapath.csr.csr_data [3]),
    .Q(\datapath.regcsralu [3])
);

DFFPOSX1 _10826_ (
    .CLK(CLK_bF$buf45),
    .D(\datapath.csr.csr_data [4]),
    .Q(\datapath.regcsralu [4])
);

DFFPOSX1 _10827_ (
    .CLK(CLK_bF$buf44),
    .D(\datapath.csr.csr_data [5]),
    .Q(\datapath.regcsralu [5])
);

DFFPOSX1 _10828_ (
    .CLK(CLK_bF$buf43),
    .D(\datapath.csr.csr_data [6]),
    .Q(\datapath.regcsralu [6])
);

DFFPOSX1 _10829_ (
    .CLK(CLK_bF$buf42),
    .D(\datapath.csr.csr_data [7]),
    .Q(\datapath.regcsralu [7])
);

DFFPOSX1 _10830_ (
    .CLK(CLK_bF$buf41),
    .D(\datapath.csr.csr_data [8]),
    .Q(\datapath.regcsralu [8])
);

DFFPOSX1 _10831_ (
    .CLK(CLK_bF$buf40),
    .D(\datapath.csr.csr_data [9]),
    .Q(\datapath.regcsralu [9])
);

DFFPOSX1 _10832_ (
    .CLK(CLK_bF$buf39),
    .D(\datapath.csr.csr_data [10]),
    .Q(\datapath.regcsralu [10])
);

DFFPOSX1 _10833_ (
    .CLK(CLK_bF$buf38),
    .D(\datapath.csr.csr_data [11]),
    .Q(\datapath.regcsralu [11])
);

DFFPOSX1 _10834_ (
    .CLK(CLK_bF$buf37),
    .D(\datapath.csr.csr_data [12]),
    .Q(\datapath.regcsralu [12])
);

DFFPOSX1 _10835_ (
    .CLK(CLK_bF$buf36),
    .D(\datapath.csr.csr_data [13]),
    .Q(\datapath.regcsralu [13])
);

DFFPOSX1 _10836_ (
    .CLK(CLK_bF$buf35),
    .D(\datapath.csr.csr_data [14]),
    .Q(\datapath.regcsralu [14])
);

DFFPOSX1 _10837_ (
    .CLK(CLK_bF$buf34),
    .D(\datapath.csr.csr_data [15]),
    .Q(\datapath.regcsralu [15])
);

DFFPOSX1 _10838_ (
    .CLK(CLK_bF$buf33),
    .D(\datapath.csr.csr_data [16]),
    .Q(\datapath.regcsralu [16])
);

DFFPOSX1 _10839_ (
    .CLK(CLK_bF$buf32),
    .D(\datapath.csr.csr_data [17]),
    .Q(\datapath.regcsralu [17])
);

DFFPOSX1 _10840_ (
    .CLK(CLK_bF$buf31),
    .D(\datapath.csr.csr_data [18]),
    .Q(\datapath.regcsralu [18])
);

DFFPOSX1 _10841_ (
    .CLK(CLK_bF$buf30),
    .D(\datapath.csr.csr_data [19]),
    .Q(\datapath.regcsralu [19])
);

DFFPOSX1 _10842_ (
    .CLK(CLK_bF$buf29),
    .D(\datapath.csr.csr_data [20]),
    .Q(\datapath.regcsralu [20])
);

DFFPOSX1 _10843_ (
    .CLK(CLK_bF$buf28),
    .D(\datapath.csr.csr_data [21]),
    .Q(\datapath.regcsralu [21])
);

DFFPOSX1 _10844_ (
    .CLK(CLK_bF$buf27),
    .D(\datapath.csr.csr_data [22]),
    .Q(\datapath.regcsralu [22])
);

DFFPOSX1 _10845_ (
    .CLK(CLK_bF$buf26),
    .D(\datapath.csr.csr_data [23]),
    .Q(\datapath.regcsralu [23])
);

DFFPOSX1 _10846_ (
    .CLK(CLK_bF$buf25),
    .D(\datapath.csr.csr_data [24]),
    .Q(\datapath.regcsralu [24])
);

DFFPOSX1 _10847_ (
    .CLK(CLK_bF$buf24),
    .D(\datapath.csr.csr_data [25]),
    .Q(\datapath.regcsralu [25])
);

DFFPOSX1 _10848_ (
    .CLK(CLK_bF$buf23),
    .D(\datapath.csr.csr_data [26]),
    .Q(\datapath.regcsralu [26])
);

DFFPOSX1 _10849_ (
    .CLK(CLK_bF$buf22),
    .D(\datapath.csr.csr_data [27]),
    .Q(\datapath.regcsralu [27])
);

DFFPOSX1 _10850_ (
    .CLK(CLK_bF$buf21),
    .D(\datapath.csr.csr_data [28]),
    .Q(\datapath.regcsralu [28])
);

DFFPOSX1 _10851_ (
    .CLK(CLK_bF$buf20),
    .D(\datapath.csr.csr_data [29]),
    .Q(\datapath.regcsralu [29])
);

DFFPOSX1 _10852_ (
    .CLK(CLK_bF$buf19),
    .D(\datapath.csr.csr_data [30]),
    .Q(\datapath.regcsralu [30])
);

DFFPOSX1 _10853_ (
    .CLK(CLK_bF$buf18),
    .D(\datapath.csr.csr_data [31]),
    .Q(\datapath.regcsralu [31])
);

DFFPOSX1 _10854_ (
    .CLK(CLK_bF$buf17),
    .D(\datapath.registers.regb_data [0]),
    .Q(\datapath.regrs2alu [0])
);

DFFPOSX1 _10855_ (
    .CLK(CLK_bF$buf16),
    .D(\datapath.registers.regb_data [1]),
    .Q(\datapath.regrs2alu [1])
);

DFFPOSX1 _10856_ (
    .CLK(CLK_bF$buf15),
    .D(\datapath.registers.regb_data [2]),
    .Q(\datapath.regrs2alu [2])
);

DFFPOSX1 _10857_ (
    .CLK(CLK_bF$buf14),
    .D(\datapath.registers.regb_data [3]),
    .Q(\datapath.regrs2alu [3])
);

DFFPOSX1 _10858_ (
    .CLK(CLK_bF$buf13),
    .D(\datapath.registers.regb_data [4]),
    .Q(\datapath.regrs2alu [4])
);

DFFPOSX1 _10859_ (
    .CLK(CLK_bF$buf12),
    .D(\datapath.registers.regb_data [5]),
    .Q(\datapath.regrs2alu [5])
);

DFFPOSX1 _10860_ (
    .CLK(CLK_bF$buf11),
    .D(\datapath.registers.regb_data [6]),
    .Q(\datapath.regrs2alu [6])
);

DFFPOSX1 _10861_ (
    .CLK(CLK_bF$buf10),
    .D(\datapath.registers.regb_data [7]),
    .Q(\datapath.regrs2alu [7])
);

DFFPOSX1 _10862_ (
    .CLK(CLK_bF$buf9),
    .D(\datapath.registers.regb_data [8]),
    .Q(\datapath.regrs2alu [8])
);

DFFPOSX1 _10863_ (
    .CLK(CLK_bF$buf8),
    .D(\datapath.registers.regb_data [9]),
    .Q(\datapath.regrs2alu [9])
);

DFFPOSX1 _10864_ (
    .CLK(CLK_bF$buf7),
    .D(\datapath.registers.regb_data [10]),
    .Q(\datapath.regrs2alu [10])
);

DFFPOSX1 _10865_ (
    .CLK(CLK_bF$buf6),
    .D(\datapath.registers.regb_data [11]),
    .Q(\datapath.regrs2alu [11])
);

DFFPOSX1 _10866_ (
    .CLK(CLK_bF$buf5),
    .D(\datapath.registers.regb_data [12]),
    .Q(\datapath.regrs2alu [12])
);

DFFPOSX1 _10867_ (
    .CLK(CLK_bF$buf4),
    .D(\datapath.registers.regb_data [13]),
    .Q(\datapath.regrs2alu [13])
);

DFFPOSX1 _10868_ (
    .CLK(CLK_bF$buf3),
    .D(\datapath.registers.regb_data [14]),
    .Q(\datapath.regrs2alu [14])
);

DFFPOSX1 _10869_ (
    .CLK(CLK_bF$buf2),
    .D(\datapath.registers.regb_data [15]),
    .Q(\datapath.regrs2alu [15])
);

DFFPOSX1 _10870_ (
    .CLK(CLK_bF$buf1),
    .D(\datapath.registers.regb_data [16]),
    .Q(\datapath.regrs2alu [16])
);

DFFPOSX1 _10871_ (
    .CLK(CLK_bF$buf0),
    .D(\datapath.registers.regb_data [17]),
    .Q(\datapath.regrs2alu [17])
);

DFFPOSX1 _10872_ (
    .CLK(CLK_bF$buf151),
    .D(\datapath.registers.regb_data [18]),
    .Q(\datapath.regrs2alu [18])
);

DFFPOSX1 _10873_ (
    .CLK(CLK_bF$buf150),
    .D(\datapath.registers.regb_data [19]),
    .Q(\datapath.regrs2alu [19])
);

DFFPOSX1 _10874_ (
    .CLK(CLK_bF$buf149),
    .D(\datapath.registers.regb_data [20]),
    .Q(\datapath.regrs2alu [20])
);

DFFPOSX1 _10875_ (
    .CLK(CLK_bF$buf148),
    .D(\datapath.registers.regb_data [21]),
    .Q(\datapath.regrs2alu [21])
);

DFFPOSX1 _10876_ (
    .CLK(CLK_bF$buf147),
    .D(\datapath.registers.regb_data [22]),
    .Q(\datapath.regrs2alu [22])
);

DFFPOSX1 _10877_ (
    .CLK(CLK_bF$buf146),
    .D(\datapath.registers.regb_data [23]),
    .Q(\datapath.regrs2alu [23])
);

DFFPOSX1 _10878_ (
    .CLK(CLK_bF$buf145),
    .D(\datapath.registers.regb_data [24]),
    .Q(\datapath.regrs2alu [24])
);

DFFPOSX1 _10879_ (
    .CLK(CLK_bF$buf144),
    .D(\datapath.registers.regb_data [25]),
    .Q(\datapath.regrs2alu [25])
);

DFFPOSX1 _10880_ (
    .CLK(CLK_bF$buf143),
    .D(\datapath.registers.regb_data [26]),
    .Q(\datapath.regrs2alu [26])
);

DFFPOSX1 _10881_ (
    .CLK(CLK_bF$buf142),
    .D(\datapath.registers.regb_data [27]),
    .Q(\datapath.regrs2alu [27])
);

DFFPOSX1 _10882_ (
    .CLK(CLK_bF$buf141),
    .D(\datapath.registers.regb_data [28]),
    .Q(\datapath.regrs2alu [28])
);

DFFPOSX1 _10883_ (
    .CLK(CLK_bF$buf140),
    .D(\datapath.registers.regb_data [29]),
    .Q(\datapath.regrs2alu [29])
);

DFFPOSX1 _10884_ (
    .CLK(CLK_bF$buf139),
    .D(\datapath.registers.regb_data [30]),
    .Q(\datapath.regrs2alu [30])
);

DFFPOSX1 _10885_ (
    .CLK(CLK_bF$buf138),
    .D(\datapath.registers.regb_data [31]),
    .Q(\datapath.regrs2alu [31])
);

DFFPOSX1 _10886_ (
    .CLK(CLK_bF$buf137),
    .D(\datapath.muxbval [0]),
    .Q(\datapath.alu.b [0])
);

DFFPOSX1 _10887_ (
    .CLK(CLK_bF$buf136),
    .D(\datapath.muxbval [1]),
    .Q(\datapath.alu.b [1])
);

DFFPOSX1 _10888_ (
    .CLK(CLK_bF$buf135),
    .D(\datapath.muxbval [2]),
    .Q(\datapath.alu.b [2])
);

DFFPOSX1 _10889_ (
    .CLK(CLK_bF$buf134),
    .D(\datapath.muxbval [3]),
    .Q(\datapath.alu.b [3])
);

DFFPOSX1 _10890_ (
    .CLK(CLK_bF$buf133),
    .D(\datapath.muxbval [4]),
    .Q(\datapath.alu.b [4])
);

DFFPOSX1 _10891_ (
    .CLK(CLK_bF$buf132),
    .D(\datapath.muxbval [5]),
    .Q(\datapath.alu.b [5])
);

DFFPOSX1 _10892_ (
    .CLK(CLK_bF$buf131),
    .D(\datapath.muxbval [6]),
    .Q(\datapath.alu.b [6])
);

DFFPOSX1 _10893_ (
    .CLK(CLK_bF$buf130),
    .D(\datapath.muxbval [7]),
    .Q(\datapath.alu.b [7])
);

DFFPOSX1 _10894_ (
    .CLK(CLK_bF$buf129),
    .D(\datapath.muxbval [8]),
    .Q(\datapath.alu.b [8])
);

DFFPOSX1 _10895_ (
    .CLK(CLK_bF$buf128),
    .D(\datapath.muxbval [9]),
    .Q(\datapath.alu.b [9])
);

DFFPOSX1 _10896_ (
    .CLK(CLK_bF$buf127),
    .D(\datapath.muxbval [10]),
    .Q(\datapath.alu.b [10])
);

DFFPOSX1 _10897_ (
    .CLK(CLK_bF$buf126),
    .D(\datapath.muxbval [11]),
    .Q(\datapath.alu.b [11])
);

DFFPOSX1 _10898_ (
    .CLK(CLK_bF$buf125),
    .D(\datapath.muxbval [12]),
    .Q(\datapath.alu.b [12])
);

DFFPOSX1 _10899_ (
    .CLK(CLK_bF$buf124),
    .D(\datapath.muxbval [13]),
    .Q(\datapath.alu.b [13])
);

DFFPOSX1 _10900_ (
    .CLK(CLK_bF$buf123),
    .D(\datapath.muxbval [14]),
    .Q(\datapath.alu.b [14])
);

DFFPOSX1 _10901_ (
    .CLK(CLK_bF$buf122),
    .D(\datapath.muxbval [15]),
    .Q(\datapath.alu.b [15])
);

DFFPOSX1 _10902_ (
    .CLK(CLK_bF$buf121),
    .D(\datapath.muxbval [16]),
    .Q(\datapath.alu.b [16])
);

DFFPOSX1 _10903_ (
    .CLK(CLK_bF$buf120),
    .D(\datapath.muxbval [17]),
    .Q(\datapath.alu.b [17])
);

DFFPOSX1 _10904_ (
    .CLK(CLK_bF$buf119),
    .D(\datapath.muxbval [18]),
    .Q(\datapath.alu.b [18])
);

DFFPOSX1 _10905_ (
    .CLK(CLK_bF$buf118),
    .D(\datapath.muxbval [19]),
    .Q(\datapath.alu.b [19])
);

DFFPOSX1 _10906_ (
    .CLK(CLK_bF$buf117),
    .D(\datapath.muxbval [20]),
    .Q(\datapath.alu.b [20])
);

DFFPOSX1 _10907_ (
    .CLK(CLK_bF$buf116),
    .D(\datapath.muxbval [21]),
    .Q(\datapath.alu.b [21])
);

DFFPOSX1 _10908_ (
    .CLK(CLK_bF$buf115),
    .D(\datapath.muxbval [22]),
    .Q(\datapath.alu.b [22])
);

DFFPOSX1 _10909_ (
    .CLK(CLK_bF$buf114),
    .D(\datapath.muxbval [23]),
    .Q(\datapath.alu.b [23])
);

DFFPOSX1 _10910_ (
    .CLK(CLK_bF$buf113),
    .D(\datapath.muxbval [24]),
    .Q(\datapath.alu.b [24])
);

DFFPOSX1 _10911_ (
    .CLK(CLK_bF$buf112),
    .D(\datapath.muxbval [25]),
    .Q(\datapath.alu.b [25])
);

DFFPOSX1 _10912_ (
    .CLK(CLK_bF$buf111),
    .D(\datapath.muxbval [26]),
    .Q(\datapath.alu.b [26])
);

DFFPOSX1 _10913_ (
    .CLK(CLK_bF$buf110),
    .D(\datapath.muxbval [27]),
    .Q(\datapath.alu.b [27])
);

DFFPOSX1 _10914_ (
    .CLK(CLK_bF$buf109),
    .D(\datapath.muxbval [28]),
    .Q(\datapath.alu.b [28])
);

DFFPOSX1 _10915_ (
    .CLK(CLK_bF$buf108),
    .D(\datapath.muxbval [29]),
    .Q(\datapath.alu.b [29])
);

DFFPOSX1 _10916_ (
    .CLK(CLK_bF$buf107),
    .D(\datapath.muxbval [30]),
    .Q(\datapath.alu.b [30])
);

DFFPOSX1 _10917_ (
    .CLK(CLK_bF$buf106),
    .D(\datapath.muxbval [31]),
    .Q(\datapath.alu.b [31])
);

DFFPOSX1 _10918_ (
    .CLK(CLK_bF$buf105),
    .D(\datapath.muxaval [0]),
    .Q(\datapath.alu.a [0])
);

DFFPOSX1 _10919_ (
    .CLK(CLK_bF$buf104),
    .D(\datapath.muxaval [1]),
    .Q(\datapath.alu.a [1])
);

DFFPOSX1 _10920_ (
    .CLK(CLK_bF$buf103),
    .D(\datapath.muxaval [2]),
    .Q(\datapath.alu.a [2])
);

DFFPOSX1 _10921_ (
    .CLK(CLK_bF$buf102),
    .D(\datapath.muxaval [3]),
    .Q(\datapath.alu.a [3])
);

DFFPOSX1 _10922_ (
    .CLK(CLK_bF$buf101),
    .D(\datapath.muxaval [4]),
    .Q(\datapath.alu.a [4])
);

DFFPOSX1 _10923_ (
    .CLK(CLK_bF$buf100),
    .D(\datapath.muxaval [5]),
    .Q(\datapath.alu.a [5])
);

DFFPOSX1 _10924_ (
    .CLK(CLK_bF$buf99),
    .D(\datapath.muxaval [6]),
    .Q(\datapath.alu.a [6])
);

DFFPOSX1 _10925_ (
    .CLK(CLK_bF$buf98),
    .D(\datapath.muxaval [7]),
    .Q(\datapath.alu.a [7])
);

DFFPOSX1 _10926_ (
    .CLK(CLK_bF$buf97),
    .D(\datapath.muxaval [8]),
    .Q(\datapath.alu.a [8])
);

DFFPOSX1 _10927_ (
    .CLK(CLK_bF$buf96),
    .D(\datapath.muxaval [9]),
    .Q(\datapath.alu.a [9])
);

DFFPOSX1 _10928_ (
    .CLK(CLK_bF$buf95),
    .D(\datapath.muxaval [10]),
    .Q(\datapath.alu.a [10])
);

DFFPOSX1 _10929_ (
    .CLK(CLK_bF$buf94),
    .D(\datapath.muxaval [11]),
    .Q(\datapath.alu.a [11])
);

DFFPOSX1 _10930_ (
    .CLK(CLK_bF$buf93),
    .D(\datapath.muxaval [12]),
    .Q(\datapath.alu.a [12])
);

DFFPOSX1 _10931_ (
    .CLK(CLK_bF$buf92),
    .D(\datapath.muxaval [13]),
    .Q(\datapath.alu.a [13])
);

DFFPOSX1 _10932_ (
    .CLK(CLK_bF$buf91),
    .D(\datapath.muxaval [14]),
    .Q(\datapath.alu.a [14])
);

DFFPOSX1 _10933_ (
    .CLK(CLK_bF$buf90),
    .D(\datapath.muxaval [15]),
    .Q(\datapath.alu.a [15])
);

DFFPOSX1 _10934_ (
    .CLK(CLK_bF$buf89),
    .D(\datapath.muxaval [16]),
    .Q(\datapath.alu.a [16])
);

DFFPOSX1 _10935_ (
    .CLK(CLK_bF$buf88),
    .D(\datapath.muxaval [17]),
    .Q(\datapath.alu.a [17])
);

DFFPOSX1 _10936_ (
    .CLK(CLK_bF$buf87),
    .D(\datapath.muxaval [18]),
    .Q(\datapath.alu.a [18])
);

DFFPOSX1 _10937_ (
    .CLK(CLK_bF$buf86),
    .D(\datapath.muxaval [19]),
    .Q(\datapath.alu.a [19])
);

DFFPOSX1 _10938_ (
    .CLK(CLK_bF$buf85),
    .D(\datapath.muxaval [20]),
    .Q(\datapath.alu.a [20])
);

DFFPOSX1 _10939_ (
    .CLK(CLK_bF$buf84),
    .D(\datapath.muxaval [21]),
    .Q(\datapath.alu.a [21])
);

DFFPOSX1 _10940_ (
    .CLK(CLK_bF$buf83),
    .D(\datapath.muxaval [22]),
    .Q(\datapath.alu.a [22])
);

DFFPOSX1 _10941_ (
    .CLK(CLK_bF$buf82),
    .D(\datapath.muxaval [23]),
    .Q(\datapath.alu.a [23])
);

DFFPOSX1 _10942_ (
    .CLK(CLK_bF$buf81),
    .D(\datapath.muxaval [24]),
    .Q(\datapath.alu.a [24])
);

DFFPOSX1 _10943_ (
    .CLK(CLK_bF$buf80),
    .D(\datapath.muxaval [25]),
    .Q(\datapath.alu.a [25])
);

DFFPOSX1 _10944_ (
    .CLK(CLK_bF$buf79),
    .D(\datapath.muxaval [26]),
    .Q(\datapath.alu.a [26])
);

DFFPOSX1 _10945_ (
    .CLK(CLK_bF$buf78),
    .D(\datapath.muxaval [27]),
    .Q(\datapath.alu.a [27])
);

DFFPOSX1 _10946_ (
    .CLK(CLK_bF$buf77),
    .D(\datapath.muxaval [28]),
    .Q(\datapath.alu.a [28])
);

DFFPOSX1 _10947_ (
    .CLK(CLK_bF$buf76),
    .D(\datapath.muxaval [29]),
    .Q(\datapath.alu.a [29])
);

DFFPOSX1 _10948_ (
    .CLK(CLK_bF$buf75),
    .D(\datapath.muxaval [30]),
    .Q(\datapath.alu.a [30])
);

DFFPOSX1 _10949_ (
    .CLK(CLK_bF$buf74),
    .D(\datapath.muxaval [31]),
    .Q(\datapath.alu.a [31])
);

DFFPOSX1 _10950_ (
    .CLK(CLK_bF$buf73),
    .D(alusel[0]),
    .Q(\datapath.alu.funsel [0])
);

DFFPOSX1 _10951_ (
    .CLK(CLK_bF$buf72),
    .D(alusel[1]),
    .Q(\datapath.alu.funsel [1])
);

DFFPOSX1 _10952_ (
    .CLK(CLK_bF$buf71),
    .D(alusel[2]),
    .Q(\datapath.alu.funsel [2])
);

DFFPOSX1 _10953_ (
    .CLK(CLK_bF$buf70),
    .D(alusel[3]),
    .Q(\datapath.alu.funsel [3])
);

DFFPOSX1 _10954_ (
    .CLK(CLK_bF$buf69),
    .D(\controlunit.ill_op ),
    .Q(\datapath.aluexecptions [0])
);

DFFPOSX1 _10955_ (
    .CLK(CLK_bF$buf68),
    .D(\controlunit.ebreak ),
    .Q(\datapath.aluexecptions [1])
);

DFFPOSX1 _10956_ (
    .CLK(CLK_bF$buf67),
    .D(\controlunit.ecall ),
    .Q(\datapath.aluexecptions [2])
);

DFFPOSX1 _10957_ (
    .CLK(CLK_bF$buf66),
    .D(\datapath.idinstr [0]),
    .Q(\datapath.aluinstr [0])
);

DFFPOSX1 _10958_ (
    .CLK(CLK_bF$buf65),
    .D(\datapath.idinstr [1]),
    .Q(\datapath.aluinstr [1])
);

DFFPOSX1 _10959_ (
    .CLK(CLK_bF$buf64),
    .D(\datapath.idinstr [2]),
    .Q(\datapath.aluinstr [2])
);

DFFPOSX1 _10960_ (
    .CLK(CLK_bF$buf63),
    .D(\datapath.idinstr [3]),
    .Q(\datapath.aluinstr [3])
);

DFFPOSX1 _10961_ (
    .CLK(CLK_bF$buf62),
    .D(\datapath.idinstr [4]),
    .Q(\datapath.aluinstr [4])
);

DFFPOSX1 _10962_ (
    .CLK(CLK_bF$buf61),
    .D(\datapath.idinstr [5]),
    .Q(\datapath.aluinstr [5])
);

DFFPOSX1 _10963_ (
    .CLK(CLK_bF$buf60),
    .D(\datapath.idinstr [6]),
    .Q(\datapath.aluinstr [6])
);

DFFPOSX1 _10964_ (
    .CLK(CLK_bF$buf59),
    .D(\datapath.idinstr [7]),
    .Q(\datapath.aluinstr [7])
);

DFFPOSX1 _10965_ (
    .CLK(CLK_bF$buf58),
    .D(\datapath.idinstr [8]),
    .Q(\datapath.aluinstr [8])
);

DFFPOSX1 _10966_ (
    .CLK(CLK_bF$buf57),
    .D(\datapath.idinstr [9]),
    .Q(\datapath.aluinstr [9])
);

DFFPOSX1 _10967_ (
    .CLK(CLK_bF$buf56),
    .D(\datapath.idinstr [10]),
    .Q(\datapath.aluinstr [10])
);

DFFPOSX1 _10968_ (
    .CLK(CLK_bF$buf55),
    .D(\datapath.idinstr [11]),
    .Q(\datapath.aluinstr [11])
);

DFFPOSX1 _10969_ (
    .CLK(CLK_bF$buf54),
    .D(\datapath.idinstr [12]),
    .Q(\datapath.aluinstr [12])
);

DFFPOSX1 _10970_ (
    .CLK(CLK_bF$buf53),
    .D(\datapath.idinstr [13]),
    .Q(\datapath.aluinstr [13])
);

DFFPOSX1 _10971_ (
    .CLK(CLK_bF$buf52),
    .D(\datapath.idinstr [14]),
    .Q(\datapath.aluinstr [14])
);

DFFPOSX1 _10972_ (
    .CLK(CLK_bF$buf51),
    .D(\datapath.idinstr_15_bF$buf54 ),
    .Q(\datapath.aluinstr [15])
);

DFFPOSX1 _10973_ (
    .CLK(CLK_bF$buf50),
    .D(\datapath.idinstr_16_bF$buf51 ),
    .Q(\datapath.aluinstr [16])
);

DFFPOSX1 _10974_ (
    .CLK(CLK_bF$buf49),
    .D(\datapath.idinstr_17_bF$buf15 ),
    .Q(\datapath.aluinstr [17])
);

DFFPOSX1 _10975_ (
    .CLK(CLK_bF$buf48),
    .D(\datapath.idinstr_18_bF$buf6 ),
    .Q(\datapath.aluinstr [18])
);

DFFPOSX1 _10976_ (
    .CLK(CLK_bF$buf47),
    .D(\datapath.idinstr_19_bF$buf5 ),
    .Q(\datapath.aluinstr [19])
);

DFFPOSX1 _10977_ (
    .CLK(CLK_bF$buf46),
    .D(\datapath.idinstr_20_bF$buf55 ),
    .Q(\datapath.aluinstr [20])
);

DFFPOSX1 _10978_ (
    .CLK(CLK_bF$buf45),
    .D(\datapath.idinstr_21_bF$buf51 ),
    .Q(\datapath.aluinstr [21])
);

DFFPOSX1 _10979_ (
    .CLK(CLK_bF$buf44),
    .D(\datapath.idinstr_22_bF$buf41 ),
    .Q(\datapath.aluinstr [22])
);

DFFPOSX1 _10980_ (
    .CLK(CLK_bF$buf43),
    .D(\datapath.idinstr_23_bF$buf6 ),
    .Q(\datapath.aluinstr [23])
);

DFFPOSX1 _10981_ (
    .CLK(CLK_bF$buf42),
    .D(\datapath.idinstr_24_bF$buf5 ),
    .Q(\datapath.aluinstr [24])
);

DFFPOSX1 _10982_ (
    .CLK(CLK_bF$buf41),
    .D(\datapath.idinstr [25]),
    .Q(\datapath.aluinstr [25])
);

DFFPOSX1 _10983_ (
    .CLK(CLK_bF$buf40),
    .D(\datapath.idinstr [26]),
    .Q(\datapath.aluinstr [26])
);

DFFPOSX1 _10984_ (
    .CLK(CLK_bF$buf39),
    .D(\datapath.idinstr [27]),
    .Q(\datapath.aluinstr [27])
);

DFFPOSX1 _10985_ (
    .CLK(CLK_bF$buf38),
    .D(\datapath.idinstr [28]),
    .Q(\datapath.aluinstr [28])
);

DFFPOSX1 _10986_ (
    .CLK(CLK_bF$buf37),
    .D(\datapath.idinstr [29]),
    .Q(\datapath.aluinstr [29])
);

DFFPOSX1 _10987_ (
    .CLK(CLK_bF$buf36),
    .D(\datapath.idinstr [30]),
    .Q(\datapath.aluinstr [30])
);

DFFPOSX1 _10988_ (
    .CLK(CLK_bF$buf35),
    .D(\datapath.idinstr [31]),
    .Q(\datapath.aluinstr [31])
);

DFFPOSX1 _10989_ (
    .CLK(CLK_bF$buf34),
    .D(\datapath.idpc_4 [0]),
    .Q(\datapath.alupc_4 [0])
);

DFFPOSX1 _10990_ (
    .CLK(CLK_bF$buf33),
    .D(\datapath.idpc_4 [1]),
    .Q(\datapath.alupc_4 [1])
);

DFFPOSX1 _10991_ (
    .CLK(CLK_bF$buf32),
    .D(\datapath.idpc_4 [2]),
    .Q(\datapath.alupc_4 [2])
);

DFFPOSX1 _10992_ (
    .CLK(CLK_bF$buf31),
    .D(\datapath.idpc_4 [3]),
    .Q(\datapath.alupc_4 [3])
);

DFFPOSX1 _10993_ (
    .CLK(CLK_bF$buf30),
    .D(\datapath.idpc_4 [4]),
    .Q(\datapath.alupc_4 [4])
);

DFFPOSX1 _10994_ (
    .CLK(CLK_bF$buf29),
    .D(\datapath.idpc_4 [5]),
    .Q(\datapath.alupc_4 [5])
);

DFFPOSX1 _10995_ (
    .CLK(CLK_bF$buf28),
    .D(\datapath.idpc_4 [6]),
    .Q(\datapath.alupc_4 [6])
);

DFFPOSX1 _10996_ (
    .CLK(CLK_bF$buf27),
    .D(\datapath.idpc_4 [7]),
    .Q(\datapath.alupc_4 [7])
);

DFFPOSX1 _10997_ (
    .CLK(CLK_bF$buf26),
    .D(\datapath.idpc_4 [8]),
    .Q(\datapath.alupc_4 [8])
);

DFFPOSX1 _10998_ (
    .CLK(CLK_bF$buf25),
    .D(\datapath.idpc_4 [9]),
    .Q(\datapath.alupc_4 [9])
);

DFFPOSX1 _10999_ (
    .CLK(CLK_bF$buf24),
    .D(\datapath.idpc_4 [10]),
    .Q(\datapath.alupc_4 [10])
);

DFFPOSX1 _11000_ (
    .CLK(CLK_bF$buf23),
    .D(\datapath.idpc_4 [11]),
    .Q(\datapath.alupc_4 [11])
);

DFFPOSX1 _11001_ (
    .CLK(CLK_bF$buf22),
    .D(\datapath.idpc_4 [12]),
    .Q(\datapath.alupc_4 [12])
);

DFFPOSX1 _11002_ (
    .CLK(CLK_bF$buf21),
    .D(\datapath.idpc_4 [13]),
    .Q(\datapath.alupc_4 [13])
);

DFFPOSX1 _11003_ (
    .CLK(CLK_bF$buf20),
    .D(\datapath.idpc_4 [14]),
    .Q(\datapath.alupc_4 [14])
);

DFFPOSX1 _11004_ (
    .CLK(CLK_bF$buf19),
    .D(\datapath.idpc_4 [15]),
    .Q(\datapath.alupc_4 [15])
);

DFFPOSX1 _11005_ (
    .CLK(CLK_bF$buf18),
    .D(\datapath.idpc_4 [16]),
    .Q(\datapath.alupc_4 [16])
);

DFFPOSX1 _11006_ (
    .CLK(CLK_bF$buf17),
    .D(\datapath.idpc_4 [17]),
    .Q(\datapath.alupc_4 [17])
);

DFFPOSX1 _11007_ (
    .CLK(CLK_bF$buf16),
    .D(\datapath.idpc_4 [18]),
    .Q(\datapath.alupc_4 [18])
);

DFFPOSX1 _11008_ (
    .CLK(CLK_bF$buf15),
    .D(\datapath.idpc_4 [19]),
    .Q(\datapath.alupc_4 [19])
);

DFFPOSX1 _11009_ (
    .CLK(CLK_bF$buf14),
    .D(\datapath.idpc_4 [20]),
    .Q(\datapath.alupc_4 [20])
);

DFFPOSX1 _11010_ (
    .CLK(CLK_bF$buf13),
    .D(\datapath.idpc_4 [21]),
    .Q(\datapath.alupc_4 [21])
);

DFFPOSX1 _11011_ (
    .CLK(CLK_bF$buf12),
    .D(\datapath.idpc_4 [22]),
    .Q(\datapath.alupc_4 [22])
);

DFFPOSX1 _11012_ (
    .CLK(CLK_bF$buf11),
    .D(\datapath.idpc_4 [23]),
    .Q(\datapath.alupc_4 [23])
);

DFFPOSX1 _11013_ (
    .CLK(CLK_bF$buf10),
    .D(\datapath.idpc_4 [24]),
    .Q(\datapath.alupc_4 [24])
);

DFFPOSX1 _11014_ (
    .CLK(CLK_bF$buf9),
    .D(\datapath.idpc_4 [25]),
    .Q(\datapath.alupc_4 [25])
);

DFFPOSX1 _11015_ (
    .CLK(CLK_bF$buf8),
    .D(\datapath.idpc_4 [26]),
    .Q(\datapath.alupc_4 [26])
);

DFFPOSX1 _11016_ (
    .CLK(CLK_bF$buf7),
    .D(\datapath.idpc_4 [27]),
    .Q(\datapath.alupc_4 [27])
);

DFFPOSX1 _11017_ (
    .CLK(CLK_bF$buf6),
    .D(\datapath.idpc_4 [28]),
    .Q(\datapath.alupc_4 [28])
);

DFFPOSX1 _11018_ (
    .CLK(CLK_bF$buf5),
    .D(\datapath.idpc_4 [29]),
    .Q(\datapath.alupc_4 [29])
);

DFFPOSX1 _11019_ (
    .CLK(CLK_bF$buf4),
    .D(\datapath.idpc_4 [30]),
    .Q(\datapath.alupc_4 [30])
);

DFFPOSX1 _11020_ (
    .CLK(CLK_bF$buf3),
    .D(\datapath.idpc_4 [31]),
    .Q(\datapath.alupc_4 [31])
);

DFFPOSX1 _11021_ (
    .CLK(CLK_bF$buf2),
    .D(\datapath.idpc [0]),
    .Q(\datapath.alupc [0])
);

DFFPOSX1 _11022_ (
    .CLK(CLK_bF$buf1),
    .D(\datapath.idpc [1]),
    .Q(\datapath.alupc [1])
);

DFFPOSX1 _11023_ (
    .CLK(CLK_bF$buf0),
    .D(\datapath.idpc [2]),
    .Q(\datapath.alupc [2])
);

DFFPOSX1 _11024_ (
    .CLK(CLK_bF$buf151),
    .D(\datapath.idpc [3]),
    .Q(\datapath.alupc [3])
);

DFFPOSX1 _11025_ (
    .CLK(CLK_bF$buf150),
    .D(\datapath.idpc [4]),
    .Q(\datapath.alupc [4])
);

DFFPOSX1 _11026_ (
    .CLK(CLK_bF$buf149),
    .D(\datapath.idpc [5]),
    .Q(\datapath.alupc [5])
);

DFFPOSX1 _11027_ (
    .CLK(CLK_bF$buf148),
    .D(\datapath.idpc [6]),
    .Q(\datapath.alupc [6])
);

DFFPOSX1 _11028_ (
    .CLK(CLK_bF$buf147),
    .D(\datapath.idpc [7]),
    .Q(\datapath.alupc [7])
);

DFFPOSX1 _11029_ (
    .CLK(CLK_bF$buf146),
    .D(\datapath.idpc [8]),
    .Q(\datapath.alupc [8])
);

DFFPOSX1 _11030_ (
    .CLK(CLK_bF$buf145),
    .D(\datapath.idpc [9]),
    .Q(\datapath.alupc [9])
);

DFFPOSX1 _11031_ (
    .CLK(CLK_bF$buf144),
    .D(\datapath.idpc [10]),
    .Q(\datapath.alupc [10])
);

DFFPOSX1 _11032_ (
    .CLK(CLK_bF$buf143),
    .D(\datapath.idpc [11]),
    .Q(\datapath.alupc [11])
);

DFFPOSX1 _11033_ (
    .CLK(CLK_bF$buf142),
    .D(\datapath.idpc [12]),
    .Q(\datapath.alupc [12])
);

DFFPOSX1 _11034_ (
    .CLK(CLK_bF$buf141),
    .D(\datapath.idpc [13]),
    .Q(\datapath.alupc [13])
);

DFFPOSX1 _11035_ (
    .CLK(CLK_bF$buf140),
    .D(\datapath.idpc [14]),
    .Q(\datapath.alupc [14])
);

DFFPOSX1 _11036_ (
    .CLK(CLK_bF$buf139),
    .D(\datapath.idpc [15]),
    .Q(\datapath.alupc [15])
);

DFFPOSX1 _11037_ (
    .CLK(CLK_bF$buf138),
    .D(\datapath.idpc [16]),
    .Q(\datapath.alupc [16])
);

DFFPOSX1 _11038_ (
    .CLK(CLK_bF$buf137),
    .D(\datapath.idpc [17]),
    .Q(\datapath.alupc [17])
);

DFFPOSX1 _11039_ (
    .CLK(CLK_bF$buf136),
    .D(\datapath.idpc [18]),
    .Q(\datapath.alupc [18])
);

DFFPOSX1 _11040_ (
    .CLK(CLK_bF$buf135),
    .D(\datapath.idpc [19]),
    .Q(\datapath.alupc [19])
);

DFFPOSX1 _11041_ (
    .CLK(CLK_bF$buf134),
    .D(\datapath.idpc [20]),
    .Q(\datapath.alupc [20])
);

DFFPOSX1 _11042_ (
    .CLK(CLK_bF$buf133),
    .D(\datapath.idpc [21]),
    .Q(\datapath.alupc [21])
);

DFFPOSX1 _11043_ (
    .CLK(CLK_bF$buf132),
    .D(\datapath.idpc [22]),
    .Q(\datapath.alupc [22])
);

DFFPOSX1 _11044_ (
    .CLK(CLK_bF$buf131),
    .D(\datapath.idpc [23]),
    .Q(\datapath.alupc [23])
);

DFFPOSX1 _11045_ (
    .CLK(CLK_bF$buf130),
    .D(\datapath.idpc [24]),
    .Q(\datapath.alupc [24])
);

DFFPOSX1 _11046_ (
    .CLK(CLK_bF$buf129),
    .D(\datapath.idpc [25]),
    .Q(\datapath.alupc [25])
);

DFFPOSX1 _11047_ (
    .CLK(CLK_bF$buf128),
    .D(\datapath.idpc [26]),
    .Q(\datapath.alupc [26])
);

DFFPOSX1 _11048_ (
    .CLK(CLK_bF$buf127),
    .D(\datapath.idpc [27]),
    .Q(\datapath.alupc [27])
);

DFFPOSX1 _11049_ (
    .CLK(CLK_bF$buf126),
    .D(\datapath.idpc [28]),
    .Q(\datapath.alupc [28])
);

DFFPOSX1 _11050_ (
    .CLK(CLK_bF$buf125),
    .D(\datapath.idpc [29]),
    .Q(\datapath.alupc [29])
);

DFFPOSX1 _11051_ (
    .CLK(CLK_bF$buf124),
    .D(\datapath.idpc [30]),
    .Q(\datapath.alupc [30])
);

DFFPOSX1 _11052_ (
    .CLK(CLK_bF$buf123),
    .D(\datapath.idpc [31]),
    .Q(\datapath.alupc [31])
);

DFFPOSX1 _11053_ (
    .CLK(CLK_bF$buf122),
    .D(\datapath._05_ [0]),
    .Q(\datapath.idinstr [0])
);

DFFPOSX1 _11054_ (
    .CLK(CLK_bF$buf121),
    .D(\datapath._05_ [1]),
    .Q(\datapath.idinstr [1])
);

DFFPOSX1 _11055_ (
    .CLK(CLK_bF$buf120),
    .D(\datapath._05_ [2]),
    .Q(\datapath.idinstr [2])
);

DFFPOSX1 _11056_ (
    .CLK(CLK_bF$buf119),
    .D(\datapath._05_ [3]),
    .Q(\datapath.idinstr [3])
);

DFFPOSX1 _11057_ (
    .CLK(CLK_bF$buf118),
    .D(\datapath._05_ [4]),
    .Q(\datapath.idinstr [4])
);

DFFPOSX1 _11058_ (
    .CLK(CLK_bF$buf117),
    .D(\datapath._05_ [5]),
    .Q(\datapath.idinstr [5])
);

DFFPOSX1 _11059_ (
    .CLK(CLK_bF$buf116),
    .D(\datapath._05_ [6]),
    .Q(\datapath.idinstr [6])
);

DFFPOSX1 _11060_ (
    .CLK(CLK_bF$buf115),
    .D(\datapath._05_ [7]),
    .Q(\datapath.idinstr [7])
);

DFFPOSX1 _11061_ (
    .CLK(CLK_bF$buf114),
    .D(\datapath._05_ [8]),
    .Q(\datapath.idinstr [8])
);

DFFPOSX1 _11062_ (
    .CLK(CLK_bF$buf113),
    .D(\datapath._05_ [9]),
    .Q(\datapath.idinstr [9])
);

DFFPOSX1 _11063_ (
    .CLK(CLK_bF$buf112),
    .D(\datapath._05_ [10]),
    .Q(\datapath.idinstr [10])
);

DFFPOSX1 _11064_ (
    .CLK(CLK_bF$buf111),
    .D(\datapath._05_ [11]),
    .Q(\datapath.idinstr [11])
);

DFFPOSX1 _11065_ (
    .CLK(CLK_bF$buf110),
    .D(\datapath._05_ [12]),
    .Q(\datapath.idinstr [12])
);

DFFPOSX1 _11066_ (
    .CLK(CLK_bF$buf109),
    .D(\datapath._05_ [13]),
    .Q(\datapath.idinstr [13])
);

DFFPOSX1 _11067_ (
    .CLK(CLK_bF$buf108),
    .D(\datapath._05_ [14]),
    .Q(\datapath.idinstr [14])
);

DFFPOSX1 _11068_ (
    .CLK(CLK_bF$buf107),
    .D(\datapath._05_ [15]),
    .Q(\datapath.idinstr [15])
);

DFFPOSX1 _11069_ (
    .CLK(CLK_bF$buf106),
    .D(\datapath._05_ [16]),
    .Q(\datapath.idinstr [16])
);

DFFPOSX1 _11070_ (
    .CLK(CLK_bF$buf105),
    .D(\datapath._05_ [17]),
    .Q(\datapath.idinstr [17])
);

DFFPOSX1 _11071_ (
    .CLK(CLK_bF$buf104),
    .D(\datapath._05_ [18]),
    .Q(\datapath.idinstr [18])
);

DFFPOSX1 _11072_ (
    .CLK(CLK_bF$buf103),
    .D(\datapath._05_ [19]),
    .Q(\datapath.idinstr [19])
);

DFFPOSX1 _11073_ (
    .CLK(CLK_bF$buf102),
    .D(\datapath._05_ [20]),
    .Q(\datapath.idinstr [20])
);

DFFPOSX1 _11074_ (
    .CLK(CLK_bF$buf101),
    .D(\datapath._05_ [21]),
    .Q(\datapath.idinstr [21])
);

DFFPOSX1 _11075_ (
    .CLK(CLK_bF$buf100),
    .D(\datapath._05_ [22]),
    .Q(\datapath.idinstr [22])
);

DFFPOSX1 _11076_ (
    .CLK(CLK_bF$buf99),
    .D(\datapath._05_ [23]),
    .Q(\datapath.idinstr [23])
);

DFFPOSX1 _11077_ (
    .CLK(CLK_bF$buf98),
    .D(\datapath._05_ [24]),
    .Q(\datapath.idinstr [24])
);

DFFPOSX1 _11078_ (
    .CLK(CLK_bF$buf97),
    .D(\datapath._05_ [25]),
    .Q(\datapath.idinstr [25])
);

DFFPOSX1 _11079_ (
    .CLK(CLK_bF$buf96),
    .D(\datapath._05_ [26]),
    .Q(\datapath.idinstr [26])
);

DFFPOSX1 _11080_ (
    .CLK(CLK_bF$buf95),
    .D(\datapath._05_ [27]),
    .Q(\datapath.idinstr [27])
);

DFFPOSX1 _11081_ (
    .CLK(CLK_bF$buf94),
    .D(\datapath._05_ [28]),
    .Q(\datapath.idinstr [28])
);

DFFPOSX1 _11082_ (
    .CLK(CLK_bF$buf93),
    .D(\datapath._05_ [29]),
    .Q(\datapath.idinstr [29])
);

DFFPOSX1 _11083_ (
    .CLK(CLK_bF$buf92),
    .D(\datapath._05_ [30]),
    .Q(\datapath.idinstr [30])
);

DFFPOSX1 _11084_ (
    .CLK(CLK_bF$buf91),
    .D(\datapath._05_ [31]),
    .Q(\datapath.idinstr [31])
);

DFFPOSX1 _11085_ (
    .CLK(CLK_bF$buf90),
    .D(\datapath._04_ [0]),
    .Q(\datapath.idpc_4 [0])
);

DFFPOSX1 _11086_ (
    .CLK(CLK_bF$buf89),
    .D(\datapath._04_ [1]),
    .Q(\datapath.idpc_4 [1])
);

DFFPOSX1 _11087_ (
    .CLK(CLK_bF$buf88),
    .D(\datapath._04_ [2]),
    .Q(\datapath.idpc_4 [2])
);

DFFPOSX1 _11088_ (
    .CLK(CLK_bF$buf87),
    .D(\datapath._04_ [3]),
    .Q(\datapath.idpc_4 [3])
);

DFFPOSX1 _11089_ (
    .CLK(CLK_bF$buf86),
    .D(\datapath._04_ [4]),
    .Q(\datapath.idpc_4 [4])
);

DFFPOSX1 _11090_ (
    .CLK(CLK_bF$buf85),
    .D(\datapath._04_ [5]),
    .Q(\datapath.idpc_4 [5])
);

DFFPOSX1 _11091_ (
    .CLK(CLK_bF$buf84),
    .D(\datapath._04_ [6]),
    .Q(\datapath.idpc_4 [6])
);

DFFPOSX1 _11092_ (
    .CLK(CLK_bF$buf83),
    .D(\datapath._04_ [7]),
    .Q(\datapath.idpc_4 [7])
);

DFFPOSX1 _11093_ (
    .CLK(CLK_bF$buf82),
    .D(\datapath._04_ [8]),
    .Q(\datapath.idpc_4 [8])
);

DFFPOSX1 _11094_ (
    .CLK(CLK_bF$buf81),
    .D(\datapath._04_ [9]),
    .Q(\datapath.idpc_4 [9])
);

DFFPOSX1 _11095_ (
    .CLK(CLK_bF$buf80),
    .D(\datapath._04_ [10]),
    .Q(\datapath.idpc_4 [10])
);

DFFPOSX1 _11096_ (
    .CLK(CLK_bF$buf79),
    .D(\datapath._04_ [11]),
    .Q(\datapath.idpc_4 [11])
);

DFFPOSX1 _11097_ (
    .CLK(CLK_bF$buf78),
    .D(\datapath._04_ [12]),
    .Q(\datapath.idpc_4 [12])
);

DFFPOSX1 _11098_ (
    .CLK(CLK_bF$buf77),
    .D(\datapath._04_ [13]),
    .Q(\datapath.idpc_4 [13])
);

DFFPOSX1 _11099_ (
    .CLK(CLK_bF$buf76),
    .D(\datapath._04_ [14]),
    .Q(\datapath.idpc_4 [14])
);

DFFPOSX1 _11100_ (
    .CLK(CLK_bF$buf75),
    .D(\datapath._04_ [15]),
    .Q(\datapath.idpc_4 [15])
);

DFFPOSX1 _11101_ (
    .CLK(CLK_bF$buf74),
    .D(\datapath._04_ [16]),
    .Q(\datapath.idpc_4 [16])
);

DFFPOSX1 _11102_ (
    .CLK(CLK_bF$buf73),
    .D(\datapath._04_ [17]),
    .Q(\datapath.idpc_4 [17])
);

DFFPOSX1 _11103_ (
    .CLK(CLK_bF$buf72),
    .D(\datapath._04_ [18]),
    .Q(\datapath.idpc_4 [18])
);

DFFPOSX1 _11104_ (
    .CLK(CLK_bF$buf71),
    .D(\datapath._04_ [19]),
    .Q(\datapath.idpc_4 [19])
);

DFFPOSX1 _11105_ (
    .CLK(CLK_bF$buf70),
    .D(\datapath._04_ [20]),
    .Q(\datapath.idpc_4 [20])
);

DFFPOSX1 _11106_ (
    .CLK(CLK_bF$buf69),
    .D(\datapath._04_ [21]),
    .Q(\datapath.idpc_4 [21])
);

DFFPOSX1 _11107_ (
    .CLK(CLK_bF$buf68),
    .D(\datapath._04_ [22]),
    .Q(\datapath.idpc_4 [22])
);

DFFPOSX1 _11108_ (
    .CLK(CLK_bF$buf67),
    .D(\datapath._04_ [23]),
    .Q(\datapath.idpc_4 [23])
);

DFFPOSX1 _11109_ (
    .CLK(CLK_bF$buf66),
    .D(\datapath._04_ [24]),
    .Q(\datapath.idpc_4 [24])
);

DFFPOSX1 _11110_ (
    .CLK(CLK_bF$buf65),
    .D(\datapath._04_ [25]),
    .Q(\datapath.idpc_4 [25])
);

DFFPOSX1 _11111_ (
    .CLK(CLK_bF$buf64),
    .D(\datapath._04_ [26]),
    .Q(\datapath.idpc_4 [26])
);

DFFPOSX1 _11112_ (
    .CLK(CLK_bF$buf63),
    .D(\datapath._04_ [27]),
    .Q(\datapath.idpc_4 [27])
);

DFFPOSX1 _11113_ (
    .CLK(CLK_bF$buf62),
    .D(\datapath._04_ [28]),
    .Q(\datapath.idpc_4 [28])
);

DFFPOSX1 _11114_ (
    .CLK(CLK_bF$buf61),
    .D(\datapath._04_ [29]),
    .Q(\datapath.idpc_4 [29])
);

DFFPOSX1 _11115_ (
    .CLK(CLK_bF$buf60),
    .D(\datapath._04_ [30]),
    .Q(\datapath.idpc_4 [30])
);

DFFPOSX1 _11116_ (
    .CLK(CLK_bF$buf59),
    .D(\datapath._04_ [31]),
    .Q(\datapath.idpc_4 [31])
);

DFFPOSX1 _11117_ (
    .CLK(CLK_bF$buf58),
    .D(\datapath._03_ [0]),
    .Q(\datapath.idpc [0])
);

DFFPOSX1 _11118_ (
    .CLK(CLK_bF$buf57),
    .D(\datapath._03_ [1]),
    .Q(\datapath.idpc [1])
);

DFFPOSX1 _11119_ (
    .CLK(CLK_bF$buf56),
    .D(\datapath._03_ [2]),
    .Q(\datapath.idpc [2])
);

DFFPOSX1 _11120_ (
    .CLK(CLK_bF$buf55),
    .D(\datapath._03_ [3]),
    .Q(\datapath.idpc [3])
);

DFFPOSX1 _11121_ (
    .CLK(CLK_bF$buf54),
    .D(\datapath._03_ [4]),
    .Q(\datapath.idpc [4])
);

DFFPOSX1 _11122_ (
    .CLK(CLK_bF$buf53),
    .D(\datapath._03_ [5]),
    .Q(\datapath.idpc [5])
);

DFFPOSX1 _11123_ (
    .CLK(CLK_bF$buf52),
    .D(\datapath._03_ [6]),
    .Q(\datapath.idpc [6])
);

DFFPOSX1 _11124_ (
    .CLK(CLK_bF$buf51),
    .D(\datapath._03_ [7]),
    .Q(\datapath.idpc [7])
);

DFFPOSX1 _11125_ (
    .CLK(CLK_bF$buf50),
    .D(\datapath._03_ [8]),
    .Q(\datapath.idpc [8])
);

DFFPOSX1 _11126_ (
    .CLK(CLK_bF$buf49),
    .D(\datapath._03_ [9]),
    .Q(\datapath.idpc [9])
);

DFFPOSX1 _11127_ (
    .CLK(CLK_bF$buf48),
    .D(\datapath._03_ [10]),
    .Q(\datapath.idpc [10])
);

DFFPOSX1 _11128_ (
    .CLK(CLK_bF$buf47),
    .D(\datapath._03_ [11]),
    .Q(\datapath.idpc [11])
);

DFFPOSX1 _11129_ (
    .CLK(CLK_bF$buf46),
    .D(\datapath._03_ [12]),
    .Q(\datapath.idpc [12])
);

DFFPOSX1 _11130_ (
    .CLK(CLK_bF$buf45),
    .D(\datapath._03_ [13]),
    .Q(\datapath.idpc [13])
);

DFFPOSX1 _11131_ (
    .CLK(CLK_bF$buf44),
    .D(\datapath._03_ [14]),
    .Q(\datapath.idpc [14])
);

DFFPOSX1 _11132_ (
    .CLK(CLK_bF$buf43),
    .D(\datapath._03_ [15]),
    .Q(\datapath.idpc [15])
);

DFFPOSX1 _11133_ (
    .CLK(CLK_bF$buf42),
    .D(\datapath._03_ [16]),
    .Q(\datapath.idpc [16])
);

DFFPOSX1 _11134_ (
    .CLK(CLK_bF$buf41),
    .D(\datapath._03_ [17]),
    .Q(\datapath.idpc [17])
);

DFFPOSX1 _11135_ (
    .CLK(CLK_bF$buf40),
    .D(\datapath._03_ [18]),
    .Q(\datapath.idpc [18])
);

DFFPOSX1 _11136_ (
    .CLK(CLK_bF$buf39),
    .D(\datapath._03_ [19]),
    .Q(\datapath.idpc [19])
);

DFFPOSX1 _11137_ (
    .CLK(CLK_bF$buf38),
    .D(\datapath._03_ [20]),
    .Q(\datapath.idpc [20])
);

DFFPOSX1 _11138_ (
    .CLK(CLK_bF$buf37),
    .D(\datapath._03_ [21]),
    .Q(\datapath.idpc [21])
);

DFFPOSX1 _11139_ (
    .CLK(CLK_bF$buf36),
    .D(\datapath._03_ [22]),
    .Q(\datapath.idpc [22])
);

DFFPOSX1 _11140_ (
    .CLK(CLK_bF$buf35),
    .D(\datapath._03_ [23]),
    .Q(\datapath.idpc [23])
);

DFFPOSX1 _11141_ (
    .CLK(CLK_bF$buf34),
    .D(\datapath._03_ [24]),
    .Q(\datapath.idpc [24])
);

DFFPOSX1 _11142_ (
    .CLK(CLK_bF$buf33),
    .D(\datapath._03_ [25]),
    .Q(\datapath.idpc [25])
);

DFFPOSX1 _11143_ (
    .CLK(CLK_bF$buf32),
    .D(\datapath._03_ [26]),
    .Q(\datapath.idpc [26])
);

DFFPOSX1 _11144_ (
    .CLK(CLK_bF$buf31),
    .D(\datapath._03_ [27]),
    .Q(\datapath.idpc [27])
);

DFFPOSX1 _11145_ (
    .CLK(CLK_bF$buf30),
    .D(\datapath._03_ [28]),
    .Q(\datapath.idpc [28])
);

DFFPOSX1 _11146_ (
    .CLK(CLK_bF$buf29),
    .D(\datapath._03_ [29]),
    .Q(\datapath.idpc [29])
);

DFFPOSX1 _11147_ (
    .CLK(CLK_bF$buf28),
    .D(\datapath._03_ [30]),
    .Q(\datapath.idpc [30])
);

DFFPOSX1 _11148_ (
    .CLK(CLK_bF$buf27),
    .D(\datapath._03_ [31]),
    .Q(\datapath.idpc [31])
);

NAND2X1 _11149_ (
    .A(\datapath.alu.a [31]),
    .B(\datapath.alu.b [31]),
    .Y(_903_)
);

INVX2 _11150_ (
    .A(\datapath.alu.a [31]),
    .Y(_913_)
);

INVX1 _11151_ (
    .A(\datapath.alu.b [31]),
    .Y(_924_)
);

NAND2X1 _11152_ (
    .A(_913_),
    .B(_924_),
    .Y(_935_)
);

NAND2X1 _11153_ (
    .A(_903_),
    .B(_935_),
    .Y(_946_)
);

NAND2X1 _11154_ (
    .A(\datapath.alu.a [23]),
    .B(\datapath.alu.b [23]),
    .Y(_956_)
);

INVX2 _11155_ (
    .A(\datapath.alu.a [23]),
    .Y(_967_)
);

INVX1 _11156_ (
    .A(\datapath.alu.b [23]),
    .Y(_978_)
);

NAND2X1 _11157_ (
    .A(_967_),
    .B(_978_),
    .Y(_989_)
);

NAND2X1 _11158_ (
    .A(_956_),
    .B(_989_),
    .Y(_1000_)
);

INVX2 _11159_ (
    .A(\datapath.alu.a [22]),
    .Y(_1010_)
);

INVX1 _11160_ (
    .A(\datapath.alu.b [22]),
    .Y(_1021_)
);

NAND2X1 _11161_ (
    .A(_1010_),
    .B(_1021_),
    .Y(_1032_)
);

NAND2X1 _11162_ (
    .A(\datapath.alu.a [22]),
    .B(\datapath.alu.b [22]),
    .Y(_1042_)
);

NAND2X1 _11163_ (
    .A(_1042_),
    .B(_1032_),
    .Y(_1053_)
);

NAND2X1 _11164_ (
    .A(_1000_),
    .B(_1053_),
    .Y(_1064_)
);

NAND2X1 _11165_ (
    .A(\datapath.alu.a [21]),
    .B(\datapath.alu.b [21]),
    .Y(_1075_)
);

INVX2 _11166_ (
    .A(\datapath.alu.a [21]),
    .Y(_1086_)
);

INVX1 _11167_ (
    .A(\datapath.alu.b [21]),
    .Y(_1096_)
);

NAND2X1 _11168_ (
    .A(_1086_),
    .B(_1096_),
    .Y(_1107_)
);

NAND2X1 _11169_ (
    .A(_1075_),
    .B(_1107_),
    .Y(_1118_)
);

INVX2 _11170_ (
    .A(\datapath.alu.a [20]),
    .Y(_1128_)
);

INVX1 _11171_ (
    .A(\datapath.alu.b [20]),
    .Y(_1139_)
);

NAND2X1 _11172_ (
    .A(_1128_),
    .B(_1139_),
    .Y(_1150_)
);

NAND2X1 _11173_ (
    .A(\datapath.alu.a [20]),
    .B(\datapath.alu.b [20]),
    .Y(_1161_)
);

NAND2X1 _11174_ (
    .A(_1161_),
    .B(_1150_),
    .Y(_1172_)
);

NAND2X1 _11175_ (
    .A(_1118_),
    .B(_1172_),
    .Y(_1183_)
);

NOR2X1 _11176_ (
    .A(_1064_),
    .B(_1183_),
    .Y(_1193_)
);

INVX1 _11177_ (
    .A(\datapath.alu.a [19]),
    .Y(_1204_)
);

INVX1 _11178_ (
    .A(\datapath.alu.b [19]),
    .Y(_1215_)
);

NOR2X1 _11179_ (
    .A(_1204_),
    .B(_1215_),
    .Y(_1225_)
);

NOR2X1 _11180_ (
    .A(\datapath.alu.a [19]),
    .B(\datapath.alu.b [19]),
    .Y(_1236_)
);

INVX2 _11181_ (
    .A(\datapath.alu.a [18]),
    .Y(_1247_)
);

INVX1 _11182_ (
    .A(\datapath.alu.b [18]),
    .Y(_1258_)
);

NAND2X1 _11183_ (
    .A(_1247_),
    .B(_1258_),
    .Y(_1268_)
);

NAND2X1 _11184_ (
    .A(\datapath.alu.a [18]),
    .B(\datapath.alu.b [18]),
    .Y(_1279_)
);

NAND2X1 _11185_ (
    .A(_1279_),
    .B(_1268_),
    .Y(_1290_)
);

OAI21X1 _11186_ (
    .A(_1225_),
    .B(_1236_),
    .C(_1290_),
    .Y(_1300_)
);

NAND2X1 _11187_ (
    .A(\datapath.alu.a [17]),
    .B(\datapath.alu.b [17]),
    .Y(_1311_)
);

INVX2 _11188_ (
    .A(\datapath.alu.a [17]),
    .Y(_1322_)
);

INVX2 _11189_ (
    .A(\datapath.alu.b [17]),
    .Y(_1333_)
);

NAND2X1 _11190_ (
    .A(_1322_),
    .B(_1333_),
    .Y(_1343_)
);

NAND2X1 _11191_ (
    .A(_1311_),
    .B(_1343_),
    .Y(_1354_)
);

INVX2 _11192_ (
    .A(\datapath.alu.a [16]),
    .Y(_1365_)
);

INVX1 _11193_ (
    .A(\datapath.alu.b [16]),
    .Y(_1375_)
);

NAND2X1 _11194_ (
    .A(_1365_),
    .B(_1375_),
    .Y(_1386_)
);

NAND2X1 _11195_ (
    .A(\datapath.alu.a [16]),
    .B(\datapath.alu.b [16]),
    .Y(_1397_)
);

NAND2X1 _11196_ (
    .A(_1397_),
    .B(_1386_),
    .Y(_1408_)
);

NAND2X1 _11197_ (
    .A(_1354_),
    .B(_1408_),
    .Y(_1418_)
);

NOR2X1 _11198_ (
    .A(_1418_),
    .B(_1300_),
    .Y(_1429_)
);

NAND2X1 _11199_ (
    .A(_1193_),
    .B(_1429_),
    .Y(_1440_)
);

INVX2 _11200_ (
    .A(\datapath.alu.a [30]),
    .Y(_1450_)
);

INVX1 _11201_ (
    .A(\datapath.alu.b [30]),
    .Y(_1461_)
);

NAND2X1 _11202_ (
    .A(_1450_),
    .B(_1461_),
    .Y(_1472_)
);

NAND2X1 _11203_ (
    .A(\datapath.alu.a [30]),
    .B(\datapath.alu.b [30]),
    .Y(_1483_)
);

NAND2X1 _11204_ (
    .A(_1483_),
    .B(_1472_),
    .Y(_1494_)
);

NAND2X1 _11205_ (
    .A(_946_),
    .B(_1494_),
    .Y(_1504_)
);

NAND2X1 _11206_ (
    .A(\datapath.alu.a [29]),
    .B(\datapath.alu.b [29]),
    .Y(_1515_)
);

INVX2 _11207_ (
    .A(\datapath.alu.a [29]),
    .Y(_1526_)
);

INVX1 _11208_ (
    .A(\datapath.alu.b [29]),
    .Y(_1536_)
);

NAND2X1 _11209_ (
    .A(_1526_),
    .B(_1536_),
    .Y(_1547_)
);

NAND2X1 _11210_ (
    .A(_1515_),
    .B(_1547_),
    .Y(_1558_)
);

INVX2 _11211_ (
    .A(\datapath.alu.a [28]),
    .Y(_1568_)
);

INVX1 _11212_ (
    .A(\datapath.alu.b [28]),
    .Y(_1579_)
);

NAND2X1 _11213_ (
    .A(_1568_),
    .B(_1579_),
    .Y(_1590_)
);

NAND2X1 _11214_ (
    .A(\datapath.alu.a [28]),
    .B(\datapath.alu.b [28]),
    .Y(_1601_)
);

NAND2X1 _11215_ (
    .A(_1601_),
    .B(_1590_),
    .Y(_1611_)
);

NAND2X1 _11216_ (
    .A(_1558_),
    .B(_1611_),
    .Y(_1622_)
);

NOR2X1 _11217_ (
    .A(_1504_),
    .B(_1622_),
    .Y(_1633_)
);

INVX2 _11218_ (
    .A(\datapath.alu.a [27]),
    .Y(_1643_)
);

INVX1 _11219_ (
    .A(\datapath.alu.b [27]),
    .Y(_1654_)
);

NOR2X1 _11220_ (
    .A(_1643_),
    .B(_1654_),
    .Y(_1665_)
);

NOR2X1 _11221_ (
    .A(\datapath.alu.a [27]),
    .B(\datapath.alu.b [27]),
    .Y(_1676_)
);

INVX2 _11222_ (
    .A(\datapath.alu.a [26]),
    .Y(_1686_)
);

INVX1 _11223_ (
    .A(\datapath.alu.b [26]),
    .Y(_1697_)
);

NAND2X1 _11224_ (
    .A(_1686_),
    .B(_1697_),
    .Y(_1708_)
);

NAND2X1 _11225_ (
    .A(\datapath.alu.a [26]),
    .B(\datapath.alu.b [26]),
    .Y(_1718_)
);

NAND2X1 _11226_ (
    .A(_1718_),
    .B(_1708_),
    .Y(_1729_)
);

OAI21X1 _11227_ (
    .A(_1665_),
    .B(_1676_),
    .C(_1729_),
    .Y(_1740_)
);

NAND2X1 _11228_ (
    .A(\datapath.alu.a [25]),
    .B(\datapath.alu.b [25]),
    .Y(_1750_)
);

INVX2 _11229_ (
    .A(\datapath.alu.a [25]),
    .Y(_1760_)
);

INVX1 _11230_ (
    .A(\datapath.alu.b [25]),
    .Y(_1761_)
);

NAND2X1 _11231_ (
    .A(_1760_),
    .B(_1761_),
    .Y(_1762_)
);

NAND2X1 _11232_ (
    .A(_1750_),
    .B(_1762_),
    .Y(_1763_)
);

NOR2X1 _11233_ (
    .A(\datapath.alu.a [24]),
    .B(\datapath.alu.b [24]),
    .Y(_1764_)
);

INVX2 _11234_ (
    .A(\datapath.alu.a [24]),
    .Y(_1765_)
);

INVX1 _11235_ (
    .A(\datapath.alu.b [24]),
    .Y(_1766_)
);

NOR2X1 _11236_ (
    .A(_1765_),
    .B(_1766_),
    .Y(_1767_)
);

OAI21X1 _11237_ (
    .A(_1764_),
    .B(_1767_),
    .C(_1763_),
    .Y(_1768_)
);

NOR2X1 _11238_ (
    .A(_1740_),
    .B(_1768_),
    .Y(_1769_)
);

NAND2X1 _11239_ (
    .A(_1633_),
    .B(_1769_),
    .Y(_1770_)
);

NOR2X1 _11240_ (
    .A(_1440_),
    .B(_1770_),
    .Y(_1771_)
);

NAND2X1 _11241_ (
    .A(\datapath.alu.a [15]),
    .B(\datapath.alu.b [15]),
    .Y(_1772_)
);

INVX2 _11242_ (
    .A(\datapath.alu.a [15]),
    .Y(_1773_)
);

INVX2 _11243_ (
    .A(\datapath.alu.b [15]),
    .Y(_1774_)
);

NAND2X1 _11244_ (
    .A(_1773_),
    .B(_1774_),
    .Y(_1775_)
);

NAND2X1 _11245_ (
    .A(_1772_),
    .B(_1775_),
    .Y(_1776_)
);

INVX2 _11246_ (
    .A(\datapath.alu.a [14]),
    .Y(_1777_)
);

NAND2X1 _11247_ (
    .A(\datapath.alu.b [14]),
    .B(_1777_),
    .Y(_1778_)
);

INVX1 _11248_ (
    .A(\datapath.alu.b [14]),
    .Y(_1779_)
);

NAND2X1 _11249_ (
    .A(\datapath.alu.a [14]),
    .B(_1779_),
    .Y(_1780_)
);

AND2X2 _11250_ (
    .A(_1778_),
    .B(_1780_),
    .Y(_1781_)
);

NAND2X1 _11251_ (
    .A(_1776_),
    .B(_1781_),
    .Y(_1782_)
);

INVX1 _11252_ (
    .A(\datapath.alu.a [12]),
    .Y(_1783_)
);

INVX2 _11253_ (
    .A(\datapath.alu.a [13]),
    .Y(_1784_)
);

AOI22X1 _11254_ (
    .A(_1783_),
    .B(\datapath.alu.b [12]),
    .C(_1784_),
    .D(\datapath.alu.b [13]),
    .Y(_1785_)
);

INVX1 _11255_ (
    .A(\datapath.alu.b [13]),
    .Y(_1786_)
);

NAND2X1 _11256_ (
    .A(\datapath.alu.a [13]),
    .B(_1786_),
    .Y(_1787_)
);

INVX1 _11257_ (
    .A(\datapath.alu.b [12]),
    .Y(_1788_)
);

NAND2X1 _11258_ (
    .A(\datapath.alu.a [12]),
    .B(_1788_),
    .Y(_1789_)
);

NAND3X1 _11259_ (
    .A(_1787_),
    .B(_1789_),
    .C(_1785_),
    .Y(_1790_)
);

NOR2X1 _11260_ (
    .A(_1790_),
    .B(_1782_),
    .Y(_1791_)
);

NAND2X1 _11261_ (
    .A(\datapath.alu.a [11]),
    .B(\datapath.alu.b [11]),
    .Y(_1792_)
);

INVX2 _11262_ (
    .A(\datapath.alu.a [11]),
    .Y(_1793_)
);

INVX1 _11263_ (
    .A(\datapath.alu.b [11]),
    .Y(_1794_)
);

NAND2X1 _11264_ (
    .A(_1793_),
    .B(_1794_),
    .Y(_1795_)
);

NAND2X1 _11265_ (
    .A(_1792_),
    .B(_1795_),
    .Y(_1796_)
);

XNOR2X1 _11266_ (
    .A(\datapath.alu.a [10]),
    .B(\datapath.alu.b [10]),
    .Y(_1797_)
);

NAND2X1 _11267_ (
    .A(_1797_),
    .B(_1796_),
    .Y(_1798_)
);

INVX1 _11268_ (
    .A(\datapath.alu.a [9]),
    .Y(_1799_)
);

NAND2X1 _11269_ (
    .A(\datapath.alu.b [9]),
    .B(_1799_),
    .Y(_1800_)
);

INVX1 _11270_ (
    .A(\datapath.alu.b [9]),
    .Y(_1801_)
);

NAND2X1 _11271_ (
    .A(\datapath.alu.a [9]),
    .B(_1801_),
    .Y(_1802_)
);

AND2X2 _11272_ (
    .A(_1800_),
    .B(_1802_),
    .Y(_1803_)
);

INVX1 _11273_ (
    .A(\datapath.alu.b [8]),
    .Y(_1804_)
);

NOR2X1 _11274_ (
    .A(\datapath.alu.a [8]),
    .B(_1804_),
    .Y(_1805_)
);

INVX1 _11275_ (
    .A(\datapath.alu.a [8]),
    .Y(_1806_)
);

NOR2X1 _11276_ (
    .A(\datapath.alu.b [8]),
    .B(_1806_),
    .Y(_1807_)
);

NOR2X1 _11277_ (
    .A(_1805_),
    .B(_1807_),
    .Y(_1808_)
);

NAND2X1 _11278_ (
    .A(_1803_),
    .B(_1808_),
    .Y(_1809_)
);

NOR2X1 _11279_ (
    .A(_1798_),
    .B(_1809_),
    .Y(_1810_)
);

NAND2X1 _11280_ (
    .A(_1791_),
    .B(_1810_),
    .Y(_1811_)
);

NAND2X1 _11281_ (
    .A(\datapath.alu.a [7]),
    .B(\datapath.alu.b [7]),
    .Y(_1812_)
);

INVX2 _11282_ (
    .A(\datapath.alu.a [7]),
    .Y(_1813_)
);

INVX2 _11283_ (
    .A(\datapath.alu.b [7]),
    .Y(_1814_)
);

NAND2X1 _11284_ (
    .A(_1813_),
    .B(_1814_),
    .Y(_1815_)
);

NAND2X1 _11285_ (
    .A(_1812_),
    .B(_1815_),
    .Y(_1816_)
);

XNOR2X1 _11286_ (
    .A(\datapath.alu.a [6]),
    .B(\datapath.alu.b [6]),
    .Y(_1817_)
);

NAND2X1 _11287_ (
    .A(_1817_),
    .B(_1816_),
    .Y(_1818_)
);

INVX1 _11288_ (
    .A(\datapath.alu.a [4]),
    .Y(_1819_)
);

INVX2 _11289_ (
    .A(\datapath.alu.a [5]),
    .Y(_1820_)
);

AOI22X1 _11290_ (
    .A(_1819_),
    .B(\datapath.alu.b_4_bF$buf4 ),
    .C(_1820_),
    .D(\datapath.alu.b [5]),
    .Y(_1821_)
);

INVX2 _11291_ (
    .A(\datapath.alu.b [5]),
    .Y(_1822_)
);

NAND2X1 _11292_ (
    .A(\datapath.alu.a [5]),
    .B(_1822_),
    .Y(_1823_)
);

INVX8 _11293_ (
    .A(\datapath.alu.b_4_bF$buf3 ),
    .Y(_1824_)
);

NAND2X1 _11294_ (
    .A(\datapath.alu.a [4]),
    .B(_1824__bF$buf5),
    .Y(_1825_)
);

NAND3X1 _11295_ (
    .A(_1823_),
    .B(_1825_),
    .C(_1821_),
    .Y(_1826_)
);

NOR2X1 _11296_ (
    .A(_1826_),
    .B(_1818_),
    .Y(_1827_)
);

NAND2X1 _11297_ (
    .A(\datapath.alu.b_3_bF$buf7 ),
    .B(\datapath.alu.a [3]),
    .Y(_1828_)
);

OR2X2 _11298_ (
    .A(\datapath.alu.b_3_bF$buf6 ),
    .B(\datapath.alu.a [3]),
    .Y(_1829_)
);

NAND2X1 _11299_ (
    .A(_1828_),
    .B(_1829_),
    .Y(_1830_)
);

XNOR2X1 _11300_ (
    .A(\datapath.alu.b_2_bF$buf7 ),
    .B(\datapath.alu.a [2]),
    .Y(_1831_)
);

NAND2X1 _11301_ (
    .A(_1830_),
    .B(_1831_),
    .Y(_1832_)
);

INVX8 _11302_ (
    .A(\datapath.alu.b_1_bF$buf6 ),
    .Y(_1833_)
);

NAND2X1 _11303_ (
    .A(\datapath.alu.a [1]),
    .B(_1833__bF$buf7),
    .Y(_1834_)
);

INVX4 _11304_ (
    .A(\datapath.alu.b_0_bF$buf9 ),
    .Y(_1835_)
);

NAND2X1 _11305_ (
    .A(\datapath.alu.a [0]),
    .B(_1835_),
    .Y(_1836_)
);

NOR2X1 _11306_ (
    .A(\datapath.alu.a [1]),
    .B(_1833__bF$buf6),
    .Y(_1837_)
);

OAI21X1 _11307_ (
    .A(_1836_),
    .B(_1837_),
    .C(_1834_),
    .Y(_1838_)
);

INVX8 _11308_ (
    .A(\datapath.alu.b_2_bF$buf6 ),
    .Y(_1839_)
);

NOR2X1 _11309_ (
    .A(\datapath.alu.a [2]),
    .B(_1839__bF$buf6),
    .Y(_1840_)
);

INVX8 _11310_ (
    .A(\datapath.alu.b_3_bF$buf5 ),
    .Y(_1841_)
);

NOR2X1 _11311_ (
    .A(\datapath.alu.a [3]),
    .B(_1841__bF$buf7),
    .Y(_1842_)
);

NAND2X1 _11312_ (
    .A(\datapath.alu.a [3]),
    .B(_1841__bF$buf6),
    .Y(_1843_)
);

AOI21X1 _11313_ (
    .A(_1840_),
    .B(_1843_),
    .C(_1842_),
    .Y(_1844_)
);

OAI21X1 _11314_ (
    .A(_1838_),
    .B(_1832_),
    .C(_1844_),
    .Y(_1845_)
);

INVX1 _11315_ (
    .A(\datapath.alu.a [6]),
    .Y(_1846_)
);

NAND2X1 _11316_ (
    .A(\datapath.alu.b [6]),
    .B(_1846_),
    .Y(_1847_)
);

INVX1 _11317_ (
    .A(_1847_),
    .Y(_1848_)
);

NOR2X1 _11318_ (
    .A(\datapath.alu.b [7]),
    .B(_1813_),
    .Y(_1849_)
);

INVX1 _11319_ (
    .A(_1849_),
    .Y(_1850_)
);

NOR2X1 _11320_ (
    .A(\datapath.alu.a [7]),
    .B(_1814_),
    .Y(_1851_)
);

OAI21X1 _11321_ (
    .A(_1851_),
    .B(_1848_),
    .C(_1850_),
    .Y(_1852_)
);

NOR2X1 _11322_ (
    .A(\datapath.alu.a [5]),
    .B(_1822_),
    .Y(_1853_)
);

NOR2X1 _11323_ (
    .A(\datapath.alu.a [4]),
    .B(_1824__bF$buf4),
    .Y(_1854_)
);

OAI21X1 _11324_ (
    .A(_1853_),
    .B(_1854_),
    .C(_1823_),
    .Y(_1855_)
);

OAI21X1 _11325_ (
    .A(_1855_),
    .B(_1818_),
    .C(_1852_),
    .Y(_1856_)
);

AOI21X1 _11326_ (
    .A(_1845_),
    .B(_1827_),
    .C(_1856_),
    .Y(_1857_)
);

NOR2X1 _11327_ (
    .A(\datapath.alu.a [9]),
    .B(_1801_),
    .Y(_1858_)
);

OAI21X1 _11328_ (
    .A(_1858_),
    .B(_1805_),
    .C(_1802_),
    .Y(_1859_)
);

INVX2 _11329_ (
    .A(\datapath.alu.a [10]),
    .Y(_1860_)
);

NAND2X1 _11330_ (
    .A(\datapath.alu.b [10]),
    .B(_1860_),
    .Y(_1861_)
);

INVX1 _11331_ (
    .A(_1861_),
    .Y(_1862_)
);

NOR2X1 _11332_ (
    .A(\datapath.alu.a [11]),
    .B(_1794_),
    .Y(_1863_)
);

AOI21X1 _11333_ (
    .A(_1796_),
    .B(_1862_),
    .C(_1863_),
    .Y(_1864_)
);

OAI21X1 _11334_ (
    .A(_1859_),
    .B(_1798_),
    .C(_1864_),
    .Y(_1865_)
);

NAND2X1 _11335_ (
    .A(\datapath.alu.b [13]),
    .B(_1784_),
    .Y(_1866_)
);

INVX1 _11336_ (
    .A(_1866_),
    .Y(_1867_)
);

NAND2X1 _11337_ (
    .A(\datapath.alu.b [12]),
    .B(_1783_),
    .Y(_1868_)
);

INVX1 _11338_ (
    .A(_1868_),
    .Y(_1869_)
);

OAI21X1 _11339_ (
    .A(_1867_),
    .B(_1869_),
    .C(_1787_),
    .Y(_1870_)
);

OAI21X1 _11340_ (
    .A(\datapath.alu.a [15]),
    .B(_1774_),
    .C(_1778_),
    .Y(_1871_)
);

OAI21X1 _11341_ (
    .A(_1773_),
    .B(\datapath.alu.b [15]),
    .C(_1871_),
    .Y(_1872_)
);

OAI21X1 _11342_ (
    .A(_1870_),
    .B(_1782_),
    .C(_1872_),
    .Y(_1873_)
);

AOI21X1 _11343_ (
    .A(_1791_),
    .B(_1865_),
    .C(_1873_),
    .Y(_1874_)
);

OAI21X1 _11344_ (
    .A(_1857_),
    .B(_1811_),
    .C(_1874_),
    .Y(_1875_)
);

NAND2X1 _11345_ (
    .A(\datapath.alu.b [16]),
    .B(_1365_),
    .Y(_1876_)
);

OAI21X1 _11346_ (
    .A(\datapath.alu.a [17]),
    .B(_1333_),
    .C(_1876_),
    .Y(_1877_)
);

OAI21X1 _11347_ (
    .A(_1322_),
    .B(\datapath.alu.b [17]),
    .C(_1877_),
    .Y(_1878_)
);

NAND2X1 _11348_ (
    .A(\datapath.alu.a [19]),
    .B(_1215_),
    .Y(_1879_)
);

NOR2X1 _11349_ (
    .A(\datapath.alu.a [18]),
    .B(_1258_),
    .Y(_1880_)
);

NOR2X1 _11350_ (
    .A(\datapath.alu.a [19]),
    .B(_1215_),
    .Y(_1881_)
);

OAI21X1 _11351_ (
    .A(_1880_),
    .B(_1881_),
    .C(_1879_),
    .Y(_1882_)
);

OAI21X1 _11352_ (
    .A(_1300_),
    .B(_1878_),
    .C(_1882_),
    .Y(_1883_)
);

OAI22X1 _11353_ (
    .A(\datapath.alu.a [20]),
    .B(_1139_),
    .C(\datapath.alu.a [21]),
    .D(_1096_),
    .Y(_1884_)
);

OAI21X1 _11354_ (
    .A(_1086_),
    .B(\datapath.alu.b [21]),
    .C(_1884_),
    .Y(_1885_)
);

NAND2X1 _11355_ (
    .A(\datapath.alu.a [23]),
    .B(_978_),
    .Y(_1886_)
);

NOR2X1 _11356_ (
    .A(\datapath.alu.a [22]),
    .B(_1021_),
    .Y(_1887_)
);

NOR2X1 _11357_ (
    .A(\datapath.alu.a [23]),
    .B(_978_),
    .Y(_1888_)
);

OAI21X1 _11358_ (
    .A(_1887_),
    .B(_1888_),
    .C(_1886_),
    .Y(_1889_)
);

OAI21X1 _11359_ (
    .A(_1885_),
    .B(_1064_),
    .C(_1889_),
    .Y(_1890_)
);

AOI21X1 _11360_ (
    .A(_1883_),
    .B(_1193_),
    .C(_1890_),
    .Y(_1891_)
);

NOR2X1 _11361_ (
    .A(\datapath.alu.a [25]),
    .B(_1761_),
    .Y(_1892_)
);

NOR2X1 _11362_ (
    .A(\datapath.alu.a [24]),
    .B(_1766_),
    .Y(_1893_)
);

AOI21X1 _11363_ (
    .A(_1763_),
    .B(_1893_),
    .C(_1892_),
    .Y(_1894_)
);

NAND2X1 _11364_ (
    .A(\datapath.alu.a [27]),
    .B(_1654_),
    .Y(_1895_)
);

NOR2X1 _11365_ (
    .A(\datapath.alu.a [26]),
    .B(_1697_),
    .Y(_1896_)
);

NOR2X1 _11366_ (
    .A(\datapath.alu.a [27]),
    .B(_1654_),
    .Y(_1897_)
);

OAI21X1 _11367_ (
    .A(_1896_),
    .B(_1897_),
    .C(_1895_),
    .Y(_1898_)
);

OAI21X1 _11368_ (
    .A(_1740_),
    .B(_1894_),
    .C(_1898_),
    .Y(_1899_)
);

NOR2X1 _11369_ (
    .A(\datapath.alu.a [29]),
    .B(_1536_),
    .Y(_1900_)
);

NOR2X1 _11370_ (
    .A(\datapath.alu.a [28]),
    .B(_1579_),
    .Y(_1901_)
);

AOI21X1 _11371_ (
    .A(_1558_),
    .B(_1901_),
    .C(_1900_),
    .Y(_1902_)
);

NOR2X1 _11372_ (
    .A(\datapath.alu.a [31]),
    .B(_924_),
    .Y(_1903_)
);

NOR2X1 _11373_ (
    .A(\datapath.alu.a [30]),
    .B(_1461_),
    .Y(_1904_)
);

AOI21X1 _11374_ (
    .A(_946_),
    .B(_1904_),
    .C(_1903_),
    .Y(_1905_)
);

OAI21X1 _11375_ (
    .A(_1504_),
    .B(_1902_),
    .C(_1905_),
    .Y(_1906_)
);

AOI21X1 _11376_ (
    .A(_1899_),
    .B(_1633_),
    .C(_1906_),
    .Y(_1907_)
);

OAI21X1 _11377_ (
    .A(_1770_),
    .B(_1891_),
    .C(_1907_),
    .Y(_1908_)
);

AOI21X1 _11378_ (
    .A(_1875_),
    .B(_1771_),
    .C(_1908_),
    .Y(_1909_)
);

NAND2X1 _11379_ (
    .A(_946_),
    .B(_1909_),
    .Y(_1910_)
);

OR2X2 _11380_ (
    .A(_1440_),
    .B(_1770_),
    .Y(_1911_)
);

NAND2X1 _11381_ (
    .A(_1778_),
    .B(_1780_),
    .Y(_1912_)
);

AOI21X1 _11382_ (
    .A(_1772_),
    .B(_1775_),
    .C(_1912_),
    .Y(_1913_)
);

INVX1 _11383_ (
    .A(_1790_),
    .Y(_1914_)
);

NAND2X1 _11384_ (
    .A(_1913_),
    .B(_1914_),
    .Y(_1915_)
);

INVX2 _11385_ (
    .A(\datapath.alu.b [10]),
    .Y(_1916_)
);

NAND2X1 _11386_ (
    .A(\datapath.alu.a [10]),
    .B(_1916_),
    .Y(_1917_)
);

NAND2X1 _11387_ (
    .A(_1861_),
    .B(_1917_),
    .Y(_1918_)
);

AOI21X1 _11388_ (
    .A(_1792_),
    .B(_1795_),
    .C(_1918_),
    .Y(_1919_)
);

NAND2X1 _11389_ (
    .A(_1800_),
    .B(_1802_),
    .Y(_1920_)
);

NAND2X1 _11390_ (
    .A(\datapath.alu.b [8]),
    .B(_1806_),
    .Y(_1921_)
);

NAND2X1 _11391_ (
    .A(\datapath.alu.a [8]),
    .B(_1804_),
    .Y(_1922_)
);

NAND2X1 _11392_ (
    .A(_1921_),
    .B(_1922_),
    .Y(_1923_)
);

NOR2X1 _11393_ (
    .A(_1920_),
    .B(_1923_),
    .Y(_1924_)
);

NAND2X1 _11394_ (
    .A(_1919_),
    .B(_1924_),
    .Y(_1925_)
);

NOR2X1 _11395_ (
    .A(_1925_),
    .B(_1915_),
    .Y(_1926_)
);

XNOR2X1 _11396_ (
    .A(\datapath.alu.b_1_bF$buf5 ),
    .B(\datapath.alu.a [1]),
    .Y(_1927_)
);

NOR2X1 _11397_ (
    .A(\datapath.alu.b_0_bF$buf8 ),
    .B(\datapath.alu.a [0]),
    .Y(_1928_)
);

NAND2X1 _11398_ (
    .A(\datapath.alu.b_0_bF$buf7 ),
    .B(\datapath.alu.a [0]),
    .Y(_1929_)
);

INVX1 _11399_ (
    .A(_1929_),
    .Y(_1930_)
);

OAI21X1 _11400_ (
    .A(_1928_),
    .B(_1930_),
    .C(_1927_),
    .Y(_1931_)
);

NOR2X1 _11401_ (
    .A(_1832_),
    .B(_1931_),
    .Y(_1932_)
);

NAND3X1 _11402_ (
    .A(_1827_),
    .B(_1932_),
    .C(_1926_),
    .Y(_1933_)
);

NOR2X1 _11403_ (
    .A(_1933_),
    .B(_1911_),
    .Y(_1934_)
);

INVX1 _11404_ (
    .A(\datapath.alu.funsel [1]),
    .Y(_1935_)
);

NOR2X1 _11405_ (
    .A(\datapath.alu.funsel [0]),
    .B(_1935_),
    .Y(_1936_)
);

NOR2X1 _11406_ (
    .A(\datapath.alu.funsel [2]),
    .B(_1903_),
    .Y(_1937_)
);

NAND2X1 _11407_ (
    .A(_1936_),
    .B(_1937_),
    .Y(_1938_)
);

NOR2X1 _11408_ (
    .A(_1938_),
    .B(_1934_),
    .Y(_1939_)
);

NAND2X1 _11409_ (
    .A(\datapath.alu.funsel [0]),
    .B(\datapath.alu.funsel [1]),
    .Y(_1940_)
);

NOR2X1 _11410_ (
    .A(\datapath.alu.funsel [2]),
    .B(_1940_),
    .Y(_1941_)
);

OAI21X1 _11411_ (
    .A(_1933_),
    .B(_1911_),
    .C(_1941_),
    .Y(_1942_)
);

INVX1 _11412_ (
    .A(\datapath.alu.a [0]),
    .Y(_1943_)
);

NAND2X1 _11413_ (
    .A(\datapath.alu.b_0_bF$buf6 ),
    .B(\datapath.alu.a [1]),
    .Y(_1944_)
);

OAI21X1 _11414_ (
    .A(\datapath.alu.b_0_bF$buf5 ),
    .B(_1943_),
    .C(_1944_),
    .Y(_1945_)
);

MUX2X1 _11415_ (
    .A(\datapath.alu.a [3]),
    .B(\datapath.alu.a [2]),
    .S(\datapath.alu.b_0_bF$buf4 ),
    .Y(_1946_)
);

NAND2X1 _11416_ (
    .A(\datapath.alu.b_1_bF$buf4 ),
    .B(_1946_),
    .Y(_1947_)
);

OAI21X1 _11417_ (
    .A(\datapath.alu.b_1_bF$buf3 ),
    .B(_1945_),
    .C(_1947_),
    .Y(_1948_)
);

NAND2X1 _11418_ (
    .A(_1839__bF$buf5),
    .B(_1948_),
    .Y(_1949_)
);

MUX2X1 _11419_ (
    .A(\datapath.alu.a [7]),
    .B(\datapath.alu.a [6]),
    .S(\datapath.alu.b_0_bF$buf3 ),
    .Y(_1950_)
);

NAND2X1 _11420_ (
    .A(\datapath.alu.b_1_bF$buf2 ),
    .B(_1950_),
    .Y(_1951_)
);

MUX2X1 _11421_ (
    .A(\datapath.alu.a [5]),
    .B(\datapath.alu.a [4]),
    .S(\datapath.alu.b_0_bF$buf2 ),
    .Y(_1952_)
);

NAND2X1 _11422_ (
    .A(_1833__bF$buf5),
    .B(_1952_),
    .Y(_1953_)
);

NAND2X1 _11423_ (
    .A(_1951_),
    .B(_1953_),
    .Y(_1954_)
);

NAND2X1 _11424_ (
    .A(\datapath.alu.b_2_bF$buf5 ),
    .B(_1954_),
    .Y(_1955_)
);

NAND3X1 _11425_ (
    .A(_1841__bF$buf5),
    .B(_1955_),
    .C(_1949_),
    .Y(_1956_)
);

NAND2X1 _11426_ (
    .A(\datapath.alu.a [14]),
    .B(_1835_),
    .Y(_1957_)
);

NAND2X1 _11427_ (
    .A(\datapath.alu.b_0_bF$buf1 ),
    .B(\datapath.alu.a [15]),
    .Y(_1958_)
);

NAND3X1 _11428_ (
    .A(\datapath.alu.b_1_bF$buf1 ),
    .B(_1958_),
    .C(_1957_),
    .Y(_1959_)
);

NAND2X1 _11429_ (
    .A(\datapath.alu.a [12]),
    .B(_1835_),
    .Y(_1960_)
);

NAND2X1 _11430_ (
    .A(\datapath.alu.b_0_bF$buf0 ),
    .B(\datapath.alu.a [13]),
    .Y(_1961_)
);

NAND3X1 _11431_ (
    .A(_1833__bF$buf4),
    .B(_1961_),
    .C(_1960_),
    .Y(_1962_)
);

NAND2X1 _11432_ (
    .A(_1959_),
    .B(_1962_),
    .Y(_1963_)
);

MUX2X1 _11433_ (
    .A(\datapath.alu.a [11]),
    .B(\datapath.alu.a [10]),
    .S(\datapath.alu.b_0_bF$buf9 ),
    .Y(_1964_)
);

NAND2X1 _11434_ (
    .A(\datapath.alu.b_1_bF$buf0 ),
    .B(_1964_),
    .Y(_1965_)
);

MUX2X1 _11435_ (
    .A(\datapath.alu.a [9]),
    .B(\datapath.alu.a [8]),
    .S(\datapath.alu.b_0_bF$buf8 ),
    .Y(_1966_)
);

NAND2X1 _11436_ (
    .A(_1833__bF$buf3),
    .B(_1966_),
    .Y(_1967_)
);

NAND3X1 _11437_ (
    .A(_1839__bF$buf4),
    .B(_1965_),
    .C(_1967_),
    .Y(_1968_)
);

OAI21X1 _11438_ (
    .A(_1839__bF$buf3),
    .B(_1963_),
    .C(_1968_),
    .Y(_1969_)
);

NAND2X1 _11439_ (
    .A(\datapath.alu.b_3_bF$buf4 ),
    .B(_1969_),
    .Y(_1970_)
);

INVX1 _11440_ (
    .A(\datapath.alu.funsel [2]),
    .Y(_1971_)
);

NAND2X1 _11441_ (
    .A(\datapath.alu.funsel [0]),
    .B(_1935_),
    .Y(_1972_)
);

NOR2X1 _11442_ (
    .A(_1971_),
    .B(_1972_),
    .Y(_1973_)
);

INVX2 _11443_ (
    .A(_1973_),
    .Y(_1974_)
);

NOR2X1 _11444_ (
    .A(\datapath.alu.b_4_bF$buf2 ),
    .B(_1974_),
    .Y(_1975_)
);

INVX2 _11445_ (
    .A(_1975_),
    .Y(_1976_)
);

AOI21X1 _11446_ (
    .A(_1970_),
    .B(_1956_),
    .C(_1976_),
    .Y(_1977_)
);

NAND2X1 _11447_ (
    .A(\datapath.alu.a [26]),
    .B(_1835_),
    .Y(_1978_)
);

NAND2X1 _11448_ (
    .A(\datapath.alu.b_0_bF$buf7 ),
    .B(\datapath.alu.a [27]),
    .Y(_1979_)
);

NAND3X1 _11449_ (
    .A(\datapath.alu.b_1_bF$buf6 ),
    .B(_1979_),
    .C(_1978_),
    .Y(_1980_)
);

NAND2X1 _11450_ (
    .A(\datapath.alu.a [24]),
    .B(_1835_),
    .Y(_1981_)
);

NAND2X1 _11451_ (
    .A(\datapath.alu.b_0_bF$buf6 ),
    .B(\datapath.alu.a [25]),
    .Y(_1982_)
);

NAND3X1 _11452_ (
    .A(_1833__bF$buf2),
    .B(_1982_),
    .C(_1981_),
    .Y(_1983_)
);

NAND3X1 _11453_ (
    .A(_1839__bF$buf2),
    .B(_1980_),
    .C(_1983_),
    .Y(_1984_)
);

NAND2X1 _11454_ (
    .A(\datapath.alu.a [30]),
    .B(_1835_),
    .Y(_1985_)
);

NAND2X1 _11455_ (
    .A(\datapath.alu.b_0_bF$buf5 ),
    .B(\datapath.alu.a [31]),
    .Y(_1986_)
);

NAND3X1 _11456_ (
    .A(\datapath.alu.b_1_bF$buf5 ),
    .B(_1986_),
    .C(_1985_),
    .Y(_1987_)
);

NAND2X1 _11457_ (
    .A(\datapath.alu.a [28]),
    .B(_1835_),
    .Y(_1988_)
);

NAND2X1 _11458_ (
    .A(\datapath.alu.b_0_bF$buf4 ),
    .B(\datapath.alu.a [29]),
    .Y(_1989_)
);

NAND3X1 _11459_ (
    .A(_1833__bF$buf1),
    .B(_1989_),
    .C(_1988_),
    .Y(_1990_)
);

NAND3X1 _11460_ (
    .A(\datapath.alu.b_2_bF$buf4 ),
    .B(_1987_),
    .C(_1990_),
    .Y(_1991_)
);

NAND3X1 _11461_ (
    .A(\datapath.alu.b_3_bF$buf3 ),
    .B(_1991_),
    .C(_1984_),
    .Y(_1992_)
);

NAND2X1 _11462_ (
    .A(\datapath.alu.a [18]),
    .B(_1835_),
    .Y(_1993_)
);

NAND2X1 _11463_ (
    .A(\datapath.alu.b_0_bF$buf3 ),
    .B(\datapath.alu.a [19]),
    .Y(_1994_)
);

NAND3X1 _11464_ (
    .A(\datapath.alu.b_1_bF$buf4 ),
    .B(_1994_),
    .C(_1993_),
    .Y(_1995_)
);

NAND2X1 _11465_ (
    .A(\datapath.alu.a [16]),
    .B(_1835_),
    .Y(_1996_)
);

NAND2X1 _11466_ (
    .A(\datapath.alu.b_0_bF$buf2 ),
    .B(\datapath.alu.a [17]),
    .Y(_1997_)
);

NAND3X1 _11467_ (
    .A(_1833__bF$buf0),
    .B(_1997_),
    .C(_1996_),
    .Y(_1998_)
);

NAND3X1 _11468_ (
    .A(_1839__bF$buf1),
    .B(_1995_),
    .C(_1998_),
    .Y(_1999_)
);

NAND2X1 _11469_ (
    .A(\datapath.alu.a [22]),
    .B(_1835_),
    .Y(_2000_)
);

NAND2X1 _11470_ (
    .A(\datapath.alu.b_0_bF$buf1 ),
    .B(\datapath.alu.a [23]),
    .Y(_2001_)
);

NAND3X1 _11471_ (
    .A(\datapath.alu.b_1_bF$buf3 ),
    .B(_2001_),
    .C(_2000_),
    .Y(_2002_)
);

NAND2X1 _11472_ (
    .A(\datapath.alu.a [20]),
    .B(_1835_),
    .Y(_2003_)
);

NAND2X1 _11473_ (
    .A(\datapath.alu.b_0_bF$buf0 ),
    .B(\datapath.alu.a [21]),
    .Y(_2004_)
);

NAND3X1 _11474_ (
    .A(_1833__bF$buf7),
    .B(_2004_),
    .C(_2003_),
    .Y(_2005_)
);

NAND3X1 _11475_ (
    .A(\datapath.alu.b_2_bF$buf3 ),
    .B(_2002_),
    .C(_2005_),
    .Y(_2006_)
);

NAND3X1 _11476_ (
    .A(_1841__bF$buf4),
    .B(_1999_),
    .C(_2006_),
    .Y(_2007_)
);

NAND2X1 _11477_ (
    .A(_1992_),
    .B(_2007_),
    .Y(_2008_)
);

NOR2X1 _11478_ (
    .A(_1824__bF$buf3),
    .B(_1974_),
    .Y(_2009_)
);

INVX1 _11479_ (
    .A(_2009_),
    .Y(_2010_)
);

NOR2X1 _11480_ (
    .A(_2010_),
    .B(_2008_),
    .Y(_2011_)
);

INVX1 _11481_ (
    .A(_1940_),
    .Y(_2012_)
);

NOR2X1 _11482_ (
    .A(\datapath.alu.funsel [3]),
    .B(_1971_),
    .Y(_2013_)
);

NAND2X1 _11483_ (
    .A(_2012_),
    .B(_2013_),
    .Y(_2014_)
);

NAND2X1 _11484_ (
    .A(\datapath.alu.funsel [3]),
    .B(\datapath.alu.funsel [2]),
    .Y(_2015_)
);

NOR2X1 _11485_ (
    .A(_1940_),
    .B(_2015_),
    .Y(_2016_)
);

INVX8 _11486_ (
    .A(_2016__bF$buf3),
    .Y(_2017_)
);

NAND2X1 _11487_ (
    .A(\datapath.alu.b_0_bF$buf9 ),
    .B(_1943_),
    .Y(_2018_)
);

OAI22X1 _11488_ (
    .A(_1929_),
    .B(_2014__bF$buf3),
    .C(_2018_),
    .D(_2017_),
    .Y(_2019_)
);

INVX1 _11489_ (
    .A(\datapath.alu.funsel [0]),
    .Y(_2020_)
);

NAND2X1 _11490_ (
    .A(_2020_),
    .B(_1935_),
    .Y(_2021_)
);

NOR2X1 _11491_ (
    .A(_2015_),
    .B(_2021_),
    .Y(_2022_)
);

NAND2X1 _11492_ (
    .A(\datapath.alu.a [0]),
    .B(_2022_),
    .Y(_2023_)
);

NAND2X1 _11493_ (
    .A(\datapath.alu.funsel [1]),
    .B(_2020_),
    .Y(_2024_)
);

INVX1 _11494_ (
    .A(\datapath.alu.funsel [3]),
    .Y(_2025_)
);

NAND2X1 _11495_ (
    .A(\datapath.alu.funsel [2]),
    .B(_2025_),
    .Y(_2026_)
);

NOR2X1 _11496_ (
    .A(_2024_),
    .B(_2026_),
    .Y(_2027_)
);

OAI21X1 _11497_ (
    .A(\datapath.alu.b_0_bF$buf8 ),
    .B(\datapath.alu.a [0]),
    .C(_2027__bF$buf3),
    .Y(_2028_)
);

NOR2X1 _11498_ (
    .A(_2015_),
    .B(_2024_),
    .Y(_2029_)
);

NAND2X1 _11499_ (
    .A(\datapath.alu.b_0_bF$buf7 ),
    .B(_2029_),
    .Y(_2030_)
);

NAND3X1 _11500_ (
    .A(_2030_),
    .B(_2023_),
    .C(_2028_),
    .Y(_2031_)
);

NOR2X1 _11501_ (
    .A(_2019_),
    .B(_2031_),
    .Y(_2032_)
);

NOR2X1 _11502_ (
    .A(\datapath.alu.b_1_bF$buf2 ),
    .B(_1836_),
    .Y(_2033_)
);

NAND2X1 _11503_ (
    .A(_1839__bF$buf0),
    .B(_2033_),
    .Y(_2034_)
);

NOR2X1 _11504_ (
    .A(\datapath.alu.b_3_bF$buf2 ),
    .B(_2034_),
    .Y(_2035_)
);

NOR2X1 _11505_ (
    .A(\datapath.alu.funsel [1]),
    .B(\datapath.alu.funsel [2]),
    .Y(_2036_)
);

INVX2 _11506_ (
    .A(_2036_),
    .Y(_2037_)
);

NAND2X1 _11507_ (
    .A(\datapath.alu.funsel [0]),
    .B(_2025_),
    .Y(_2038_)
);

OR2X2 _11508_ (
    .A(_2037_),
    .B(_2038_),
    .Y(_2039_)
);

NOR2X1 _11509_ (
    .A(\datapath.alu.b_4_bF$buf1 ),
    .B(_2039_),
    .Y(_2040_)
);

NAND2X1 _11510_ (
    .A(_2040_),
    .B(_2035_),
    .Y(_2041_)
);

NOR2X1 _11511_ (
    .A(_1928_),
    .B(_1930_),
    .Y(_2042_)
);

NAND2X1 _11512_ (
    .A(\datapath.alu.funsel [3]),
    .B(_2020_),
    .Y(_2043_)
);

NAND2X1 _11513_ (
    .A(_2038_),
    .B(_2043_),
    .Y(_2044_)
);

NOR2X1 _11514_ (
    .A(_2037_),
    .B(_2044_),
    .Y(_2045_)
);

NOR2X1 _11515_ (
    .A(\datapath.alu.funsel [0]),
    .B(\datapath.alu.funsel [1]),
    .Y(_2046_)
);

NAND2X1 _11516_ (
    .A(_2046_),
    .B(_2013_),
    .Y(_2047_)
);

OAI21X1 _11517_ (
    .A(_2037_),
    .B(_2043_),
    .C(_2047__bF$buf3),
    .Y(_2048_)
);

OAI21X1 _11518_ (
    .A(_2045_),
    .B(_2048_),
    .C(_2042_),
    .Y(_2049_)
);

NAND3X1 _11519_ (
    .A(_2041_),
    .B(_2049_),
    .C(_2032_),
    .Y(_2050_)
);

NOR3X1 _11520_ (
    .A(_2050_),
    .B(_2011_),
    .C(_1977_),
    .Y(_2051_)
);

OAI21X1 _11521_ (
    .A(_1942_),
    .B(_1909_),
    .C(_2051_),
    .Y(_2052_)
);

AOI21X1 _11522_ (
    .A(_1910_),
    .B(_1939_),
    .C(_2052_),
    .Y(_2053_)
);

INVX1 _11523_ (
    .A(_2053_),
    .Y(\datapath.alu.condtrue )
);

NOR2X1 _11524_ (
    .A(_2015_),
    .B(_1972_),
    .Y(_2054_)
);

NAND2X1 _11525_ (
    .A(\datapath.alu.b_0_bF$buf6 ),
    .B(\datapath.alu.a [24]),
    .Y(_2055_)
);

OAI21X1 _11526_ (
    .A(\datapath.alu.b_0_bF$buf5 ),
    .B(_967_),
    .C(_2055_),
    .Y(_2056_)
);

NAND2X1 _11527_ (
    .A(\datapath.alu.b_0_bF$buf4 ),
    .B(\datapath.alu.a [22]),
    .Y(_2057_)
);

OAI21X1 _11528_ (
    .A(\datapath.alu.b_0_bF$buf3 ),
    .B(_1086_),
    .C(_2057_),
    .Y(_2058_)
);

MUX2X1 _11529_ (
    .A(_2058_),
    .B(_2056_),
    .S(_1833__bF$buf6),
    .Y(_2059_)
);

NAND2X1 _11530_ (
    .A(\datapath.alu.b_2_bF$buf2 ),
    .B(_2059_),
    .Y(_2060_)
);

NOR2X1 _11531_ (
    .A(\datapath.alu.b_0_bF$buf2 ),
    .B(\datapath.alu.a [19]),
    .Y(_2061_)
);

NOR2X1 _11532_ (
    .A(\datapath.alu.a [20]),
    .B(_1835_),
    .Y(_2062_)
);

OAI21X1 _11533_ (
    .A(_2061_),
    .B(_2062_),
    .C(\datapath.alu.b_1_bF$buf1 ),
    .Y(_2063_)
);

NOR2X1 _11534_ (
    .A(\datapath.alu.b_0_bF$buf1 ),
    .B(\datapath.alu.a [17]),
    .Y(_2064_)
);

NOR2X1 _11535_ (
    .A(\datapath.alu.a [18]),
    .B(_1835_),
    .Y(_2065_)
);

OAI21X1 _11536_ (
    .A(_2064_),
    .B(_2065_),
    .C(_1833__bF$buf5),
    .Y(_2066_)
);

AND2X2 _11537_ (
    .A(_2063_),
    .B(_2066_),
    .Y(_2067_)
);

OAI21X1 _11538_ (
    .A(\datapath.alu.b_2_bF$buf1 ),
    .B(_2067_),
    .C(_2060_),
    .Y(_2068_)
);

NOR2X1 _11539_ (
    .A(\datapath.alu.b_3_bF$buf1 ),
    .B(_2068_),
    .Y(_2069_)
);

NAND2X1 _11540_ (
    .A(\datapath.alu.b_0_bF$buf0 ),
    .B(\datapath.alu.a [28]),
    .Y(_2070_)
);

OAI21X1 _11541_ (
    .A(\datapath.alu.b_0_bF$buf9 ),
    .B(_1643_),
    .C(_2070_),
    .Y(_2071_)
);

NAND2X1 _11542_ (
    .A(\datapath.alu.b_0_bF$buf8 ),
    .B(\datapath.alu.a [26]),
    .Y(_2072_)
);

OAI21X1 _11543_ (
    .A(\datapath.alu.b_0_bF$buf7 ),
    .B(_1760_),
    .C(_2072_),
    .Y(_2073_)
);

MUX2X1 _11544_ (
    .A(_2073_),
    .B(_2071_),
    .S(_1833__bF$buf4),
    .Y(_2074_)
);

NOR2X1 _11545_ (
    .A(\datapath.alu.b_2_bF$buf0 ),
    .B(_2074_),
    .Y(_2075_)
);

NAND2X1 _11546_ (
    .A(\datapath.alu.b_0_bF$buf6 ),
    .B(\datapath.alu.a [30]),
    .Y(_2076_)
);

OAI21X1 _11547_ (
    .A(\datapath.alu.b_0_bF$buf5 ),
    .B(_1526_),
    .C(_2076_),
    .Y(_2077_)
);

NAND2X1 _11548_ (
    .A(_1833__bF$buf3),
    .B(_2077_),
    .Y(_2078_)
);

OAI21X1 _11549_ (
    .A(_1833__bF$buf2),
    .B(_913_),
    .C(_2078_),
    .Y(_2079_)
);

AOI21X1 _11550_ (
    .A(\datapath.alu.b_2_bF$buf7 ),
    .B(_2079_),
    .C(_2075_),
    .Y(_2080_)
);

NOR2X1 _11551_ (
    .A(_1841__bF$buf3),
    .B(_2080_),
    .Y(_2081_)
);

OAI21X1 _11552_ (
    .A(_2081_),
    .B(_2069_),
    .C(_2054_),
    .Y(_2082_)
);

NOR2X1 _11553_ (
    .A(_1972_),
    .B(_2026_),
    .Y(_2083_)
);

NOR2X1 _11554_ (
    .A(\datapath.alu.b_0_bF$buf4 ),
    .B(_913_),
    .Y(_2084_)
);

MUX2X1 _11555_ (
    .A(_2077_),
    .B(_2084_),
    .S(_1833__bF$buf1),
    .Y(_2085_)
);

MUX2X1 _11556_ (
    .A(_2074_),
    .B(_2085_),
    .S(_1839__bF$buf6),
    .Y(_2086_)
);

AND2X2 _11557_ (
    .A(_2086_),
    .B(\datapath.alu.b_3_bF$buf0 ),
    .Y(_2087_)
);

OAI21X1 _11558_ (
    .A(_2087_),
    .B(_2069_),
    .C(_2083_),
    .Y(_2088_)
);

AOI21X1 _11559_ (
    .A(_2088_),
    .B(_2082_),
    .C(_1824__bF$buf2),
    .Y(_2089_)
);

MUX2X1 _11560_ (
    .A(\datapath.alu.a [8]),
    .B(\datapath.alu.a [7]),
    .S(\datapath.alu.b_0_bF$buf3 ),
    .Y(_2090_)
);

MUX2X1 _11561_ (
    .A(\datapath.alu.a [6]),
    .B(\datapath.alu.a [5]),
    .S(\datapath.alu.b_0_bF$buf2 ),
    .Y(_2091_)
);

MUX2X1 _11562_ (
    .A(_2091_),
    .B(_2090_),
    .S(_1833__bF$buf0),
    .Y(_2092_)
);

MUX2X1 _11563_ (
    .A(\datapath.alu.a [2]),
    .B(\datapath.alu.a [1]),
    .S(\datapath.alu.b_0_bF$buf1 ),
    .Y(_2093_)
);

INVX1 _11564_ (
    .A(\datapath.alu.a [3]),
    .Y(_2094_)
);

NAND2X1 _11565_ (
    .A(\datapath.alu.b_0_bF$buf0 ),
    .B(\datapath.alu.a [4]),
    .Y(_2095_)
);

OAI21X1 _11566_ (
    .A(\datapath.alu.b_0_bF$buf9 ),
    .B(_2094_),
    .C(_2095_),
    .Y(_2096_)
);

OAI21X1 _11567_ (
    .A(_1833__bF$buf7),
    .B(_2096_),
    .C(_1839__bF$buf5),
    .Y(_2097_)
);

AOI21X1 _11568_ (
    .A(_1833__bF$buf6),
    .B(_2093_),
    .C(_2097_),
    .Y(_2098_)
);

AOI21X1 _11569_ (
    .A(\datapath.alu.b_2_bF$buf6 ),
    .B(_2092_),
    .C(_2098_),
    .Y(_2099_)
);

NOR2X1 _11570_ (
    .A(\datapath.alu.a [16]),
    .B(_1835_),
    .Y(_2100_)
);

NOR2X1 _11571_ (
    .A(\datapath.alu.b_0_bF$buf8 ),
    .B(\datapath.alu.a [15]),
    .Y(_2101_)
);

OAI21X1 _11572_ (
    .A(_2101_),
    .B(_2100_),
    .C(\datapath.alu.b_1_bF$buf0 ),
    .Y(_2102_)
);

NAND2X1 _11573_ (
    .A(\datapath.alu.b_0_bF$buf7 ),
    .B(\datapath.alu.a [14]),
    .Y(_2103_)
);

OAI21X1 _11574_ (
    .A(\datapath.alu.b_0_bF$buf6 ),
    .B(_1784_),
    .C(_2103_),
    .Y(_2104_)
);

OAI21X1 _11575_ (
    .A(\datapath.alu.b_1_bF$buf6 ),
    .B(_2104_),
    .C(_2102_),
    .Y(_2105_)
);

MUX2X1 _11576_ (
    .A(\datapath.alu.a [12]),
    .B(\datapath.alu.a [11]),
    .S(\datapath.alu.b_0_bF$buf5 ),
    .Y(_2106_)
);

MUX2X1 _11577_ (
    .A(\datapath.alu.a [10]),
    .B(\datapath.alu.a [9]),
    .S(\datapath.alu.b_0_bF$buf4 ),
    .Y(_2107_)
);

MUX2X1 _11578_ (
    .A(_2107_),
    .B(_2106_),
    .S(_1833__bF$buf5),
    .Y(_2108_)
);

NAND2X1 _11579_ (
    .A(_1839__bF$buf4),
    .B(_2108_),
    .Y(_2109_)
);

OAI21X1 _11580_ (
    .A(_1839__bF$buf3),
    .B(_2105_),
    .C(_2109_),
    .Y(_2110_)
);

NAND2X1 _11581_ (
    .A(\datapath.alu.b_3_bF$buf7 ),
    .B(_2110_),
    .Y(_2111_)
);

OAI21X1 _11582_ (
    .A(\datapath.alu.b_3_bF$buf6 ),
    .B(_2099_),
    .C(_2111_),
    .Y(_2112_)
);

NAND2X1 _11583_ (
    .A(_1975_),
    .B(_2112_),
    .Y(_2113_)
);

OAI21X1 _11584_ (
    .A(_1927_),
    .B(_1929_),
    .C(_2045_),
    .Y(_2114_)
);

AOI21X1 _11585_ (
    .A(_1927_),
    .B(_1929_),
    .C(_2114_),
    .Y(_2115_)
);

INVX1 _11586_ (
    .A(_2115_),
    .Y(_2116_)
);

INVX1 _11587_ (
    .A(_2015_),
    .Y(_2117_)
);

NAND2X1 _11588_ (
    .A(_2046_),
    .B(_2117_),
    .Y(_2118_)
);

OAI21X1 _11589_ (
    .A(_1833__bF$buf4),
    .B(_2014__bF$buf2),
    .C(_2118__bF$buf3),
    .Y(_2119_)
);

INVX2 _11590_ (
    .A(\datapath.alu.a [1]),
    .Y(_2120_)
);

NAND2X1 _11591_ (
    .A(_1833__bF$buf3),
    .B(_2120_),
    .Y(_2121_)
);

NAND2X1 _11592_ (
    .A(_1936_),
    .B(_2013_),
    .Y(_2122_)
);

NOR2X1 _11593_ (
    .A(_1833__bF$buf2),
    .B(_2120_),
    .Y(_2123_)
);

OAI21X1 _11594_ (
    .A(_2123_),
    .B(_2047__bF$buf2),
    .C(_2122_),
    .Y(_2124_)
);

AOI22X1 _11595_ (
    .A(_2124_),
    .B(_2121_),
    .C(\datapath.alu.a [1]),
    .D(_2119_),
    .Y(_2125_)
);

AND2X2 _11596_ (
    .A(_2116_),
    .B(_2125_),
    .Y(_2126_)
);

INVX2 _11597_ (
    .A(_2040_),
    .Y(_2127_)
);

OAI21X1 _11598_ (
    .A(\datapath.alu.b_0_bF$buf3 ),
    .B(_2120_),
    .C(_1929_),
    .Y(_2128_)
);

NAND2X1 _11599_ (
    .A(_1833__bF$buf1),
    .B(_2128_),
    .Y(_2129_)
);

NOR2X1 _11600_ (
    .A(\datapath.alu.b_2_bF$buf5 ),
    .B(_2129_),
    .Y(_2130_)
);

NAND2X1 _11601_ (
    .A(_1841__bF$buf2),
    .B(_2130_),
    .Y(_2131_)
);

NOR2X1 _11602_ (
    .A(_2131_),
    .B(_2127_),
    .Y(_2132_)
);

NOR2X1 _11603_ (
    .A(_2043_),
    .B(_2037_),
    .Y(_2133_)
);

INVX4 _11604_ (
    .A(_2133__bF$buf3),
    .Y(_2134_)
);

AOI21X1 _11605_ (
    .A(_1927_),
    .B(_2018_),
    .C(_2134_),
    .Y(_2135_)
);

OAI21X1 _11606_ (
    .A(_1927_),
    .B(_2018_),
    .C(_2135_),
    .Y(_2136_)
);

AOI21X1 _11607_ (
    .A(_2120_),
    .B(_2016__bF$buf2),
    .C(_2029_),
    .Y(_2137_)
);

OAI21X1 _11608_ (
    .A(_1833__bF$buf0),
    .B(_2137_),
    .C(_2136_),
    .Y(_2138_)
);

NOR2X1 _11609_ (
    .A(_2132_),
    .B(_2138_),
    .Y(_2139_)
);

NAND3X1 _11610_ (
    .A(_2126_),
    .B(_2139_),
    .C(_2113_),
    .Y(_2140_)
);

NOR2X1 _11611_ (
    .A(_2140_),
    .B(_2089_),
    .Y(_2141_)
);

INVX1 _11612_ (
    .A(_2141_),
    .Y(\datapath.alu.c [1])
);

INVX4 _11613_ (
    .A(_2083_),
    .Y(_2142_)
);

INVX4 _11614_ (
    .A(_2054_),
    .Y(_2143_)
);

OAI21X1 _11615_ (
    .A(\datapath.alu.b_0_bF$buf2 ),
    .B(_1765_),
    .C(_1982_),
    .Y(_2144_)
);

OAI21X1 _11616_ (
    .A(\datapath.alu.b_0_bF$buf1 ),
    .B(_1010_),
    .C(_2001_),
    .Y(_2145_)
);

MUX2X1 _11617_ (
    .A(_2145_),
    .B(_2144_),
    .S(_1833__bF$buf7),
    .Y(_2146_)
);

OAI21X1 _11618_ (
    .A(\datapath.alu.b_0_bF$buf0 ),
    .B(_1128_),
    .C(_2004_),
    .Y(_2147_)
);

OAI21X1 _11619_ (
    .A(\datapath.alu.b_0_bF$buf9 ),
    .B(_1247_),
    .C(_1994_),
    .Y(_2148_)
);

MUX2X1 _11620_ (
    .A(_2148_),
    .B(_2147_),
    .S(_1833__bF$buf6),
    .Y(_2149_)
);

MUX2X1 _11621_ (
    .A(_2149_),
    .B(_2146_),
    .S(_1839__bF$buf2),
    .Y(_2150_)
);

OAI21X1 _11622_ (
    .A(\datapath.alu.b_0_bF$buf8 ),
    .B(_1568_),
    .C(_1989_),
    .Y(_2151_)
);

OAI21X1 _11623_ (
    .A(\datapath.alu.b_0_bF$buf7 ),
    .B(_1686_),
    .C(_1979_),
    .Y(_2152_)
);

MUX2X1 _11624_ (
    .A(_2152_),
    .B(_2151_),
    .S(_1833__bF$buf5),
    .Y(_2153_)
);

OAI21X1 _11625_ (
    .A(\datapath.alu.b_0_bF$buf6 ),
    .B(_1450_),
    .C(_1986_),
    .Y(_2154_)
);

MUX2X1 _11626_ (
    .A(_2154_),
    .B(\datapath.alu.a [31]),
    .S(_1833__bF$buf4),
    .Y(_2155_)
);

MUX2X1 _11627_ (
    .A(_2153_),
    .B(_2155_),
    .S(_1839__bF$buf1),
    .Y(_2156_)
);

MUX2X1 _11628_ (
    .A(_2150_),
    .B(_2156_),
    .S(_1841__bF$buf1),
    .Y(_2157_)
);

NAND2X1 _11629_ (
    .A(_1833__bF$buf3),
    .B(_2154_),
    .Y(_2158_)
);

MUX2X1 _11630_ (
    .A(_2153_),
    .B(_2158_),
    .S(_1839__bF$buf0),
    .Y(_2159_)
);

MUX2X1 _11631_ (
    .A(_2150_),
    .B(_2159_),
    .S(_1841__bF$buf0),
    .Y(_2160_)
);

OAI22X1 _11632_ (
    .A(_2142_),
    .B(_2160_),
    .C(_2143_),
    .D(_2157_),
    .Y(_2161_)
);

NAND3X1 _11633_ (
    .A(\datapath.alu.b_1_bF$buf5 ),
    .B(_1961_),
    .C(_1960_),
    .Y(_2162_)
);

NAND2X1 _11634_ (
    .A(_1833__bF$buf2),
    .B(_1964_),
    .Y(_2163_)
);

NAND3X1 _11635_ (
    .A(_1839__bF$buf6),
    .B(_2162_),
    .C(_2163_),
    .Y(_2164_)
);

NAND3X1 _11636_ (
    .A(\datapath.alu.b_1_bF$buf4 ),
    .B(_1997_),
    .C(_1996_),
    .Y(_2165_)
);

NAND3X1 _11637_ (
    .A(_1833__bF$buf1),
    .B(_1958_),
    .C(_1957_),
    .Y(_2166_)
);

NAND3X1 _11638_ (
    .A(\datapath.alu.b_2_bF$buf4 ),
    .B(_2165_),
    .C(_2166_),
    .Y(_2167_)
);

NAND3X1 _11639_ (
    .A(\datapath.alu.b_3_bF$buf5 ),
    .B(_2164_),
    .C(_2167_),
    .Y(_2168_)
);

MUX2X1 _11640_ (
    .A(_1966_),
    .B(_1950_),
    .S(\datapath.alu.b_1_bF$buf3 ),
    .Y(_2169_)
);

NOR2X1 _11641_ (
    .A(_1839__bF$buf5),
    .B(_2169_),
    .Y(_2170_)
);

INVX1 _11642_ (
    .A(_1952_),
    .Y(_2171_)
);

OAI21X1 _11643_ (
    .A(\datapath.alu.b_1_bF$buf2 ),
    .B(_1946_),
    .C(_1839__bF$buf4),
    .Y(_2172_)
);

AOI21X1 _11644_ (
    .A(\datapath.alu.b_1_bF$buf1 ),
    .B(_2171_),
    .C(_2172_),
    .Y(_2173_)
);

OAI21X1 _11645_ (
    .A(_2173_),
    .B(_2170_),
    .C(_1841__bF$buf7),
    .Y(_2174_)
);

NAND3X1 _11646_ (
    .A(_1973_),
    .B(_2168_),
    .C(_2174_),
    .Y(_2175_)
);

OAI21X1 _11647_ (
    .A(\datapath.alu.b_0_bF$buf5 ),
    .B(_1943_),
    .C(\datapath.alu.b_1_bF$buf0 ),
    .Y(_2176_)
);

INVX1 _11648_ (
    .A(\datapath.alu.a [2]),
    .Y(_2177_)
);

OAI21X1 _11649_ (
    .A(\datapath.alu.b_0_bF$buf4 ),
    .B(_2177_),
    .C(_1944_),
    .Y(_2178_)
);

OAI21X1 _11650_ (
    .A(\datapath.alu.b_1_bF$buf6 ),
    .B(_2178_),
    .C(_2176_),
    .Y(_2179_)
);

NOR2X1 _11651_ (
    .A(\datapath.alu.b_2_bF$buf3 ),
    .B(_2179_),
    .Y(_2180_)
);

NOR2X1 _11652_ (
    .A(\datapath.alu.b_3_bF$buf4 ),
    .B(_2039_),
    .Y(_2181_)
);

AOI21X1 _11653_ (
    .A(_2181_),
    .B(_2180_),
    .C(_2009_),
    .Y(_2182_)
);

NAND2X1 _11654_ (
    .A(_2182_),
    .B(_2175_),
    .Y(_2183_)
);

OAI21X1 _11655_ (
    .A(_1824__bF$buf1),
    .B(_2161_),
    .C(_2183_),
    .Y(_2184_)
);

XOR2X1 _11656_ (
    .A(\datapath.alu.b_2_bF$buf2 ),
    .B(\datapath.alu.a [2]),
    .Y(_2185_)
);

NOR2X1 _11657_ (
    .A(\datapath.alu.b_1_bF$buf5 ),
    .B(_2120_),
    .Y(_2186_)
);

NAND2X1 _11658_ (
    .A(\datapath.alu.b_1_bF$buf4 ),
    .B(_2120_),
    .Y(_2187_)
);

AOI21X1 _11659_ (
    .A(_2187_),
    .B(_2018_),
    .C(_2186_),
    .Y(_2188_)
);

AOI21X1 _11660_ (
    .A(_2185_),
    .B(_2188_),
    .C(_2134_),
    .Y(_2189_)
);

OAI21X1 _11661_ (
    .A(_2185_),
    .B(_2188_),
    .C(_2189_),
    .Y(_2190_)
);

OAI21X1 _11662_ (
    .A(_2186_),
    .B(_1837_),
    .C(_1930_),
    .Y(_2191_)
);

INVX1 _11663_ (
    .A(_2123_),
    .Y(_2192_)
);

AOI21X1 _11664_ (
    .A(_2191_),
    .B(_2192_),
    .C(_1831_),
    .Y(_2193_)
);

OAI21X1 _11665_ (
    .A(_1929_),
    .B(_1927_),
    .C(_2192_),
    .Y(_2194_)
);

OAI21X1 _11666_ (
    .A(_2185_),
    .B(_2194_),
    .C(_2045_),
    .Y(_2195_)
);

NOR2X1 _11667_ (
    .A(_2193_),
    .B(_2195_),
    .Y(_2196_)
);

NOR2X1 _11668_ (
    .A(_1940_),
    .B(_2026_),
    .Y(_2197_)
);

NAND2X1 _11669_ (
    .A(\datapath.alu.b_2_bF$buf1 ),
    .B(\datapath.alu.a [2]),
    .Y(_2198_)
);

INVX1 _11670_ (
    .A(_2198_),
    .Y(_2199_)
);

AOI22X1 _11671_ (
    .A(_1840_),
    .B(_2016__bF$buf1),
    .C(_2199_),
    .D(_2197_),
    .Y(_2200_)
);

AOI22X1 _11672_ (
    .A(_2029_),
    .B(\datapath.alu.b_2_bF$buf0 ),
    .C(\datapath.alu.a [2]),
    .D(_2022_),
    .Y(_2201_)
);

OAI21X1 _11673_ (
    .A(_2199_),
    .B(_2047__bF$buf1),
    .C(_2122_),
    .Y(_2202_)
);

OAI21X1 _11674_ (
    .A(\datapath.alu.b_2_bF$buf7 ),
    .B(\datapath.alu.a [2]),
    .C(_2202_),
    .Y(_2203_)
);

NAND3X1 _11675_ (
    .A(_2200_),
    .B(_2201_),
    .C(_2203_),
    .Y(_2204_)
);

NOR2X1 _11676_ (
    .A(_2204_),
    .B(_2196_),
    .Y(_2205_)
);

AND2X2 _11677_ (
    .A(_2205_),
    .B(_2190_),
    .Y(_2206_)
);

NAND2X1 _11678_ (
    .A(_2206_),
    .B(_2184_),
    .Y(\datapath.alu.c [2])
);

NAND2X1 _11679_ (
    .A(\datapath.alu.b_0_bF$buf3 ),
    .B(\datapath.alu.a [6]),
    .Y(_2207_)
);

OAI21X1 _11680_ (
    .A(\datapath.alu.b_0_bF$buf2 ),
    .B(_1820_),
    .C(_2207_),
    .Y(_2208_)
);

MUX2X1 _11681_ (
    .A(_2208_),
    .B(_2096_),
    .S(\datapath.alu.b_1_bF$buf3 ),
    .Y(_2209_)
);

NOR2X1 _11682_ (
    .A(\datapath.alu.b_2_bF$buf6 ),
    .B(_2209_),
    .Y(_2210_)
);

NAND2X1 _11683_ (
    .A(\datapath.alu.b_0_bF$buf1 ),
    .B(\datapath.alu.a [8]),
    .Y(_2211_)
);

OAI21X1 _11684_ (
    .A(\datapath.alu.b_0_bF$buf0 ),
    .B(_1813_),
    .C(_2211_),
    .Y(_2212_)
);

NAND2X1 _11685_ (
    .A(\datapath.alu.b_0_bF$buf9 ),
    .B(\datapath.alu.a [10]),
    .Y(_2213_)
);

OAI21X1 _11686_ (
    .A(\datapath.alu.b_0_bF$buf8 ),
    .B(_1799_),
    .C(_2213_),
    .Y(_2214_)
);

MUX2X1 _11687_ (
    .A(_2214_),
    .B(_2212_),
    .S(\datapath.alu.b_1_bF$buf2 ),
    .Y(_2215_)
);

NOR2X1 _11688_ (
    .A(_1839__bF$buf3),
    .B(_2215_),
    .Y(_2216_)
);

OAI21X1 _11689_ (
    .A(_2210_),
    .B(_2216_),
    .C(_1841__bF$buf6),
    .Y(_2217_)
);

AOI21X1 _11690_ (
    .A(\datapath.alu.b_0_bF$buf7 ),
    .B(_1247_),
    .C(_2064_),
    .Y(_2218_)
);

NOR2X1 _11691_ (
    .A(_1833__bF$buf0),
    .B(_2218_),
    .Y(_2219_)
);

AOI21X1 _11692_ (
    .A(\datapath.alu.b_0_bF$buf6 ),
    .B(_1365_),
    .C(_2101_),
    .Y(_2220_)
);

NOR2X1 _11693_ (
    .A(\datapath.alu.b_1_bF$buf1 ),
    .B(_2220_),
    .Y(_2221_)
);

OAI21X1 _11694_ (
    .A(_2219_),
    .B(_2221_),
    .C(\datapath.alu.b_2_bF$buf5 ),
    .Y(_2222_)
);

NAND2X1 _11695_ (
    .A(_1833__bF$buf7),
    .B(_2106_),
    .Y(_2223_)
);

OAI21X1 _11696_ (
    .A(_1833__bF$buf6),
    .B(_2104_),
    .C(_2223_),
    .Y(_2224_)
);

NAND2X1 _11697_ (
    .A(_1839__bF$buf2),
    .B(_2224_),
    .Y(_2225_)
);

NAND3X1 _11698_ (
    .A(\datapath.alu.b_3_bF$buf3 ),
    .B(_2225_),
    .C(_2222_),
    .Y(_2226_)
);

AOI21X1 _11699_ (
    .A(_2226_),
    .B(_2217_),
    .C(\datapath.alu.b_4_bF$buf0 ),
    .Y(_2227_)
);

MUX2X1 _11700_ (
    .A(_2073_),
    .B(_2056_),
    .S(\datapath.alu.b_1_bF$buf0 ),
    .Y(_2228_)
);

NAND2X1 _11701_ (
    .A(\datapath.alu.b_2_bF$buf4 ),
    .B(_2228_),
    .Y(_2229_)
);

NOR2X1 _11702_ (
    .A(_1833__bF$buf5),
    .B(_2058_),
    .Y(_2230_)
);

AOI21X1 _11703_ (
    .A(\datapath.alu.b_0_bF$buf5 ),
    .B(_1128_),
    .C(_2061_),
    .Y(_2231_)
);

NOR2X1 _11704_ (
    .A(\datapath.alu.b_1_bF$buf6 ),
    .B(_2231_),
    .Y(_2232_)
);

OAI21X1 _11705_ (
    .A(_2230_),
    .B(_2232_),
    .C(_1839__bF$buf1),
    .Y(_2233_)
);

NAND3X1 _11706_ (
    .A(_1841__bF$buf5),
    .B(_2229_),
    .C(_2233_),
    .Y(_2234_)
);

MUX2X1 _11707_ (
    .A(_2077_),
    .B(_2071_),
    .S(\datapath.alu.b_1_bF$buf5 ),
    .Y(_2235_)
);

NOR2X1 _11708_ (
    .A(\datapath.alu.b_2_bF$buf3 ),
    .B(_2235_),
    .Y(_2236_)
);

NAND2X1 _11709_ (
    .A(\datapath.alu.b_2_bF$buf2 ),
    .B(\datapath.alu.a [31]),
    .Y(_2237_)
);

INVX1 _11710_ (
    .A(_2237_),
    .Y(_2238_)
);

OAI21X1 _11711_ (
    .A(_2238_),
    .B(_2236_),
    .C(\datapath.alu.b_3_bF$buf2 ),
    .Y(_2239_)
);

AOI21X1 _11712_ (
    .A(_2234_),
    .B(_2239_),
    .C(_1824__bF$buf0),
    .Y(_2240_)
);

OAI21X1 _11713_ (
    .A(_2240_),
    .B(_2227_),
    .C(_2054_),
    .Y(_2241_)
);

NAND2X1 _11714_ (
    .A(_1833__bF$buf4),
    .B(_2084_),
    .Y(_2242_)
);

NOR2X1 _11715_ (
    .A(_1839__bF$buf0),
    .B(_2242_),
    .Y(_2243_)
);

OAI21X1 _11716_ (
    .A(_2243_),
    .B(_2236_),
    .C(\datapath.alu.b_3_bF$buf1 ),
    .Y(_2244_)
);

AOI21X1 _11717_ (
    .A(_2234_),
    .B(_2244_),
    .C(_1824__bF$buf5),
    .Y(_2245_)
);

OAI21X1 _11718_ (
    .A(_2245_),
    .B(_2227_),
    .C(_2083_),
    .Y(_2246_)
);

NAND2X1 _11719_ (
    .A(\datapath.alu.a [2]),
    .B(_1839__bF$buf6),
    .Y(_2247_)
);

OAI21X1 _11720_ (
    .A(_1840_),
    .B(_2188_),
    .C(_2247_),
    .Y(_2248_)
);

OAI21X1 _11721_ (
    .A(_1830_),
    .B(_2248_),
    .C(_2133__bF$buf2),
    .Y(_2249_)
);

AOI21X1 _11722_ (
    .A(_1830_),
    .B(_2248_),
    .C(_2249_),
    .Y(_2250_)
);

OR2X2 _11723_ (
    .A(_2044_),
    .B(_2037_),
    .Y(_2251_)
);

OAI21X1 _11724_ (
    .A(_2199_),
    .B(_2193_),
    .C(_1830_),
    .Y(_2252_)
);

AND2X2 _11725_ (
    .A(\datapath.alu.b_3_bF$buf0 ),
    .B(\datapath.alu.a [3]),
    .Y(_2253_)
);

NOR2X1 _11726_ (
    .A(\datapath.alu.b_3_bF$buf7 ),
    .B(\datapath.alu.a [3]),
    .Y(_2254_)
);

NOR2X1 _11727_ (
    .A(_2254_),
    .B(_2253_),
    .Y(_2255_)
);

AOI21X1 _11728_ (
    .A(_1834_),
    .B(_2187_),
    .C(_1929_),
    .Y(_2256_)
);

OAI21X1 _11729_ (
    .A(_2123_),
    .B(_2256_),
    .C(_2185_),
    .Y(_2257_)
);

NAND3X1 _11730_ (
    .A(_2255_),
    .B(_2198_),
    .C(_2257_),
    .Y(_2258_)
);

AOI21X1 _11731_ (
    .A(_2252_),
    .B(_2258_),
    .C(_2251__bF$buf3),
    .Y(_2259_)
);

MUX2X1 _11732_ (
    .A(\datapath.alu.a [2]),
    .B(\datapath.alu.a [3]),
    .S(\datapath.alu.b_0_bF$buf4 ),
    .Y(_2260_)
);

NAND2X1 _11733_ (
    .A(_1833__bF$buf3),
    .B(_2260_),
    .Y(_2261_)
);

OAI21X1 _11734_ (
    .A(_1833__bF$buf2),
    .B(_2128_),
    .C(_2261_),
    .Y(_2262_)
);

NOR2X1 _11735_ (
    .A(\datapath.alu.b_2_bF$buf1 ),
    .B(_2262_),
    .Y(_2263_)
);

NAND3X1 _11736_ (
    .A(_1841__bF$buf4),
    .B(_2040_),
    .C(_2263_),
    .Y(_2264_)
);

INVX1 _11737_ (
    .A(_1842_),
    .Y(_2265_)
);

OAI22X1 _11738_ (
    .A(_2094_),
    .B(_2118__bF$buf2),
    .C(_2265_),
    .D(_2017_),
    .Y(_2266_)
);

NAND2X1 _11739_ (
    .A(_2117_),
    .B(_1936_),
    .Y(_2267_)
);

OAI22X1 _11740_ (
    .A(_1830_),
    .B(_2047__bF$buf0),
    .C(_1841__bF$buf3),
    .D(_2267__bF$buf3),
    .Y(_2268_)
);

OAI22X1 _11741_ (
    .A(_1828_),
    .B(_2014__bF$buf1),
    .C(_2254_),
    .D(_2122_),
    .Y(_2269_)
);

NOR3X1 _11742_ (
    .A(_2268_),
    .B(_2266_),
    .C(_2269_),
    .Y(_2270_)
);

NAND2X1 _11743_ (
    .A(_2270_),
    .B(_2264_),
    .Y(_2271_)
);

NOR3X1 _11744_ (
    .A(_2250_),
    .B(_2271_),
    .C(_2259_),
    .Y(_2272_)
);

NAND3X1 _11745_ (
    .A(_2241_),
    .B(_2246_),
    .C(_2272_),
    .Y(\datapath.alu.c [3])
);

MUX2X1 _11746_ (
    .A(_2144_),
    .B(_2152_),
    .S(_1833__bF$buf1),
    .Y(_2273_)
);

NAND2X1 _11747_ (
    .A(\datapath.alu.b_2_bF$buf0 ),
    .B(_2273_),
    .Y(_2274_)
);

NOR2X1 _11748_ (
    .A(_1833__bF$buf0),
    .B(_2145_),
    .Y(_2275_)
);

NOR2X1 _11749_ (
    .A(\datapath.alu.b_1_bF$buf4 ),
    .B(_2147_),
    .Y(_2276_)
);

OAI21X1 _11750_ (
    .A(_2275_),
    .B(_2276_),
    .C(_1839__bF$buf5),
    .Y(_2277_)
);

NAND3X1 _11751_ (
    .A(_1841__bF$buf2),
    .B(_2274_),
    .C(_2277_),
    .Y(_2278_)
);

NAND2X1 _11752_ (
    .A(_1833__bF$buf7),
    .B(_2151_),
    .Y(_2279_)
);

NAND2X1 _11753_ (
    .A(\datapath.alu.b_1_bF$buf3 ),
    .B(_2154_),
    .Y(_2280_)
);

AOI21X1 _11754_ (
    .A(_2279_),
    .B(_2280_),
    .C(\datapath.alu.b_2_bF$buf7 ),
    .Y(_2281_)
);

OAI21X1 _11755_ (
    .A(_2238_),
    .B(_2281_),
    .C(\datapath.alu.b_3_bF$buf6 ),
    .Y(_2282_)
);

AOI21X1 _11756_ (
    .A(_2278_),
    .B(_2282_),
    .C(_2143_),
    .Y(_2283_)
);

NAND2X1 _11757_ (
    .A(\datapath.alu.b_3_bF$buf5 ),
    .B(_2281_),
    .Y(_2284_)
);

AOI21X1 _11758_ (
    .A(_2278_),
    .B(_2284_),
    .C(_2142_),
    .Y(_2285_)
);

OAI21X1 _11759_ (
    .A(_2285_),
    .B(_2283_),
    .C(\datapath.alu.b_4_bF$buf4 ),
    .Y(_2286_)
);

NAND2X1 _11760_ (
    .A(\datapath.alu.b_4_bF$buf3 ),
    .B(_1819_),
    .Y(_2287_)
);

NAND2X1 _11761_ (
    .A(_2287_),
    .B(_1825_),
    .Y(_2288_)
);

NOR2X1 _11762_ (
    .A(\datapath.alu.b_2_bF$buf6 ),
    .B(_2177_),
    .Y(_2289_)
);

OAI21X1 _11763_ (
    .A(_1840_),
    .B(_2289_),
    .C(_2255_),
    .Y(_2290_)
);

AOI21X1 _11764_ (
    .A(_2191_),
    .B(_2192_),
    .C(_2290_),
    .Y(_2291_)
);

OAI21X1 _11765_ (
    .A(_2198_),
    .B(_2254_),
    .C(_1828_),
    .Y(_2292_)
);

OAI21X1 _11766_ (
    .A(_2292_),
    .B(_2291_),
    .C(_2288_),
    .Y(_2293_)
);

INVX1 _11767_ (
    .A(_2288_),
    .Y(_2294_)
);

NAND2X1 _11768_ (
    .A(\datapath.alu.b_2_bF$buf5 ),
    .B(_2177_),
    .Y(_2295_)
);

AOI21X1 _11769_ (
    .A(_2295_),
    .B(_2247_),
    .C(_1830_),
    .Y(_2296_)
);

AOI21X1 _11770_ (
    .A(_2194_),
    .B(_2296_),
    .C(_2292_),
    .Y(_2297_)
);

AOI21X1 _11771_ (
    .A(_2297_),
    .B(_2294_),
    .C(_2251__bF$buf2),
    .Y(_2298_)
);

NAND3X1 _11772_ (
    .A(_1839__bF$buf4),
    .B(_1951_),
    .C(_1953_),
    .Y(_2299_)
);

NAND3X1 _11773_ (
    .A(\datapath.alu.b_2_bF$buf4 ),
    .B(_1965_),
    .C(_1967_),
    .Y(_2300_)
);

NAND3X1 _11774_ (
    .A(_1841__bF$buf1),
    .B(_2299_),
    .C(_2300_),
    .Y(_2301_)
);

NAND3X1 _11775_ (
    .A(_1839__bF$buf3),
    .B(_1959_),
    .C(_1962_),
    .Y(_2302_)
);

NAND3X1 _11776_ (
    .A(\datapath.alu.b_2_bF$buf3 ),
    .B(_1995_),
    .C(_1998_),
    .Y(_2303_)
);

NAND3X1 _11777_ (
    .A(\datapath.alu.b_3_bF$buf4 ),
    .B(_2302_),
    .C(_2303_),
    .Y(_2304_)
);

NAND3X1 _11778_ (
    .A(_1975_),
    .B(_2304_),
    .C(_2301_),
    .Y(_2305_)
);

INVX1 _11779_ (
    .A(_2033_),
    .Y(_2306_)
);

NAND2X1 _11780_ (
    .A(\datapath.alu.a [2]),
    .B(_1835_),
    .Y(_2307_)
);

NAND3X1 _11781_ (
    .A(\datapath.alu.b_1_bF$buf2 ),
    .B(_1944_),
    .C(_2307_),
    .Y(_2308_)
);

MUX2X1 _11782_ (
    .A(\datapath.alu.a [3]),
    .B(\datapath.alu.a [4]),
    .S(\datapath.alu.b_0_bF$buf3 ),
    .Y(_2309_)
);

NAND2X1 _11783_ (
    .A(_1833__bF$buf6),
    .B(_2309_),
    .Y(_2310_)
);

NAND3X1 _11784_ (
    .A(_1839__bF$buf2),
    .B(_2308_),
    .C(_2310_),
    .Y(_2311_)
);

OAI21X1 _11785_ (
    .A(_1839__bF$buf1),
    .B(_2306_),
    .C(_2311_),
    .Y(_2312_)
);

NAND2X1 _11786_ (
    .A(_1841__bF$buf0),
    .B(_2312_),
    .Y(_2313_)
);

OAI21X1 _11787_ (
    .A(_2127_),
    .B(_2313_),
    .C(_2305_),
    .Y(_2314_)
);

AOI21X1 _11788_ (
    .A(_2293_),
    .B(_2298_),
    .C(_2314_),
    .Y(_2315_)
);

NOR2X1 _11789_ (
    .A(\datapath.alu.b_3_bF$buf3 ),
    .B(_2094_),
    .Y(_2316_)
);

AOI21X1 _11790_ (
    .A(_1830_),
    .B(_2289_),
    .C(_2316_),
    .Y(_2317_)
);

OAI21X1 _11791_ (
    .A(_1832_),
    .B(_2188_),
    .C(_2317_),
    .Y(_2318_)
);

NAND2X1 _11792_ (
    .A(_2294_),
    .B(_2318_),
    .Y(_2319_)
);

AOI21X1 _11793_ (
    .A(_1828_),
    .B(_1829_),
    .C(_2185_),
    .Y(_2320_)
);

NOR2X1 _11794_ (
    .A(\datapath.alu.a [0]),
    .B(_1835_),
    .Y(_2321_)
);

OAI21X1 _11795_ (
    .A(_1837_),
    .B(_2321_),
    .C(_1834_),
    .Y(_2322_)
);

OAI21X1 _11796_ (
    .A(_2247_),
    .B(_2255_),
    .C(_1843_),
    .Y(_2323_)
);

AOI21X1 _11797_ (
    .A(_2320_),
    .B(_2322_),
    .C(_2323_),
    .Y(_2324_)
);

AOI21X1 _11798_ (
    .A(_2324_),
    .B(_2288_),
    .C(_2134_),
    .Y(_2325_)
);

NAND2X1 _11799_ (
    .A(\datapath.alu.b_4_bF$buf2 ),
    .B(\datapath.alu.a [4]),
    .Y(_2326_)
);

INVX1 _11800_ (
    .A(_2326_),
    .Y(_2327_)
);

AOI22X1 _11801_ (
    .A(_1854_),
    .B(_2016__bF$buf0),
    .C(_2327_),
    .D(_2197_),
    .Y(_2328_)
);

OAI21X1 _11802_ (
    .A(_2327_),
    .B(_2047__bF$buf3),
    .C(_2122_),
    .Y(_2329_)
);

OAI21X1 _11803_ (
    .A(\datapath.alu.b_4_bF$buf1 ),
    .B(\datapath.alu.a [4]),
    .C(_2329_),
    .Y(_2330_)
);

AOI22X1 _11804_ (
    .A(_2029_),
    .B(\datapath.alu.b_4_bF$buf0 ),
    .C(\datapath.alu.a [4]),
    .D(_2022_),
    .Y(_2331_)
);

NAND3X1 _11805_ (
    .A(_2328_),
    .B(_2331_),
    .C(_2330_),
    .Y(_2332_)
);

AOI21X1 _11806_ (
    .A(_2325_),
    .B(_2319_),
    .C(_2332_),
    .Y(_2333_)
);

NAND3X1 _11807_ (
    .A(_2333_),
    .B(_2286_),
    .C(_2315_),
    .Y(\datapath.alu.c [4])
);

NAND2X1 _11808_ (
    .A(\datapath.alu.b [5]),
    .B(_1820_),
    .Y(_2334_)
);

NAND2X1 _11809_ (
    .A(_2334_),
    .B(_1823_),
    .Y(_2335_)
);

OAI21X1 _11810_ (
    .A(_2294_),
    .B(_2297_),
    .C(_2326_),
    .Y(_2336_)
);

AOI21X1 _11811_ (
    .A(_2336_),
    .B(_2335_),
    .C(_2251__bF$buf1),
    .Y(_2337_)
);

OAI21X1 _11812_ (
    .A(_2335_),
    .B(_2336_),
    .C(_2337_),
    .Y(_2338_)
);

OAI21X1 _11813_ (
    .A(_1854_),
    .B(_2324_),
    .C(_1825_),
    .Y(_2339_)
);

AND2X2 _11814_ (
    .A(_2339_),
    .B(_2335_),
    .Y(_2340_)
);

NOR2X1 _11815_ (
    .A(_2335_),
    .B(_2339_),
    .Y(_2341_)
);

OAI21X1 _11816_ (
    .A(_2341_),
    .B(_2340_),
    .C(_2133__bF$buf1),
    .Y(_2342_)
);

MUX2X1 _11817_ (
    .A(_2074_),
    .B(_2059_),
    .S(\datapath.alu.b_2_bF$buf2 ),
    .Y(_2343_)
);

OAI21X1 _11818_ (
    .A(\datapath.alu.b_2_bF$buf1 ),
    .B(\datapath.alu.b_1_bF$buf1 ),
    .C(\datapath.alu.a [31]),
    .Y(_2344_)
);

OAI21X1 _11819_ (
    .A(\datapath.alu.b_2_bF$buf0 ),
    .B(_2078_),
    .C(_2344_),
    .Y(_2345_)
);

MUX2X1 _11820_ (
    .A(_2343_),
    .B(_2345_),
    .S(_1841__bF$buf7),
    .Y(_2346_)
);

NOR2X1 _11821_ (
    .A(\datapath.alu.b_2_bF$buf7 ),
    .B(_2085_),
    .Y(_2347_)
);

MUX2X1 _11822_ (
    .A(_2343_),
    .B(_2347_),
    .S(_1841__bF$buf6),
    .Y(_2348_)
);

OAI22X1 _11823_ (
    .A(_2142_),
    .B(_2348_),
    .C(_2143_),
    .D(_2346_),
    .Y(_2349_)
);

OR2X2 _11824_ (
    .A(_2104_),
    .B(\datapath.alu.b_1_bF$buf0 ),
    .Y(_2350_)
);

NAND3X1 _11825_ (
    .A(_1839__bF$buf0),
    .B(_2102_),
    .C(_2350_),
    .Y(_2351_)
);

NAND3X1 _11826_ (
    .A(\datapath.alu.b_2_bF$buf6 ),
    .B(_2063_),
    .C(_2066_),
    .Y(_2352_)
);

NAND3X1 _11827_ (
    .A(\datapath.alu.b_3_bF$buf2 ),
    .B(_2352_),
    .C(_2351_),
    .Y(_2353_)
);

MUX2X1 _11828_ (
    .A(_2108_),
    .B(_2092_),
    .S(\datapath.alu.b_2_bF$buf5 ),
    .Y(_2354_)
);

NAND2X1 _11829_ (
    .A(_1841__bF$buf5),
    .B(_2354_),
    .Y(_2355_)
);

NAND3X1 _11830_ (
    .A(_1975_),
    .B(_2355_),
    .C(_2353_),
    .Y(_2356_)
);

NAND2X1 _11831_ (
    .A(_1820_),
    .B(_1822_),
    .Y(_2357_)
);

NOR2X1 _11832_ (
    .A(_1820_),
    .B(_1822_),
    .Y(_2358_)
);

OAI21X1 _11833_ (
    .A(_2358_),
    .B(_2047__bF$buf2),
    .C(_2122_),
    .Y(_2359_)
);

AOI22X1 _11834_ (
    .A(_1853_),
    .B(_2016__bF$buf3),
    .C(_2358_),
    .D(_2197_),
    .Y(_2360_)
);

AOI22X1 _11835_ (
    .A(_2029_),
    .B(\datapath.alu.b [5]),
    .C(\datapath.alu.a [5]),
    .D(_2022_),
    .Y(_2361_)
);

NAND2X1 _11836_ (
    .A(_2360_),
    .B(_2361_),
    .Y(_2362_)
);

AOI21X1 _11837_ (
    .A(_2357_),
    .B(_2359_),
    .C(_2362_),
    .Y(_2363_)
);

NAND2X1 _11838_ (
    .A(\datapath.alu.b_1_bF$buf6 ),
    .B(_2260_),
    .Y(_2364_)
);

OAI21X1 _11839_ (
    .A(\datapath.alu.b_0_bF$buf2 ),
    .B(_1820_),
    .C(_2095_),
    .Y(_2365_)
);

OAI21X1 _11840_ (
    .A(\datapath.alu.b_1_bF$buf5 ),
    .B(_2365_),
    .C(_2364_),
    .Y(_2366_)
);

MUX2X1 _11841_ (
    .A(_2366_),
    .B(_2129_),
    .S(_1839__bF$buf6),
    .Y(_2367_)
);

NAND3X1 _11842_ (
    .A(_1841__bF$buf4),
    .B(_2040_),
    .C(_2367_),
    .Y(_2368_)
);

NAND3X1 _11843_ (
    .A(_2363_),
    .B(_2368_),
    .C(_2356_),
    .Y(_2369_)
);

AOI21X1 _11844_ (
    .A(\datapath.alu.b_4_bF$buf4 ),
    .B(_2349_),
    .C(_2369_),
    .Y(_2370_)
);

NAND3X1 _11845_ (
    .A(_2338_),
    .B(_2342_),
    .C(_2370_),
    .Y(\datapath.alu.c [5])
);

INVX1 _11846_ (
    .A(\datapath.alu.b [6]),
    .Y(_2371_)
);

NAND2X1 _11847_ (
    .A(\datapath.alu.a [6]),
    .B(_2371_),
    .Y(_2372_)
);

NAND2X1 _11848_ (
    .A(_1847_),
    .B(_2372_),
    .Y(_2373_)
);

OAI21X1 _11849_ (
    .A(_1820_),
    .B(_1822_),
    .C(_2326_),
    .Y(_2374_)
);

AND2X2 _11850_ (
    .A(_2374_),
    .B(_2357_),
    .Y(_2375_)
);

INVX1 _11851_ (
    .A(_2375_),
    .Y(_2376_)
);

AOI22X1 _11852_ (
    .A(_2334_),
    .B(_1823_),
    .C(_2287_),
    .D(_1825_),
    .Y(_2377_)
);

INVX1 _11853_ (
    .A(_2377_),
    .Y(_2378_)
);

OAI21X1 _11854_ (
    .A(_2378_),
    .B(_2297_),
    .C(_2376_),
    .Y(_2379_)
);

OAI21X1 _11855_ (
    .A(_2373_),
    .B(_2379_),
    .C(_2045_),
    .Y(_2380_)
);

AOI21X1 _11856_ (
    .A(_2373_),
    .B(_2379_),
    .C(_2380_),
    .Y(_2381_)
);

OAI21X1 _11857_ (
    .A(_1825_),
    .B(_2335_),
    .C(_1823_),
    .Y(_2382_)
);

NAND3X1 _11858_ (
    .A(_1830_),
    .B(_1831_),
    .C(_2322_),
    .Y(_2383_)
);

AOI21X1 _11859_ (
    .A(_2383_),
    .B(_2317_),
    .C(_1826_),
    .Y(_2384_)
);

OAI21X1 _11860_ (
    .A(_2382_),
    .B(_2384_),
    .C(_1817_),
    .Y(_2385_)
);

OAI21X1 _11861_ (
    .A(\datapath.alu.b_4_bF$buf3 ),
    .B(_1819_),
    .C(_1823_),
    .Y(_2386_)
);

OAI21X1 _11862_ (
    .A(\datapath.alu.a [5]),
    .B(_1822_),
    .C(_2386_),
    .Y(_2387_)
);

NOR2X1 _11863_ (
    .A(_2335_),
    .B(_2288_),
    .Y(_2388_)
);

NOR2X1 _11864_ (
    .A(_2289_),
    .B(_2316_),
    .Y(_2389_)
);

OAI21X1 _11865_ (
    .A(_2185_),
    .B(_2188_),
    .C(_2389_),
    .Y(_2390_)
);

NAND3X1 _11866_ (
    .A(_2388_),
    .B(_2265_),
    .C(_2390_),
    .Y(_2391_)
);

NAND3X1 _11867_ (
    .A(_2373_),
    .B(_2387_),
    .C(_2391_),
    .Y(_2392_)
);

NAND3X1 _11868_ (
    .A(_2133__bF$buf0),
    .B(_2392_),
    .C(_2385_),
    .Y(_2393_)
);

NAND2X1 _11869_ (
    .A(\datapath.alu.b_2_bF$buf4 ),
    .B(_2153_),
    .Y(_2394_)
);

NAND2X1 _11870_ (
    .A(_1839__bF$buf5),
    .B(_2146_),
    .Y(_2395_)
);

NAND3X1 _11871_ (
    .A(_1841__bF$buf3),
    .B(_2394_),
    .C(_2395_),
    .Y(_2396_)
);

INVX1 _11872_ (
    .A(_2344_),
    .Y(_2397_)
);

NOR2X1 _11873_ (
    .A(\datapath.alu.b_2_bF$buf3 ),
    .B(_2158_),
    .Y(_2398_)
);

OAI21X1 _11874_ (
    .A(_2397_),
    .B(_2398_),
    .C(\datapath.alu.b_3_bF$buf1 ),
    .Y(_2399_)
);

AOI21X1 _11875_ (
    .A(_2396_),
    .B(_2399_),
    .C(_2143_),
    .Y(_2400_)
);

NAND2X1 _11876_ (
    .A(\datapath.alu.b_3_bF$buf0 ),
    .B(_2398_),
    .Y(_2401_)
);

AOI21X1 _11877_ (
    .A(_2396_),
    .B(_2401_),
    .C(_2142_),
    .Y(_2402_)
);

OAI21X1 _11878_ (
    .A(_2400_),
    .B(_2402_),
    .C(\datapath.alu.b_4_bF$buf2 ),
    .Y(_2403_)
);

AND2X2 _11879_ (
    .A(_2163_),
    .B(_2162_),
    .Y(_2404_)
);

MUX2X1 _11880_ (
    .A(_2404_),
    .B(_2169_),
    .S(\datapath.alu.b_2_bF$buf2 ),
    .Y(_2405_)
);

AND2X2 _11881_ (
    .A(_2165_),
    .B(_2166_),
    .Y(_2406_)
);

NAND2X1 _11882_ (
    .A(\datapath.alu.b_2_bF$buf1 ),
    .B(_2149_),
    .Y(_2407_)
);

OAI21X1 _11883_ (
    .A(\datapath.alu.b_2_bF$buf0 ),
    .B(_2406_),
    .C(_2407_),
    .Y(_2408_)
);

MUX2X1 _11884_ (
    .A(_2405_),
    .B(_2408_),
    .S(_1841__bF$buf2),
    .Y(_2409_)
);

NAND2X1 _11885_ (
    .A(\datapath.alu.b_2_bF$buf7 ),
    .B(_2179_),
    .Y(_2410_)
);

NAND2X1 _11886_ (
    .A(\datapath.alu.b_1_bF$buf4 ),
    .B(_2309_),
    .Y(_2411_)
);

MUX2X1 _11887_ (
    .A(\datapath.alu.a [5]),
    .B(\datapath.alu.a [6]),
    .S(\datapath.alu.b_0_bF$buf1 ),
    .Y(_2412_)
);

NAND2X1 _11888_ (
    .A(_1833__bF$buf5),
    .B(_2412_),
    .Y(_2413_)
);

NAND2X1 _11889_ (
    .A(_2411_),
    .B(_2413_),
    .Y(_2414_)
);

NAND2X1 _11890_ (
    .A(_1839__bF$buf4),
    .B(_2414_),
    .Y(_2415_)
);

NAND3X1 _11891_ (
    .A(_1841__bF$buf1),
    .B(_2410_),
    .C(_2415_),
    .Y(_2416_)
);

AOI22X1 _11892_ (
    .A(_2029_),
    .B(\datapath.alu.b [6]),
    .C(\datapath.alu.a [6]),
    .D(_2022_),
    .Y(_2417_)
);

NOR2X1 _11893_ (
    .A(_1846_),
    .B(_2371_),
    .Y(_2418_)
);

AOI22X1 _11894_ (
    .A(_1848_),
    .B(_2016__bF$buf2),
    .C(_2418_),
    .D(_2197_),
    .Y(_2419_)
);

NAND2X1 _11895_ (
    .A(_2419_),
    .B(_2417_),
    .Y(_2420_)
);

NAND2X1 _11896_ (
    .A(_1846_),
    .B(_2371_),
    .Y(_2421_)
);

OAI21X1 _11897_ (
    .A(_2418_),
    .B(_2047__bF$buf1),
    .C(_2122_),
    .Y(_2422_)
);

AOI21X1 _11898_ (
    .A(_2421_),
    .B(_2422_),
    .C(_2420_),
    .Y(_2423_)
);

OAI21X1 _11899_ (
    .A(_2127_),
    .B(_2416_),
    .C(_2423_),
    .Y(_2424_)
);

AOI21X1 _11900_ (
    .A(_1975_),
    .B(_2409_),
    .C(_2424_),
    .Y(_2425_)
);

NAND3X1 _11901_ (
    .A(_2393_),
    .B(_2403_),
    .C(_2425_),
    .Y(_2426_)
);

NOR2X1 _11902_ (
    .A(_2381_),
    .B(_2426_),
    .Y(_2427_)
);

INVX1 _11903_ (
    .A(_2427_),
    .Y(\datapath.alu.c [6])
);

AOI21X1 _11904_ (
    .A(_2379_),
    .B(_2373_),
    .C(_2418_),
    .Y(_2428_)
);

OR2X2 _11905_ (
    .A(_2428_),
    .B(_1816_),
    .Y(_2429_)
);

AOI21X1 _11906_ (
    .A(_2428_),
    .B(_1816_),
    .C(_2251__bF$buf0),
    .Y(_2430_)
);

INVX1 _11907_ (
    .A(_1816_),
    .Y(_2431_)
);

NAND3X1 _11908_ (
    .A(_2431_),
    .B(_2372_),
    .C(_2385_),
    .Y(_2432_)
);

INVX1 _11909_ (
    .A(_2372_),
    .Y(_2433_)
);

AOI21X1 _11910_ (
    .A(_2391_),
    .B(_2387_),
    .C(_2373_),
    .Y(_2434_)
);

OAI21X1 _11911_ (
    .A(_2433_),
    .B(_2434_),
    .C(_1816_),
    .Y(_2435_)
);

NAND3X1 _11912_ (
    .A(_2133__bF$buf3),
    .B(_2435_),
    .C(_2432_),
    .Y(_2436_)
);

MUX2X1 _11913_ (
    .A(_2235_),
    .B(_2228_),
    .S(\datapath.alu.b_2_bF$buf6 ),
    .Y(_2437_)
);

NOR2X1 _11914_ (
    .A(_1841__bF$buf0),
    .B(_913_),
    .Y(_2438_)
);

AOI21X1 _11915_ (
    .A(_2437_),
    .B(_1841__bF$buf7),
    .C(_2438_),
    .Y(_2439_)
);

NOR2X1 _11916_ (
    .A(\datapath.alu.b_2_bF$buf5 ),
    .B(_2242_),
    .Y(_2440_)
);

MUX2X1 _11917_ (
    .A(_2437_),
    .B(_2440_),
    .S(_1841__bF$buf6),
    .Y(_2441_)
);

OAI22X1 _11918_ (
    .A(_2143_),
    .B(_2439_),
    .C(_2142_),
    .D(_2441_),
    .Y(_2442_)
);

OAI21X1 _11919_ (
    .A(_2064_),
    .B(_2065_),
    .C(\datapath.alu.b_1_bF$buf3 ),
    .Y(_2443_)
);

OAI21X1 _11920_ (
    .A(_2101_),
    .B(_2100_),
    .C(_1833__bF$buf4),
    .Y(_2444_)
);

NAND3X1 _11921_ (
    .A(_1839__bF$buf3),
    .B(_2443_),
    .C(_2444_),
    .Y(_2445_)
);

OR2X2 _11922_ (
    .A(_2058_),
    .B(_1833__bF$buf3),
    .Y(_2446_)
);

OAI21X1 _11923_ (
    .A(_2061_),
    .B(_2062_),
    .C(_1833__bF$buf2),
    .Y(_2447_)
);

NAND3X1 _11924_ (
    .A(\datapath.alu.b_2_bF$buf4 ),
    .B(_2447_),
    .C(_2446_),
    .Y(_2448_)
);

NAND3X1 _11925_ (
    .A(\datapath.alu.b_3_bF$buf7 ),
    .B(_2445_),
    .C(_2448_),
    .Y(_2449_)
);

NOR2X1 _11926_ (
    .A(\datapath.alu.b_1_bF$buf2 ),
    .B(_2090_),
    .Y(_2450_)
);

NOR2X1 _11927_ (
    .A(_1833__bF$buf1),
    .B(_2107_),
    .Y(_2451_)
);

OAI21X1 _11928_ (
    .A(_2450_),
    .B(_2451_),
    .C(_1839__bF$buf2),
    .Y(_2452_)
);

OR2X2 _11929_ (
    .A(_2104_),
    .B(_1833__bF$buf0),
    .Y(_2453_)
);

NAND3X1 _11930_ (
    .A(\datapath.alu.b_2_bF$buf3 ),
    .B(_2223_),
    .C(_2453_),
    .Y(_2454_)
);

NAND3X1 _11931_ (
    .A(_1841__bF$buf5),
    .B(_2452_),
    .C(_2454_),
    .Y(_2455_)
);

NAND3X1 _11932_ (
    .A(_1975_),
    .B(_2449_),
    .C(_2455_),
    .Y(_2456_)
);

MUX2X1 _11933_ (
    .A(\datapath.alu.a [6]),
    .B(\datapath.alu.a [7]),
    .S(\datapath.alu.b_0_bF$buf0 ),
    .Y(_2457_)
);

NAND2X1 _11934_ (
    .A(_1833__bF$buf7),
    .B(_2457_),
    .Y(_2458_)
);

OAI21X1 _11935_ (
    .A(_1833__bF$buf6),
    .B(_2365_),
    .C(_2458_),
    .Y(_2459_)
);

MUX2X1 _11936_ (
    .A(_2459_),
    .B(_2262_),
    .S(_1839__bF$buf1),
    .Y(_2460_)
);

NAND3X1 _11937_ (
    .A(_1841__bF$buf4),
    .B(_2040_),
    .C(_2460_),
    .Y(_2461_)
);

INVX1 _11938_ (
    .A(_1851_),
    .Y(_2462_)
);

OAI22X1 _11939_ (
    .A(_1814_),
    .B(_2267__bF$buf2),
    .C(_2462_),
    .D(_2017_),
    .Y(_2463_)
);

OAI21X1 _11940_ (
    .A(\datapath.alu.a [7]),
    .B(\datapath.alu.b [7]),
    .C(_2027__bF$buf2),
    .Y(_2464_)
);

OAI21X1 _11941_ (
    .A(_1816_),
    .B(_2047__bF$buf0),
    .C(_2464_),
    .Y(_2465_)
);

OAI21X1 _11942_ (
    .A(_1814_),
    .B(_2014__bF$buf0),
    .C(_2118__bF$buf1),
    .Y(_2466_)
);

AND2X2 _11943_ (
    .A(_2466_),
    .B(\datapath.alu.a [7]),
    .Y(_2467_)
);

NOR3X1 _11944_ (
    .A(_2463_),
    .B(_2465_),
    .C(_2467_),
    .Y(_2468_)
);

NAND3X1 _11945_ (
    .A(_2461_),
    .B(_2456_),
    .C(_2468_),
    .Y(_2469_)
);

AOI21X1 _11946_ (
    .A(\datapath.alu.b_4_bF$buf1 ),
    .B(_2442_),
    .C(_2469_),
    .Y(_2470_)
);

NAND2X1 _11947_ (
    .A(_2470_),
    .B(_2436_),
    .Y(_2471_)
);

AOI21X1 _11948_ (
    .A(_2430_),
    .B(_2429_),
    .C(_2471_),
    .Y(_2472_)
);

INVX1 _11949_ (
    .A(_2472_),
    .Y(\datapath.alu.c [7])
);

OAI21X1 _11950_ (
    .A(_2256_),
    .B(_2123_),
    .C(_2296_),
    .Y(_2473_)
);

INVX1 _11951_ (
    .A(_2292_),
    .Y(_2474_)
);

NOR2X1 _11952_ (
    .A(_1817_),
    .B(_1816_),
    .Y(_2475_)
);

NAND2X1 _11953_ (
    .A(_2377_),
    .B(_2475_),
    .Y(_2476_)
);

AOI21X1 _11954_ (
    .A(_2473_),
    .B(_2474_),
    .C(_2476_),
    .Y(_2477_)
);

NAND2X1 _11955_ (
    .A(_2375_),
    .B(_2475_),
    .Y(_2478_)
);

OAI21X1 _11956_ (
    .A(\datapath.alu.a [7]),
    .B(\datapath.alu.b [7]),
    .C(_2418_),
    .Y(_2479_)
);

NAND3X1 _11957_ (
    .A(_1812_),
    .B(_2479_),
    .C(_2478_),
    .Y(_2480_)
);

OAI21X1 _11958_ (
    .A(_2480_),
    .B(_2477_),
    .C(_1923_),
    .Y(_2481_)
);

NAND2X1 _11959_ (
    .A(_2474_),
    .B(_2473_),
    .Y(_2482_)
);

AND2X2 _11960_ (
    .A(_2475_),
    .B(_2377_),
    .Y(_2483_)
);

AOI21X1 _11961_ (
    .A(_2482_),
    .B(_2483_),
    .C(_2480_),
    .Y(_2484_)
);

NAND2X1 _11962_ (
    .A(_1808_),
    .B(_2484_),
    .Y(_2485_)
);

NAND3X1 _11963_ (
    .A(_2045_),
    .B(_2481_),
    .C(_2485_),
    .Y(_2486_)
);

AOI21X1 _11964_ (
    .A(_1816_),
    .B(_2433_),
    .C(_1849_),
    .Y(_2487_)
);

OAI21X1 _11965_ (
    .A(_1818_),
    .B(_2387_),
    .C(_2487_),
    .Y(_2488_)
);

AOI21X1 _11966_ (
    .A(_2318_),
    .B(_1827_),
    .C(_2488_),
    .Y(_2489_)
);

AOI21X1 _11967_ (
    .A(_2489_),
    .B(_1923_),
    .C(_2134_),
    .Y(_2490_)
);

OAI21X1 _11968_ (
    .A(_1923_),
    .B(_2489_),
    .C(_2490_),
    .Y(_2491_)
);

OAI21X1 _11969_ (
    .A(\datapath.alu.b_2_bF$buf2 ),
    .B(_2273_),
    .C(_1991_),
    .Y(_2492_)
);

NAND2X1 _11970_ (
    .A(_1841__bF$buf3),
    .B(_2492_),
    .Y(_2493_)
);

NAND2X1 _11971_ (
    .A(_2438_),
    .B(_2054_),
    .Y(_2494_)
);

AOI21X1 _11972_ (
    .A(_2493_),
    .B(_2494_),
    .C(_1974_),
    .Y(_2495_)
);

NAND2X1 _11973_ (
    .A(\datapath.alu.b_1_bF$buf1 ),
    .B(_2412_),
    .Y(_2496_)
);

MUX2X1 _11974_ (
    .A(\datapath.alu.a [7]),
    .B(\datapath.alu.a [8]),
    .S(\datapath.alu.b_0_bF$buf9 ),
    .Y(_2497_)
);

NAND2X1 _11975_ (
    .A(_1833__bF$buf5),
    .B(_2497_),
    .Y(_2498_)
);

NAND3X1 _11976_ (
    .A(_1839__bF$buf0),
    .B(_2496_),
    .C(_2498_),
    .Y(_2499_)
);

NAND3X1 _11977_ (
    .A(\datapath.alu.b_2_bF$buf1 ),
    .B(_2308_),
    .C(_2310_),
    .Y(_2500_)
);

NAND3X1 _11978_ (
    .A(_1841__bF$buf2),
    .B(_2500_),
    .C(_2499_),
    .Y(_2501_)
);

OAI21X1 _11979_ (
    .A(\datapath.alu.b_2_bF$buf0 ),
    .B(_2306_),
    .C(\datapath.alu.b_3_bF$buf6 ),
    .Y(_2502_)
);

NAND3X1 _11980_ (
    .A(_2040_),
    .B(_2502_),
    .C(_2501_),
    .Y(_2503_)
);

NAND3X1 _11981_ (
    .A(\datapath.alu.b_2_bF$buf7 ),
    .B(_1959_),
    .C(_1962_),
    .Y(_2504_)
);

AOI21X1 _11982_ (
    .A(_1968_),
    .B(_2504_),
    .C(\datapath.alu.b_3_bF$buf5 ),
    .Y(_2505_)
);

AOI21X1 _11983_ (
    .A(_1999_),
    .B(_2006_),
    .C(_1841__bF$buf1),
    .Y(_2506_)
);

OAI21X1 _11984_ (
    .A(_2506_),
    .B(_2505_),
    .C(_1975_),
    .Y(_2507_)
);

NAND2X1 _11985_ (
    .A(\datapath.alu.a [8]),
    .B(\datapath.alu.b [8]),
    .Y(_2508_)
);

INVX1 _11986_ (
    .A(_2508_),
    .Y(_2509_)
);

AOI22X1 _11987_ (
    .A(_1805_),
    .B(_2016__bF$buf1),
    .C(_2509_),
    .D(_2197_),
    .Y(_2510_)
);

AOI22X1 _11988_ (
    .A(_2029_),
    .B(\datapath.alu.b [8]),
    .C(\datapath.alu.a [8]),
    .D(_2022_),
    .Y(_2511_)
);

NAND2X1 _11989_ (
    .A(_2510_),
    .B(_2511_),
    .Y(_2512_)
);

NAND2X1 _11990_ (
    .A(_1806_),
    .B(_1804_),
    .Y(_2513_)
);

OAI21X1 _11991_ (
    .A(_2509_),
    .B(_2047__bF$buf3),
    .C(_2122_),
    .Y(_2514_)
);

AOI21X1 _11992_ (
    .A(_2513_),
    .B(_2514_),
    .C(_2512_),
    .Y(_2515_)
);

NAND3X1 _11993_ (
    .A(_2503_),
    .B(_2515_),
    .C(_2507_),
    .Y(_2516_)
);

AOI21X1 _11994_ (
    .A(\datapath.alu.b_4_bF$buf0 ),
    .B(_2495_),
    .C(_2516_),
    .Y(_2517_)
);

NAND3X1 _11995_ (
    .A(_2491_),
    .B(_2486_),
    .C(_2517_),
    .Y(\datapath.alu.c [8])
);

OAI21X1 _11996_ (
    .A(_1813_),
    .B(_1814_),
    .C(_2479_),
    .Y(_2518_)
);

AOI21X1 _11997_ (
    .A(_2475_),
    .B(_2375_),
    .C(_2518_),
    .Y(_2519_)
);

OAI21X1 _11998_ (
    .A(_2476_),
    .B(_2297_),
    .C(_2519_),
    .Y(_2520_)
);

AOI21X1 _11999_ (
    .A(_2520_),
    .B(_1923_),
    .C(_2509_),
    .Y(_2521_)
);

AOI21X1 _12000_ (
    .A(_2521_),
    .B(_1803_),
    .C(_2251__bF$buf3),
    .Y(_2522_)
);

OAI21X1 _12001_ (
    .A(_1803_),
    .B(_2521_),
    .C(_2522_),
    .Y(_2523_)
);

OAI21X1 _12002_ (
    .A(_1805_),
    .B(_2489_),
    .C(_1922_),
    .Y(_2524_)
);

AOI21X1 _12003_ (
    .A(_1812_),
    .B(_1815_),
    .C(_2373_),
    .Y(_2525_)
);

NAND2X1 _12004_ (
    .A(_2525_),
    .B(_2388_),
    .Y(_2526_)
);

OAI21X1 _12005_ (
    .A(_2372_),
    .B(_1851_),
    .C(_1850_),
    .Y(_2527_)
);

AOI21X1 _12006_ (
    .A(_2382_),
    .B(_2525_),
    .C(_2527_),
    .Y(_2528_)
);

OAI21X1 _12007_ (
    .A(_2526_),
    .B(_2324_),
    .C(_2528_),
    .Y(_2529_)
);

NAND2X1 _12008_ (
    .A(_1924_),
    .B(_2529_),
    .Y(_2530_)
);

AOI21X1 _12009_ (
    .A(_1803_),
    .B(_1807_),
    .C(_2134_),
    .Y(_2531_)
);

AND2X2 _12010_ (
    .A(_2530_),
    .B(_2531_),
    .Y(_2532_)
);

OAI21X1 _12011_ (
    .A(_1803_),
    .B(_2524_),
    .C(_2532_),
    .Y(_2533_)
);

INVX1 _12012_ (
    .A(_2438_),
    .Y(_2534_)
);

OAI21X1 _12013_ (
    .A(\datapath.alu.b_3_bF$buf4 ),
    .B(_2080_),
    .C(_2534_),
    .Y(_2535_)
);

NOR2X1 _12014_ (
    .A(\datapath.alu.b_3_bF$buf3 ),
    .B(_2142_),
    .Y(_2536_)
);

AOI22X1 _12015_ (
    .A(_2086_),
    .B(_2536_),
    .C(_2054_),
    .D(_2535_),
    .Y(_2537_)
);

NOR2X1 _12016_ (
    .A(_1824__bF$buf4),
    .B(_2537_),
    .Y(_2538_)
);

AOI21X1 _12017_ (
    .A(_2068_),
    .B(\datapath.alu.b_3_bF$buf2 ),
    .C(_1976_),
    .Y(_2539_)
);

OAI21X1 _12018_ (
    .A(\datapath.alu.b_3_bF$buf1 ),
    .B(_2110_),
    .C(_2539_),
    .Y(_2540_)
);

OAI21X1 _12019_ (
    .A(\datapath.alu.b_2_bF$buf6 ),
    .B(_2129_),
    .C(\datapath.alu.b_3_bF$buf0 ),
    .Y(_2541_)
);

NAND2X1 _12020_ (
    .A(\datapath.alu.b_2_bF$buf5 ),
    .B(_2366_),
    .Y(_2542_)
);

INVX1 _12021_ (
    .A(_2457_),
    .Y(_2543_)
);

MUX2X1 _12022_ (
    .A(\datapath.alu.a [8]),
    .B(\datapath.alu.a [9]),
    .S(\datapath.alu.b_0_bF$buf8 ),
    .Y(_2544_)
);

NAND2X1 _12023_ (
    .A(_1833__bF$buf4),
    .B(_2544_),
    .Y(_2545_)
);

OAI21X1 _12024_ (
    .A(_1833__bF$buf3),
    .B(_2543_),
    .C(_2545_),
    .Y(_2546_)
);

NAND2X1 _12025_ (
    .A(_1839__bF$buf6),
    .B(_2546_),
    .Y(_2547_)
);

NAND2X1 _12026_ (
    .A(_2542_),
    .B(_2547_),
    .Y(_2548_)
);

NAND2X1 _12027_ (
    .A(_1841__bF$buf0),
    .B(_2548_),
    .Y(_2549_)
);

NAND3X1 _12028_ (
    .A(_2040_),
    .B(_2541_),
    .C(_2549_),
    .Y(_2550_)
);

OAI21X1 _12029_ (
    .A(\datapath.alu.a [9]),
    .B(_2017_),
    .C(_2267__bF$buf1),
    .Y(_2551_)
);

NOR2X1 _12030_ (
    .A(\datapath.alu.a [9]),
    .B(\datapath.alu.b [9]),
    .Y(_2552_)
);

NOR2X1 _12031_ (
    .A(_2026_),
    .B(_2021_),
    .Y(_2553_)
);

NAND2X1 _12032_ (
    .A(\datapath.alu.a [9]),
    .B(\datapath.alu.b [9]),
    .Y(_2554_)
);

AOI21X1 _12033_ (
    .A(_2553_),
    .B(_2554_),
    .C(_2027__bF$buf1),
    .Y(_2555_)
);

AOI21X1 _12034_ (
    .A(_2197_),
    .B(\datapath.alu.b [9]),
    .C(_2022_),
    .Y(_2556_)
);

OAI22X1 _12035_ (
    .A(_1799_),
    .B(_2556_),
    .C(_2552_),
    .D(_2555_),
    .Y(_2557_)
);

AOI21X1 _12036_ (
    .A(\datapath.alu.b [9]),
    .B(_2551_),
    .C(_2557_),
    .Y(_2558_)
);

NAND3X1 _12037_ (
    .A(_2558_),
    .B(_2550_),
    .C(_2540_),
    .Y(_2559_)
);

NOR2X1 _12038_ (
    .A(_2559_),
    .B(_2538_),
    .Y(_2560_)
);

NAND3X1 _12039_ (
    .A(_2523_),
    .B(_2533_),
    .C(_2560_),
    .Y(\datapath.alu.c [9])
);

OAI21X1 _12040_ (
    .A(_2508_),
    .B(_2552_),
    .C(_2554_),
    .Y(_2561_)
);

OAI21X1 _12041_ (
    .A(_1805_),
    .B(_1807_),
    .C(_1920_),
    .Y(_2562_)
);

INVX1 _12042_ (
    .A(_2562_),
    .Y(_2563_)
);

AOI21X1 _12043_ (
    .A(_2520_),
    .B(_2563_),
    .C(_2561_),
    .Y(_2564_)
);

OR2X2 _12044_ (
    .A(_2564_),
    .B(_1797_),
    .Y(_2565_)
);

AOI21X1 _12045_ (
    .A(_2564_),
    .B(_1797_),
    .C(_2251__bF$buf2),
    .Y(_2566_)
);

INVX1 _12046_ (
    .A(_1802_),
    .Y(_2567_)
);

AOI21X1 _12047_ (
    .A(_1807_),
    .B(_1800_),
    .C(_2567_),
    .Y(_873_)
);

AOI21X1 _12048_ (
    .A(_2530_),
    .B(_873_),
    .C(_1918_),
    .Y(_874_)
);

OAI21X1 _12049_ (
    .A(_1809_),
    .B(_2489_),
    .C(_873_),
    .Y(_875_)
);

OAI21X1 _12050_ (
    .A(_1797_),
    .B(_875_),
    .C(_2133__bF$buf2),
    .Y(_876_)
);

AOI21X1 _12051_ (
    .A(_2156_),
    .B(_1841__bF$buf7),
    .C(_2438_),
    .Y(_877_)
);

NAND2X1 _12052_ (
    .A(_2159_),
    .B(_2536_),
    .Y(_878_)
);

OAI21X1 _12053_ (
    .A(_2143_),
    .B(_877_),
    .C(_878_),
    .Y(_879_)
);

AOI21X1 _12054_ (
    .A(_2164_),
    .B(_2167_),
    .C(\datapath.alu.b_3_bF$buf7 ),
    .Y(_880_)
);

NAND3X1 _12055_ (
    .A(\datapath.alu.b_1_bF$buf0 ),
    .B(_2004_),
    .C(_2003_),
    .Y(_881_)
);

NAND3X1 _12056_ (
    .A(_1833__bF$buf2),
    .B(_1994_),
    .C(_1993_),
    .Y(_882_)
);

NAND3X1 _12057_ (
    .A(_1839__bF$buf5),
    .B(_881_),
    .C(_882_),
    .Y(_883_)
);

NAND3X1 _12058_ (
    .A(\datapath.alu.b_1_bF$buf6 ),
    .B(_1982_),
    .C(_1981_),
    .Y(_884_)
);

NAND3X1 _12059_ (
    .A(_1833__bF$buf1),
    .B(_2001_),
    .C(_2000_),
    .Y(_885_)
);

NAND3X1 _12060_ (
    .A(\datapath.alu.b_2_bF$buf4 ),
    .B(_884_),
    .C(_885_),
    .Y(_886_)
);

AOI21X1 _12061_ (
    .A(_883_),
    .B(_886_),
    .C(_1841__bF$buf6),
    .Y(_887_)
);

OAI21X1 _12062_ (
    .A(_880_),
    .B(_887_),
    .C(_1975_),
    .Y(_888_)
);

OAI21X1 _12063_ (
    .A(_1860_),
    .B(_1916_),
    .C(_2553_),
    .Y(_889_)
);

AOI22X1 _12064_ (
    .A(_1860_),
    .B(_1916_),
    .C(_2122_),
    .D(_889_),
    .Y(_890_)
);

NAND2X1 _12065_ (
    .A(\datapath.alu.a [10]),
    .B(\datapath.alu.b [10]),
    .Y(_891_)
);

OAI22X1 _12066_ (
    .A(_891_),
    .B(_2014__bF$buf3),
    .C(_1861_),
    .D(_2017_),
    .Y(_892_)
);

OAI22X1 _12067_ (
    .A(_1860_),
    .B(_2118__bF$buf0),
    .C(_1916_),
    .D(_2267__bF$buf0),
    .Y(_893_)
);

NOR3X1 _12068_ (
    .A(_892_),
    .B(_893_),
    .C(_890_),
    .Y(_894_)
);

NAND2X1 _12069_ (
    .A(\datapath.alu.b_1_bF$buf5 ),
    .B(_2497_),
    .Y(_895_)
);

MUX2X1 _12070_ (
    .A(\datapath.alu.a [9]),
    .B(\datapath.alu.a [10]),
    .S(\datapath.alu.b_0_bF$buf7 ),
    .Y(_896_)
);

NAND2X1 _12071_ (
    .A(_1833__bF$buf0),
    .B(_896_),
    .Y(_897_)
);

NAND3X1 _12072_ (
    .A(_1839__bF$buf4),
    .B(_895_),
    .C(_897_),
    .Y(_898_)
);

NAND3X1 _12073_ (
    .A(\datapath.alu.b_2_bF$buf3 ),
    .B(_2411_),
    .C(_2413_),
    .Y(_899_)
);

NAND3X1 _12074_ (
    .A(_1841__bF$buf5),
    .B(_898_),
    .C(_899_),
    .Y(_900_)
);

OAI21X1 _12075_ (
    .A(\datapath.alu.b_2_bF$buf2 ),
    .B(_2179_),
    .C(\datapath.alu.b_3_bF$buf6 ),
    .Y(_901_)
);

NAND3X1 _12076_ (
    .A(_2040_),
    .B(_901_),
    .C(_900_),
    .Y(_902_)
);

NAND3X1 _12077_ (
    .A(_902_),
    .B(_888_),
    .C(_894_),
    .Y(_904_)
);

AOI21X1 _12078_ (
    .A(\datapath.alu.b_4_bF$buf4 ),
    .B(_879_),
    .C(_904_),
    .Y(_905_)
);

OAI21X1 _12079_ (
    .A(_874_),
    .B(_876_),
    .C(_905_),
    .Y(_906_)
);

AOI21X1 _12080_ (
    .A(_2565_),
    .B(_2566_),
    .C(_906_),
    .Y(_907_)
);

INVX1 _12081_ (
    .A(_907_),
    .Y(\datapath.alu.c [10])
);

AND2X2 _12082_ (
    .A(_1795_),
    .B(_1792_),
    .Y(_908_)
);

OAI21X1 _12083_ (
    .A(_1797_),
    .B(_2564_),
    .C(_891_),
    .Y(_909_)
);

OR2X2 _12084_ (
    .A(_909_),
    .B(_908_),
    .Y(_910_)
);

AOI21X1 _12085_ (
    .A(_909_),
    .B(_908_),
    .C(_2251__bF$buf1),
    .Y(_911_)
);

INVX1 _12086_ (
    .A(_1917_),
    .Y(_912_)
);

AOI21X1 _12087_ (
    .A(_875_),
    .B(_1861_),
    .C(_912_),
    .Y(_914_)
);

AND2X2 _12088_ (
    .A(_914_),
    .B(_908_),
    .Y(_915_)
);

OAI21X1 _12089_ (
    .A(_908_),
    .B(_914_),
    .C(_2133__bF$buf1),
    .Y(_916_)
);

AND2X2 _12090_ (
    .A(_2222_),
    .B(_2225_),
    .Y(_917_)
);

NAND2X1 _12091_ (
    .A(_2229_),
    .B(_2233_),
    .Y(_918_)
);

AOI21X1 _12092_ (
    .A(_918_),
    .B(\datapath.alu.b_3_bF$buf5 ),
    .C(_1976_),
    .Y(_919_)
);

OAI21X1 _12093_ (
    .A(\datapath.alu.b_3_bF$buf4 ),
    .B(_917_),
    .C(_919_),
    .Y(_920_)
);

OAI21X1 _12094_ (
    .A(_1794_),
    .B(_2267__bF$buf3),
    .C(_920_),
    .Y(_921_)
);

OAI21X1 _12095_ (
    .A(\datapath.alu.b_2_bF$buf1 ),
    .B(_2235_),
    .C(_2237_),
    .Y(_922_)
);

AOI21X1 _12096_ (
    .A(_922_),
    .B(_1841__bF$buf4),
    .C(_2438_),
    .Y(_923_)
);

OAI21X1 _12097_ (
    .A(_2243_),
    .B(_2236_),
    .C(_2536_),
    .Y(_925_)
);

OAI21X1 _12098_ (
    .A(_2143_),
    .B(_923_),
    .C(_925_),
    .Y(_926_)
);

NAND2X1 _12099_ (
    .A(\datapath.alu.b_4_bF$buf3 ),
    .B(_926_),
    .Y(_927_)
);

NAND2X1 _12100_ (
    .A(\datapath.alu.b_2_bF$buf0 ),
    .B(_2459_),
    .Y(_928_)
);

NAND2X1 _12101_ (
    .A(\datapath.alu.b_1_bF$buf4 ),
    .B(_2544_),
    .Y(_929_)
);

OAI21X1 _12102_ (
    .A(\datapath.alu.b_0_bF$buf6 ),
    .B(_1793_),
    .C(_2213_),
    .Y(_930_)
);

OAI21X1 _12103_ (
    .A(\datapath.alu.b_1_bF$buf3 ),
    .B(_930_),
    .C(_929_),
    .Y(_931_)
);

NAND2X1 _12104_ (
    .A(_1839__bF$buf3),
    .B(_931_),
    .Y(_932_)
);

NAND2X1 _12105_ (
    .A(_928_),
    .B(_932_),
    .Y(_933_)
);

NAND2X1 _12106_ (
    .A(\datapath.alu.b_3_bF$buf3 ),
    .B(_2263_),
    .Y(_934_)
);

OAI21X1 _12107_ (
    .A(\datapath.alu.b_3_bF$buf2 ),
    .B(_933_),
    .C(_934_),
    .Y(_936_)
);

NAND2X1 _12108_ (
    .A(_2040_),
    .B(_936_),
    .Y(_937_)
);

INVX1 _12109_ (
    .A(_1792_),
    .Y(_938_)
);

OAI21X1 _12110_ (
    .A(_938_),
    .B(_2047__bF$buf2),
    .C(_2122_),
    .Y(_939_)
);

AOI22X1 _12111_ (
    .A(_1863_),
    .B(_2016__bF$buf0),
    .C(_938_),
    .D(_2197_),
    .Y(_940_)
);

OAI21X1 _12112_ (
    .A(_1793_),
    .B(_2118__bF$buf3),
    .C(_940_),
    .Y(_941_)
);

AOI21X1 _12113_ (
    .A(_1795_),
    .B(_939_),
    .C(_941_),
    .Y(_942_)
);

NAND3X1 _12114_ (
    .A(_937_),
    .B(_942_),
    .C(_927_),
    .Y(_943_)
);

NOR2X1 _12115_ (
    .A(_921_),
    .B(_943_),
    .Y(_944_)
);

OAI21X1 _12116_ (
    .A(_915_),
    .B(_916_),
    .C(_944_),
    .Y(_945_)
);

AOI21X1 _12117_ (
    .A(_911_),
    .B(_910_),
    .C(_945_),
    .Y(_947_)
);

INVX1 _12118_ (
    .A(_947_),
    .Y(\datapath.alu.c [11])
);

INVX2 _12119_ (
    .A(_1789_),
    .Y(_948_)
);

NOR2X1 _12120_ (
    .A(_1797_),
    .B(_1796_),
    .Y(_949_)
);

OAI21X1 _12121_ (
    .A(_891_),
    .B(_1796_),
    .C(_1792_),
    .Y(_950_)
);

AOI21X1 _12122_ (
    .A(_949_),
    .B(_2561_),
    .C(_950_),
    .Y(_951_)
);

INVX1 _12123_ (
    .A(_951_),
    .Y(_952_)
);

OAI21X1 _12124_ (
    .A(_1862_),
    .B(_912_),
    .C(_908_),
    .Y(_953_)
);

NOR2X1 _12125_ (
    .A(_2562_),
    .B(_953_),
    .Y(_954_)
);

AOI21X1 _12126_ (
    .A(_2520_),
    .B(_954_),
    .C(_952_),
    .Y(_955_)
);

INVX1 _12127_ (
    .A(_955_),
    .Y(_957_)
);

OAI21X1 _12128_ (
    .A(_1869_),
    .B(_948_),
    .C(_957_),
    .Y(_958_)
);

NAND2X1 _12129_ (
    .A(_1868_),
    .B(_1789_),
    .Y(_959_)
);

INVX1 _12130_ (
    .A(_959_),
    .Y(_960_)
);

AOI21X1 _12131_ (
    .A(_955_),
    .B(_960_),
    .C(_2251__bF$buf0),
    .Y(_961_)
);

OAI21X1 _12132_ (
    .A(_1922_),
    .B(_1858_),
    .C(_1802_),
    .Y(_962_)
);

NOR2X1 _12133_ (
    .A(\datapath.alu.b [11]),
    .B(_1793_),
    .Y(_963_)
);

INVX1 _12134_ (
    .A(_963_),
    .Y(_964_)
);

OAI21X1 _12135_ (
    .A(_1917_),
    .B(_1863_),
    .C(_964_),
    .Y(_965_)
);

AOI21X1 _12136_ (
    .A(_1919_),
    .B(_962_),
    .C(_965_),
    .Y(_966_)
);

OAI21X1 _12137_ (
    .A(_1925_),
    .B(_2489_),
    .C(_966_),
    .Y(_968_)
);

AND2X2 _12138_ (
    .A(_968_),
    .B(_960_),
    .Y(_969_)
);

OAI21X1 _12139_ (
    .A(_960_),
    .B(_968_),
    .C(_2133__bF$buf0),
    .Y(_970_)
);

AOI21X1 _12140_ (
    .A(_2302_),
    .B(_2303_),
    .C(\datapath.alu.b_3_bF$buf1 ),
    .Y(_971_)
);

NAND3X1 _12141_ (
    .A(_1839__bF$buf2),
    .B(_2002_),
    .C(_2005_),
    .Y(_972_)
);

NAND3X1 _12142_ (
    .A(\datapath.alu.b_2_bF$buf7 ),
    .B(_1980_),
    .C(_1983_),
    .Y(_973_)
);

AOI21X1 _12143_ (
    .A(_972_),
    .B(_973_),
    .C(_1841__bF$buf3),
    .Y(_974_)
);

OAI21X1 _12144_ (
    .A(_971_),
    .B(_974_),
    .C(_1973_),
    .Y(_975_)
);

INVX1 _12145_ (
    .A(_2039_),
    .Y(_976_)
);

NAND2X1 _12146_ (
    .A(\datapath.alu.b_1_bF$buf2 ),
    .B(_896_),
    .Y(_977_)
);

NAND2X1 _12147_ (
    .A(\datapath.alu.b_0_bF$buf5 ),
    .B(\datapath.alu.a [11]),
    .Y(_979_)
);

NAND3X1 _12148_ (
    .A(_1833__bF$buf7),
    .B(_979_),
    .C(_1960_),
    .Y(_980_)
);

NAND3X1 _12149_ (
    .A(_1839__bF$buf1),
    .B(_980_),
    .C(_977_),
    .Y(_981_)
);

NAND3X1 _12150_ (
    .A(\datapath.alu.b_2_bF$buf6 ),
    .B(_2496_),
    .C(_2498_),
    .Y(_982_)
);

NAND3X1 _12151_ (
    .A(_1841__bF$buf2),
    .B(_981_),
    .C(_982_),
    .Y(_983_)
);

NAND2X1 _12152_ (
    .A(\datapath.alu.b_2_bF$buf5 ),
    .B(_2033_),
    .Y(_984_)
);

NAND3X1 _12153_ (
    .A(\datapath.alu.b_3_bF$buf0 ),
    .B(_984_),
    .C(_2311_),
    .Y(_985_)
);

NAND3X1 _12154_ (
    .A(_976_),
    .B(_985_),
    .C(_983_),
    .Y(_986_)
);

NAND3X1 _12155_ (
    .A(_1824__bF$buf3),
    .B(_986_),
    .C(_975_),
    .Y(_987_)
);

NAND3X1 _12156_ (
    .A(_1839__bF$buf0),
    .B(_1987_),
    .C(_1990_),
    .Y(_988_)
);

AOI21X1 _12157_ (
    .A(_988_),
    .B(_2237_),
    .C(\datapath.alu.b_3_bF$buf7 ),
    .Y(_990_)
);

OAI21X1 _12158_ (
    .A(_2438_),
    .B(_990_),
    .C(_2054_),
    .Y(_991_)
);

NAND2X1 _12159_ (
    .A(_2281_),
    .B(_2536_),
    .Y(_992_)
);

NAND3X1 _12160_ (
    .A(\datapath.alu.b_4_bF$buf2 ),
    .B(_992_),
    .C(_991_),
    .Y(_993_)
);

NOR2X1 _12161_ (
    .A(_1783_),
    .B(_1788_),
    .Y(_994_)
);

AOI22X1 _12162_ (
    .A(_1869_),
    .B(_2016__bF$buf3),
    .C(_994_),
    .D(_2197_),
    .Y(_995_)
);

AOI22X1 _12163_ (
    .A(_2029_),
    .B(\datapath.alu.b [12]),
    .C(\datapath.alu.a [12]),
    .D(_2022_),
    .Y(_996_)
);

OAI21X1 _12164_ (
    .A(_994_),
    .B(_2047__bF$buf1),
    .C(_2122_),
    .Y(_997_)
);

OAI21X1 _12165_ (
    .A(\datapath.alu.a [12]),
    .B(\datapath.alu.b [12]),
    .C(_997_),
    .Y(_998_)
);

NAND3X1 _12166_ (
    .A(_995_),
    .B(_996_),
    .C(_998_),
    .Y(_999_)
);

AOI21X1 _12167_ (
    .A(_987_),
    .B(_993_),
    .C(_999_),
    .Y(_1001_)
);

OAI21X1 _12168_ (
    .A(_969_),
    .B(_970_),
    .C(_1001_),
    .Y(_1002_)
);

AOI21X1 _12169_ (
    .A(_958_),
    .B(_961_),
    .C(_1002_),
    .Y(_1003_)
);

INVX1 _12170_ (
    .A(_1003_),
    .Y(\datapath.alu.c [12])
);

NAND2X1 _12171_ (
    .A(_1866_),
    .B(_1787_),
    .Y(_1004_)
);

INVX2 _12172_ (
    .A(_1004_),
    .Y(_1005_)
);

AOI21X1 _12173_ (
    .A(_957_),
    .B(_959_),
    .C(_994_),
    .Y(_1006_)
);

OR2X2 _12174_ (
    .A(_1006_),
    .B(_1005_),
    .Y(_1007_)
);

AOI21X1 _12175_ (
    .A(_1006_),
    .B(_1005_),
    .C(_2251__bF$buf3),
    .Y(_1008_)
);

NOR3X1 _12176_ (
    .A(_948_),
    .B(_1005_),
    .C(_969_),
    .Y(_1009_)
);

OAI21X1 _12177_ (
    .A(_948_),
    .B(_969_),
    .C(_1005_),
    .Y(_1011_)
);

NAND2X1 _12178_ (
    .A(_2133__bF$buf3),
    .B(_1011_),
    .Y(_1012_)
);

AOI21X1 _12179_ (
    .A(_2345_),
    .B(_1841__bF$buf1),
    .C(_2438_),
    .Y(_1013_)
);

NAND2X1 _12180_ (
    .A(_2347_),
    .B(_2536_),
    .Y(_1014_)
);

OAI21X1 _12181_ (
    .A(_2143_),
    .B(_1013_),
    .C(_1014_),
    .Y(_1015_)
);

NAND3X1 _12182_ (
    .A(_1841__bF$buf0),
    .B(_2352_),
    .C(_2351_),
    .Y(_1016_)
);

NOR2X1 _12183_ (
    .A(_1841__bF$buf7),
    .B(_2343_),
    .Y(_1017_)
);

NOR2X1 _12184_ (
    .A(_1976_),
    .B(_1017_),
    .Y(_1018_)
);

NAND2X1 _12185_ (
    .A(\datapath.alu.a [13]),
    .B(\datapath.alu.b [13]),
    .Y(_1019_)
);

AOI22X1 _12186_ (
    .A(_1867_),
    .B(_2016__bF$buf2),
    .C(\datapath.alu.b [13]),
    .D(_2029_),
    .Y(_1020_)
);

NOR2X1 _12187_ (
    .A(\datapath.alu.a [13]),
    .B(\datapath.alu.b [13]),
    .Y(_1022_)
);

AOI21X1 _12188_ (
    .A(_2553_),
    .B(_1019_),
    .C(_2027__bF$buf0),
    .Y(_1023_)
);

OAI21X1 _12189_ (
    .A(_1022_),
    .B(_1023_),
    .C(_1020_),
    .Y(_1024_)
);

AOI21X1 _12190_ (
    .A(\datapath.alu.a [13]),
    .B(_2022_),
    .C(_1024_),
    .Y(_1025_)
);

OAI21X1 _12191_ (
    .A(_2014__bF$buf2),
    .B(_1019_),
    .C(_1025_),
    .Y(_1026_)
);

AOI21X1 _12192_ (
    .A(_1016_),
    .B(_1018_),
    .C(_1026_),
    .Y(_1027_)
);

NAND2X1 _12193_ (
    .A(\datapath.alu.b_2_bF$buf4 ),
    .B(_2546_),
    .Y(_1028_)
);

NAND2X1 _12194_ (
    .A(\datapath.alu.b_0_bF$buf4 ),
    .B(\datapath.alu.a [12]),
    .Y(_1029_)
);

OAI21X1 _12195_ (
    .A(\datapath.alu.b_0_bF$buf3 ),
    .B(_1784_),
    .C(_1029_),
    .Y(_1030_)
);

INVX1 _12196_ (
    .A(_1030_),
    .Y(_1031_)
);

NAND2X1 _12197_ (
    .A(\datapath.alu.b_1_bF$buf1 ),
    .B(_930_),
    .Y(_1033_)
);

OAI21X1 _12198_ (
    .A(\datapath.alu.b_1_bF$buf0 ),
    .B(_1031_),
    .C(_1033_),
    .Y(_1034_)
);

OAI21X1 _12199_ (
    .A(\datapath.alu.b_2_bF$buf3 ),
    .B(_1034_),
    .C(_1028_),
    .Y(_1035_)
);

NAND2X1 _12200_ (
    .A(_1841__bF$buf6),
    .B(_1035_),
    .Y(_1036_)
);

OAI21X1 _12201_ (
    .A(_1841__bF$buf5),
    .B(_2367_),
    .C(_1036_),
    .Y(_1037_)
);

OAI21X1 _12202_ (
    .A(_2127_),
    .B(_1037_),
    .C(_1027_),
    .Y(_1038_)
);

AOI21X1 _12203_ (
    .A(\datapath.alu.b_4_bF$buf1 ),
    .B(_1015_),
    .C(_1038_),
    .Y(_1039_)
);

OAI21X1 _12204_ (
    .A(_1009_),
    .B(_1012_),
    .C(_1039_),
    .Y(_1040_)
);

AOI21X1 _12205_ (
    .A(_1007_),
    .B(_1008_),
    .C(_1040_),
    .Y(_1041_)
);

INVX1 _12206_ (
    .A(_1041_),
    .Y(\datapath.alu.c [13])
);

AND2X2 _12207_ (
    .A(_1004_),
    .B(_959_),
    .Y(_1043_)
);

INVX1 _12208_ (
    .A(_1043_),
    .Y(_1044_)
);

INVX1 _12209_ (
    .A(_994_),
    .Y(_1045_)
);

OAI21X1 _12210_ (
    .A(_1022_),
    .B(_1045_),
    .C(_1019_),
    .Y(_1046_)
);

INVX1 _12211_ (
    .A(_1046_),
    .Y(_1047_)
);

OAI21X1 _12212_ (
    .A(_1044_),
    .B(_955_),
    .C(_1047_),
    .Y(_1048_)
);

NAND2X1 _12213_ (
    .A(_1912_),
    .B(_1048_),
    .Y(_1049_)
);

INVX1 _12214_ (
    .A(_1048_),
    .Y(_1050_)
);

AOI21X1 _12215_ (
    .A(_1050_),
    .B(_1781_),
    .C(_2251__bF$buf2),
    .Y(_1051_)
);

OAI21X1 _12216_ (
    .A(_1789_),
    .B(_1004_),
    .C(_1787_),
    .Y(_1052_)
);

AOI21X1 _12217_ (
    .A(_968_),
    .B(_1914_),
    .C(_1052_),
    .Y(_1054_)
);

AND2X2 _12218_ (
    .A(_1054_),
    .B(_1912_),
    .Y(_1055_)
);

OAI21X1 _12219_ (
    .A(_1912_),
    .B(_1054_),
    .C(_2133__bF$buf2),
    .Y(_1056_)
);

NAND2X1 _12220_ (
    .A(_2410_),
    .B(_2415_),
    .Y(_1057_)
);

AND2X2 _12221_ (
    .A(_895_),
    .B(_897_),
    .Y(_1058_)
);

AND2X2 _12222_ (
    .A(_1960_),
    .B(_979_),
    .Y(_1059_)
);

OAI21X1 _12223_ (
    .A(\datapath.alu.b_0_bF$buf2 ),
    .B(_1777_),
    .C(_1961_),
    .Y(_1060_)
);

NAND2X1 _12224_ (
    .A(_1833__bF$buf6),
    .B(_1060_),
    .Y(_1061_)
);

OAI21X1 _12225_ (
    .A(_1833__bF$buf5),
    .B(_1059_),
    .C(_1061_),
    .Y(_1062_)
);

MUX2X1 _12226_ (
    .A(_1062_),
    .B(_1058_),
    .S(_1839__bF$buf6),
    .Y(_1063_)
);

MUX2X1 _12227_ (
    .A(_1057_),
    .B(_1063_),
    .S(\datapath.alu.b_3_bF$buf6 ),
    .Y(_1065_)
);

NAND2X1 _12228_ (
    .A(_976_),
    .B(_1065_),
    .Y(_1066_)
);

NOR2X1 _12229_ (
    .A(\datapath.alu.b_3_bF$buf5 ),
    .B(_2408_),
    .Y(_1067_)
);

NAND2X1 _12230_ (
    .A(_2394_),
    .B(_2395_),
    .Y(_1068_)
);

NOR2X1 _12231_ (
    .A(_1841__bF$buf4),
    .B(_1068_),
    .Y(_1069_)
);

OAI21X1 _12232_ (
    .A(_1069_),
    .B(_1067_),
    .C(_1973_),
    .Y(_1070_)
);

AOI21X1 _12233_ (
    .A(_1066_),
    .B(_1070_),
    .C(\datapath.alu.b_4_bF$buf0 ),
    .Y(_1071_)
);

OAI21X1 _12234_ (
    .A(_2397_),
    .B(_2398_),
    .C(_1841__bF$buf3),
    .Y(_1072_)
);

OAI21X1 _12235_ (
    .A(_1841__bF$buf2),
    .B(_913_),
    .C(_1072_),
    .Y(_1073_)
);

AOI22X1 _12236_ (
    .A(_2398_),
    .B(_2536_),
    .C(_2054_),
    .D(_1073_),
    .Y(_1074_)
);

NOR2X1 _12237_ (
    .A(_1824__bF$buf2),
    .B(_1074_),
    .Y(_1076_)
);

NOR2X1 _12238_ (
    .A(_1777_),
    .B(_1779_),
    .Y(_1077_)
);

INVX1 _12239_ (
    .A(_1077_),
    .Y(_1078_)
);

OAI22X1 _12240_ (
    .A(_1078_),
    .B(_2014__bF$buf1),
    .C(_1778_),
    .D(_2017_),
    .Y(_1079_)
);

OAI22X1 _12241_ (
    .A(_1777_),
    .B(_2118__bF$buf2),
    .C(_1779_),
    .D(_2267__bF$buf2),
    .Y(_1080_)
);

NOR2X1 _12242_ (
    .A(_1080_),
    .B(_1079_),
    .Y(_1081_)
);

OAI21X1 _12243_ (
    .A(_1077_),
    .B(_2047__bF$buf0),
    .C(_2122_),
    .Y(_1082_)
);

OAI21X1 _12244_ (
    .A(\datapath.alu.a [14]),
    .B(\datapath.alu.b [14]),
    .C(_1082_),
    .Y(_1083_)
);

NAND2X1 _12245_ (
    .A(_1083_),
    .B(_1081_),
    .Y(_1084_)
);

NOR3X1 _12246_ (
    .A(_1084_),
    .B(_1076_),
    .C(_1071_),
    .Y(_1085_)
);

OAI21X1 _12247_ (
    .A(_1055_),
    .B(_1056_),
    .C(_1085_),
    .Y(_1087_)
);

AOI21X1 _12248_ (
    .A(_1049_),
    .B(_1051_),
    .C(_1087_),
    .Y(_1088_)
);

INVX1 _12249_ (
    .A(_1088_),
    .Y(\datapath.alu.c [14])
);

INVX1 _12250_ (
    .A(_1776_),
    .Y(_1089_)
);

AND2X2 _12251_ (
    .A(_1048_),
    .B(_1912_),
    .Y(_1090_)
);

OAI21X1 _12252_ (
    .A(_1077_),
    .B(_1090_),
    .C(_1089_),
    .Y(_1091_)
);

NAND3X1 _12253_ (
    .A(_1776_),
    .B(_1078_),
    .C(_1049_),
    .Y(_1092_)
);

NAND3X1 _12254_ (
    .A(_2045_),
    .B(_1092_),
    .C(_1091_),
    .Y(_1093_)
);

OAI21X1 _12255_ (
    .A(_1912_),
    .B(_1054_),
    .C(_1780_),
    .Y(_1094_)
);

AOI21X1 _12256_ (
    .A(_1094_),
    .B(_1776_),
    .C(_2134_),
    .Y(_1095_)
);

OAI21X1 _12257_ (
    .A(_1776_),
    .B(_1094_),
    .C(_1095_),
    .Y(_1097_)
);

AOI21X1 _12258_ (
    .A(_2448_),
    .B(_2445_),
    .C(\datapath.alu.b_3_bF$buf4 ),
    .Y(_1098_)
);

AOI21X1 _12259_ (
    .A(\datapath.alu.b_3_bF$buf3 ),
    .B(_2437_),
    .C(_1098_),
    .Y(_1099_)
);

OAI21X1 _12260_ (
    .A(\datapath.alu.b_0_bF$buf1 ),
    .B(_1773_),
    .C(_2103_),
    .Y(_1100_)
);

NAND2X1 _12261_ (
    .A(_1833__bF$buf4),
    .B(_1100_),
    .Y(_1101_)
);

OAI21X1 _12262_ (
    .A(_1833__bF$buf3),
    .B(_1031_),
    .C(_1101_),
    .Y(_1102_)
);

NAND2X1 _12263_ (
    .A(_1839__bF$buf5),
    .B(_1102_),
    .Y(_1103_)
);

OAI21X1 _12264_ (
    .A(_1839__bF$buf4),
    .B(_931_),
    .C(_1103_),
    .Y(_1104_)
);

MUX2X1 _12265_ (
    .A(_1104_),
    .B(_2460_),
    .S(_1841__bF$buf1),
    .Y(_1105_)
);

OAI22X1 _12266_ (
    .A(_1974_),
    .B(_1099_),
    .C(_2039_),
    .D(_1105_),
    .Y(_1106_)
);

NAND2X1 _12267_ (
    .A(\datapath.alu.a [31]),
    .B(_2054_),
    .Y(_1108_)
);

NAND2X1 _12268_ (
    .A(_1841__bF$buf0),
    .B(_2440_),
    .Y(_1109_)
);

OAI21X1 _12269_ (
    .A(_2142_),
    .B(_1109_),
    .C(_1108_),
    .Y(_1110_)
);

NAND2X1 _12270_ (
    .A(\datapath.alu.b_4_bF$buf4 ),
    .B(_1110_),
    .Y(_1111_)
);

OAI21X1 _12271_ (
    .A(\datapath.alu.a [15]),
    .B(_2017_),
    .C(_2267__bF$buf1),
    .Y(_1112_)
);

NAND2X1 _12272_ (
    .A(\datapath.alu.b [15]),
    .B(_1112_),
    .Y(_1113_)
);

OAI21X1 _12273_ (
    .A(\datapath.alu.a [15]),
    .B(\datapath.alu.b [15]),
    .C(_2027__bF$buf3),
    .Y(_1114_)
);

OAI21X1 _12274_ (
    .A(_1776_),
    .B(_2047__bF$buf3),
    .C(_1114_),
    .Y(_1115_)
);

OAI21X1 _12275_ (
    .A(_1774_),
    .B(_2014__bF$buf0),
    .C(_2118__bF$buf1),
    .Y(_1116_)
);

AOI21X1 _12276_ (
    .A(\datapath.alu.a [15]),
    .B(_1116_),
    .C(_1115_),
    .Y(_1117_)
);

NAND3X1 _12277_ (
    .A(_1113_),
    .B(_1117_),
    .C(_1111_),
    .Y(_1119_)
);

AOI21X1 _12278_ (
    .A(_1106_),
    .B(_1824__bF$buf1),
    .C(_1119_),
    .Y(_1120_)
);

NAND3X1 _12279_ (
    .A(_1097_),
    .B(_1120_),
    .C(_1093_),
    .Y(\datapath.alu.c [15])
);

INVX2 _12280_ (
    .A(_1408_),
    .Y(_1121_)
);

OAI21X1 _12281_ (
    .A(_2291_),
    .B(_2292_),
    .C(_2483_),
    .Y(_1122_)
);

NOR2X1 _12282_ (
    .A(_1776_),
    .B(_1781_),
    .Y(_1123_)
);

AND2X2 _12283_ (
    .A(_1123_),
    .B(_1043_),
    .Y(_1124_)
);

NAND2X1 _12284_ (
    .A(_954_),
    .B(_1124_),
    .Y(_1125_)
);

AOI21X1 _12285_ (
    .A(_1122_),
    .B(_2519_),
    .C(_1125_),
    .Y(_1126_)
);

NAND2X1 _12286_ (
    .A(_1043_),
    .B(_1123_),
    .Y(_1127_)
);

OAI21X1 _12287_ (
    .A(\datapath.alu.a [15]),
    .B(\datapath.alu.b [15]),
    .C(_1077_),
    .Y(_1129_)
);

OAI21X1 _12288_ (
    .A(_1773_),
    .B(_1774_),
    .C(_1129_),
    .Y(_1130_)
);

AOI21X1 _12289_ (
    .A(_1123_),
    .B(_1046_),
    .C(_1130_),
    .Y(_1131_)
);

OAI21X1 _12290_ (
    .A(_1127_),
    .B(_951_),
    .C(_1131_),
    .Y(_1132_)
);

OAI21X1 _12291_ (
    .A(_1132_),
    .B(_1126_),
    .C(_1121_),
    .Y(_1133_)
);

NAND3X1 _12292_ (
    .A(_1920_),
    .B(_1923_),
    .C(_949_),
    .Y(_1134_)
);

NOR2X1 _12293_ (
    .A(_1134_),
    .B(_1127_),
    .Y(_1135_)
);

AOI21X1 _12294_ (
    .A(_2520_),
    .B(_1135_),
    .C(_1132_),
    .Y(_1136_)
);

AOI21X1 _12295_ (
    .A(_1136_),
    .B(_1408_),
    .C(_2251__bF$buf1),
    .Y(_1137_)
);

AOI21X1 _12296_ (
    .A(_1796_),
    .B(_912_),
    .C(_963_),
    .Y(_1138_)
);

OAI21X1 _12297_ (
    .A(_1798_),
    .B(_873_),
    .C(_1138_),
    .Y(_1140_)
);

INVX1 _12298_ (
    .A(_1787_),
    .Y(_1141_)
);

OAI21X1 _12299_ (
    .A(_1141_),
    .B(_948_),
    .C(_1866_),
    .Y(_1142_)
);

NOR2X1 _12300_ (
    .A(\datapath.alu.b [14]),
    .B(_1777_),
    .Y(_1143_)
);

NOR2X1 _12301_ (
    .A(\datapath.alu.b [15]),
    .B(_1773_),
    .Y(_1144_)
);

AOI21X1 _12302_ (
    .A(_1776_),
    .B(_1143_),
    .C(_1144_),
    .Y(_1145_)
);

OAI21X1 _12303_ (
    .A(_1142_),
    .B(_1782_),
    .C(_1145_),
    .Y(_1146_)
);

AOI21X1 _12304_ (
    .A(_1791_),
    .B(_1140_),
    .C(_1146_),
    .Y(_1147_)
);

OAI21X1 _12305_ (
    .A(_1811_),
    .B(_2489_),
    .C(_1147_),
    .Y(_1148_)
);

NOR2X1 _12306_ (
    .A(_1408_),
    .B(_1148_),
    .Y(_1149_)
);

OAI21X1 _12307_ (
    .A(\datapath.alu.a [15]),
    .B(_1774_),
    .C(_1143_),
    .Y(_1151_)
);

OAI21X1 _12308_ (
    .A(_1773_),
    .B(\datapath.alu.b [15]),
    .C(_1151_),
    .Y(_1152_)
);

AOI21X1 _12309_ (
    .A(_1052_),
    .B(_1913_),
    .C(_1152_),
    .Y(_1153_)
);

OAI21X1 _12310_ (
    .A(_1915_),
    .B(_966_),
    .C(_1153_),
    .Y(_1154_)
);

AOI21X1 _12311_ (
    .A(_2529_),
    .B(_1926_),
    .C(_1154_),
    .Y(_1155_)
);

OAI21X1 _12312_ (
    .A(_1121_),
    .B(_1155_),
    .C(_2133__bF$buf1),
    .Y(_1156_)
);

NOR2X1 _12313_ (
    .A(_1824__bF$buf0),
    .B(_1108_),
    .Y(_1157_)
);

INVX2 _12314_ (
    .A(_1157_),
    .Y(_1158_)
);

NAND3X1 _12315_ (
    .A(_1975_),
    .B(_2007_),
    .C(_1992_),
    .Y(_1159_)
);

OAI21X1 _12316_ (
    .A(_1365_),
    .B(_2014__bF$buf3),
    .C(_2267__bF$buf0),
    .Y(_1160_)
);

AND2X2 _12317_ (
    .A(_1160_),
    .B(\datapath.alu.b [16]),
    .Y(_1162_)
);

OAI21X1 _12318_ (
    .A(\datapath.alu.a [16]),
    .B(\datapath.alu.b [16]),
    .C(_2027__bF$buf2),
    .Y(_1163_)
);

OAI21X1 _12319_ (
    .A(_1876_),
    .B(_2017_),
    .C(_1163_),
    .Y(_1164_)
);

OAI22X1 _12320_ (
    .A(_1365_),
    .B(_2118__bF$buf0),
    .C(_1408_),
    .D(_2047__bF$buf2),
    .Y(_1165_)
);

NOR3X1 _12321_ (
    .A(_1165_),
    .B(_1164_),
    .C(_1162_),
    .Y(_1166_)
);

NAND3X1 _12322_ (
    .A(_1158_),
    .B(_1159_),
    .C(_1166_),
    .Y(_1167_)
);

AND2X2 _12323_ (
    .A(_977_),
    .B(_980_),
    .Y(_1168_)
);

NAND2X1 _12324_ (
    .A(\datapath.alu.b_0_bF$buf0 ),
    .B(_1773_),
    .Y(_1169_)
);

OAI21X1 _12325_ (
    .A(\datapath.alu.b_0_bF$buf9 ),
    .B(\datapath.alu.a [16]),
    .C(_1169_),
    .Y(_1170_)
);

NAND2X1 _12326_ (
    .A(_1833__bF$buf2),
    .B(_1170_),
    .Y(_1171_)
);

OAI21X1 _12327_ (
    .A(_1833__bF$buf1),
    .B(_1060_),
    .C(_1171_),
    .Y(_1173_)
);

NAND2X1 _12328_ (
    .A(_1839__bF$buf3),
    .B(_1173_),
    .Y(_1174_)
);

OAI21X1 _12329_ (
    .A(_1839__bF$buf2),
    .B(_1168_),
    .C(_1174_),
    .Y(_1175_)
);

NAND2X1 _12330_ (
    .A(_2500_),
    .B(_2499_),
    .Y(_1176_)
);

AOI21X1 _12331_ (
    .A(_1176_),
    .B(\datapath.alu.b_3_bF$buf2 ),
    .C(\datapath.alu.b_4_bF$buf3 ),
    .Y(_1177_)
);

OAI21X1 _12332_ (
    .A(\datapath.alu.b_3_bF$buf1 ),
    .B(_1175_),
    .C(_1177_),
    .Y(_1178_)
);

NOR2X1 _12333_ (
    .A(_1824__bF$buf5),
    .B(_2035_),
    .Y(_1179_)
);

NOR2X1 _12334_ (
    .A(_2039_),
    .B(_1179_),
    .Y(_1180_)
);

AOI21X1 _12335_ (
    .A(_1178_),
    .B(_1180_),
    .C(_1167_),
    .Y(_1181_)
);

OAI21X1 _12336_ (
    .A(_1149_),
    .B(_1156_),
    .C(_1181_),
    .Y(_1182_)
);

AOI21X1 _12337_ (
    .A(_1133_),
    .B(_1137_),
    .C(_1182_),
    .Y(_1184_)
);

INVX1 _12338_ (
    .A(_1184_),
    .Y(\datapath.alu.c [16])
);

AND2X2 _12339_ (
    .A(_1133_),
    .B(_1397_),
    .Y(_1185_)
);

OR2X2 _12340_ (
    .A(_1185_),
    .B(_1354_),
    .Y(_1186_)
);

AOI21X1 _12341_ (
    .A(_1185_),
    .B(_1354_),
    .C(_2251__bF$buf0),
    .Y(_1187_)
);

NAND2X1 _12342_ (
    .A(\datapath.alu.a [16]),
    .B(_1375_),
    .Y(_1188_)
);

OAI21X1 _12343_ (
    .A(_1121_),
    .B(_1155_),
    .C(_1188_),
    .Y(_1189_)
);

AND2X2 _12344_ (
    .A(_1189_),
    .B(_1354_),
    .Y(_1190_)
);

OAI21X1 _12345_ (
    .A(_1354_),
    .B(_1189_),
    .C(_2133__bF$buf0),
    .Y(_1191_)
);

NAND2X1 _12346_ (
    .A(\datapath.alu.b_2_bF$buf2 ),
    .B(_1034_),
    .Y(_1192_)
);

NAND2X1 _12347_ (
    .A(\datapath.alu.b_1_bF$buf6 ),
    .B(_1100_),
    .Y(_1194_)
);

NAND2X1 _12348_ (
    .A(\datapath.alu.b_0_bF$buf8 ),
    .B(_1365_),
    .Y(_1195_)
);

OAI21X1 _12349_ (
    .A(\datapath.alu.b_0_bF$buf7 ),
    .B(\datapath.alu.a [17]),
    .C(_1195_),
    .Y(_1196_)
);

OAI21X1 _12350_ (
    .A(\datapath.alu.b_1_bF$buf5 ),
    .B(_1196_),
    .C(_1194_),
    .Y(_1197_)
);

NAND2X1 _12351_ (
    .A(_1839__bF$buf1),
    .B(_1197_),
    .Y(_1198_)
);

AOI21X1 _12352_ (
    .A(_1192_),
    .B(_1198_),
    .C(\datapath.alu.b_3_bF$buf0 ),
    .Y(_1199_)
);

NOR2X1 _12353_ (
    .A(_1841__bF$buf7),
    .B(_2548_),
    .Y(_1200_)
);

OAI21X1 _12354_ (
    .A(_1199_),
    .B(_1200_),
    .C(_976_),
    .Y(_1201_)
);

NAND3X1 _12355_ (
    .A(_2082_),
    .B(_2088_),
    .C(_1201_),
    .Y(_1202_)
);

OAI21X1 _12356_ (
    .A(\datapath.alu.a [17]),
    .B(_2017_),
    .C(_2267__bF$buf3),
    .Y(_1203_)
);

OAI22X1 _12357_ (
    .A(_1322_),
    .B(_2118__bF$buf3),
    .C(_1311_),
    .D(_2014__bF$buf2),
    .Y(_1205_)
);

OAI21X1 _12358_ (
    .A(\datapath.alu.a [17]),
    .B(\datapath.alu.b [17]),
    .C(_2027__bF$buf1),
    .Y(_1206_)
);

OAI21X1 _12359_ (
    .A(_1354_),
    .B(_2047__bF$buf1),
    .C(_1206_),
    .Y(_1207_)
);

NOR2X1 _12360_ (
    .A(_1205_),
    .B(_1207_),
    .Y(_1208_)
);

OAI21X1 _12361_ (
    .A(_1824__bF$buf4),
    .B(_1108_),
    .C(_1208_),
    .Y(_1209_)
);

AOI21X1 _12362_ (
    .A(\datapath.alu.b [17]),
    .B(_1203_),
    .C(_1209_),
    .Y(_1210_)
);

NOR2X1 _12363_ (
    .A(_1824__bF$buf3),
    .B(_2039_),
    .Y(_1211_)
);

INVX2 _12364_ (
    .A(_1211_),
    .Y(_1212_)
);

OAI21X1 _12365_ (
    .A(_2131_),
    .B(_1212_),
    .C(_1210_),
    .Y(_1213_)
);

AOI21X1 _12366_ (
    .A(_1202_),
    .B(_1824__bF$buf2),
    .C(_1213_),
    .Y(_1214_)
);

OAI21X1 _12367_ (
    .A(_1190_),
    .B(_1191_),
    .C(_1214_),
    .Y(_1216_)
);

AOI21X1 _12368_ (
    .A(_1186_),
    .B(_1187_),
    .C(_1216_),
    .Y(_1217_)
);

INVX1 _12369_ (
    .A(_1217_),
    .Y(\datapath.alu.c [17])
);

INVX2 _12370_ (
    .A(_1290_),
    .Y(_1218_)
);

INVX1 _12371_ (
    .A(_1354_),
    .Y(_1219_)
);

NAND2X1 _12372_ (
    .A(_1219_),
    .B(_1121_),
    .Y(_1220_)
);

OAI21X1 _12373_ (
    .A(_1322_),
    .B(_1333_),
    .C(_1397_),
    .Y(_1221_)
);

OAI21X1 _12374_ (
    .A(\datapath.alu.a [17]),
    .B(\datapath.alu.b [17]),
    .C(_1221_),
    .Y(_1222_)
);

OAI21X1 _12375_ (
    .A(_1220_),
    .B(_1136_),
    .C(_1222_),
    .Y(_1223_)
);

NAND2X1 _12376_ (
    .A(_1218_),
    .B(_1223_),
    .Y(_1224_)
);

NOR2X1 _12377_ (
    .A(_1218_),
    .B(_1223_),
    .Y(_1226_)
);

NOR2X1 _12378_ (
    .A(_2251__bF$buf3),
    .B(_1226_),
    .Y(_1227_)
);

NAND2X1 _12379_ (
    .A(\datapath.alu.a [17]),
    .B(_1333_),
    .Y(_1228_)
);

OAI21X1 _12380_ (
    .A(_1365_),
    .B(\datapath.alu.b [16]),
    .C(_1228_),
    .Y(_1229_)
);

OAI21X1 _12381_ (
    .A(\datapath.alu.a [17]),
    .B(_1333_),
    .C(_1229_),
    .Y(_1230_)
);

OAI21X1 _12382_ (
    .A(_1418_),
    .B(_1155_),
    .C(_1230_),
    .Y(_1231_)
);

NOR2X1 _12383_ (
    .A(_1290_),
    .B(_1231_),
    .Y(_1232_)
);

INVX1 _12384_ (
    .A(_1418_),
    .Y(_1233_)
);

INVX1 _12385_ (
    .A(_1230_),
    .Y(_1234_)
);

AOI21X1 _12386_ (
    .A(_1148_),
    .B(_1233_),
    .C(_1234_),
    .Y(_1235_)
);

OAI21X1 _12387_ (
    .A(_1218_),
    .B(_1235_),
    .C(_2133__bF$buf3),
    .Y(_1237_)
);

INVX1 _12388_ (
    .A(_1279_),
    .Y(_1238_)
);

AOI22X1 _12389_ (
    .A(_2197_),
    .B(_1238_),
    .C(\datapath.alu.a [18]),
    .D(_2022_),
    .Y(_1239_)
);

AOI21X1 _12390_ (
    .A(_1247_),
    .B(_2016__bF$buf1),
    .C(_2029_),
    .Y(_1240_)
);

OAI21X1 _12391_ (
    .A(_1258_),
    .B(_1240_),
    .C(_1239_),
    .Y(_1241_)
);

OAI21X1 _12392_ (
    .A(\datapath.alu.a [18]),
    .B(\datapath.alu.b [18]),
    .C(_2027__bF$buf0),
    .Y(_1242_)
);

OAI21X1 _12393_ (
    .A(_1290_),
    .B(_2047__bF$buf0),
    .C(_1242_),
    .Y(_1243_)
);

NOR2X1 _12394_ (
    .A(_1243_),
    .B(_1241_),
    .Y(_1244_)
);

AND2X2 _12395_ (
    .A(_1244_),
    .B(_1158_),
    .Y(_1245_)
);

OAI21X1 _12396_ (
    .A(_1839__bF$buf0),
    .B(_2414_),
    .C(_898_),
    .Y(_1246_)
);

MUX2X1 _12397_ (
    .A(_1322_),
    .B(_1247_),
    .S(\datapath.alu.b_0_bF$buf6 ),
    .Y(_1248_)
);

NAND2X1 _12398_ (
    .A(\datapath.alu.b_1_bF$buf4 ),
    .B(_1170_),
    .Y(_1249_)
);

OAI21X1 _12399_ (
    .A(\datapath.alu.b_1_bF$buf3 ),
    .B(_1248_),
    .C(_1249_),
    .Y(_1250_)
);

NAND2X1 _12400_ (
    .A(_1839__bF$buf6),
    .B(_1250_),
    .Y(_1251_)
);

OAI21X1 _12401_ (
    .A(_1839__bF$buf5),
    .B(_1062_),
    .C(_1251_),
    .Y(_1252_)
);

OAI21X1 _12402_ (
    .A(\datapath.alu.b_3_bF$buf7 ),
    .B(_1252_),
    .C(_1824__bF$buf1),
    .Y(_1253_)
);

AOI21X1 _12403_ (
    .A(\datapath.alu.b_3_bF$buf6 ),
    .B(_1246_),
    .C(_1253_),
    .Y(_1254_)
);

AOI21X1 _12404_ (
    .A(_2181_),
    .B(_2180_),
    .C(_2040_),
    .Y(_1255_)
);

OAI21X1 _12405_ (
    .A(_1255_),
    .B(_1254_),
    .C(_1245_),
    .Y(_1256_)
);

AOI21X1 _12406_ (
    .A(_1824__bF$buf0),
    .B(_2161_),
    .C(_1256_),
    .Y(_1257_)
);

OAI21X1 _12407_ (
    .A(_1232_),
    .B(_1237_),
    .C(_1257_),
    .Y(_1259_)
);

AOI21X1 _12408_ (
    .A(_1227_),
    .B(_1224_),
    .C(_1259_),
    .Y(_1260_)
);

INVX1 _12409_ (
    .A(_1260_),
    .Y(\datapath.alu.c [18])
);

NOR2X1 _12410_ (
    .A(_1236_),
    .B(_1225_),
    .Y(_1261_)
);

AND2X2 _12411_ (
    .A(_1223_),
    .B(_1218_),
    .Y(_1262_)
);

OAI21X1 _12412_ (
    .A(_1238_),
    .B(_1262_),
    .C(_1261_),
    .Y(_1263_)
);

INVX2 _12413_ (
    .A(_1261_),
    .Y(_1264_)
);

NAND3X1 _12414_ (
    .A(_1264_),
    .B(_1279_),
    .C(_1224_),
    .Y(_1265_)
);

NAND3X1 _12415_ (
    .A(_2045_),
    .B(_1265_),
    .C(_1263_),
    .Y(_1266_)
);

NAND2X1 _12416_ (
    .A(\datapath.alu.a [18]),
    .B(_1258_),
    .Y(_1267_)
);

OAI21X1 _12417_ (
    .A(_1218_),
    .B(_1235_),
    .C(_1267_),
    .Y(_1269_)
);

AOI21X1 _12418_ (
    .A(_1269_),
    .B(_1264_),
    .C(_2134_),
    .Y(_1270_)
);

OAI21X1 _12419_ (
    .A(_1264_),
    .B(_1269_),
    .C(_1270_),
    .Y(_1271_)
);

OAI21X1 _12420_ (
    .A(\datapath.alu.b_3_bF$buf5 ),
    .B(_918_),
    .C(_2239_),
    .Y(_1272_)
);

NAND2X1 _12421_ (
    .A(_2054_),
    .B(_1272_),
    .Y(_1273_)
);

AND2X2 _12422_ (
    .A(_2234_),
    .B(_2244_),
    .Y(_1274_)
);

OAI21X1 _12423_ (
    .A(_2142_),
    .B(_1274_),
    .C(_1273_),
    .Y(_1275_)
);

OAI21X1 _12424_ (
    .A(\datapath.alu.a [19]),
    .B(_2017_),
    .C(_2267__bF$buf2),
    .Y(_1276_)
);

NAND2X1 _12425_ (
    .A(\datapath.alu.b [19]),
    .B(_1276_),
    .Y(_1277_)
);

NAND2X1 _12426_ (
    .A(_1225_),
    .B(_2197_),
    .Y(_1278_)
);

OAI21X1 _12427_ (
    .A(_1204_),
    .B(_2118__bF$buf2),
    .C(_1278_),
    .Y(_1280_)
);

OAI22X1 _12428_ (
    .A(_1236_),
    .B(_2122_),
    .C(_2047__bF$buf3),
    .D(_1264_),
    .Y(_1281_)
);

NOR2X1 _12429_ (
    .A(_1280_),
    .B(_1281_),
    .Y(_1282_)
);

NAND3X1 _12430_ (
    .A(_1277_),
    .B(_1158_),
    .C(_1282_),
    .Y(_1283_)
);

AOI21X1 _12431_ (
    .A(_1275_),
    .B(_1824__bF$buf5),
    .C(_1283_),
    .Y(_1284_)
);

NOR2X1 _12432_ (
    .A(_2061_),
    .B(_2065_),
    .Y(_1285_)
);

NAND2X1 _12433_ (
    .A(_1833__bF$buf0),
    .B(_1285_),
    .Y(_1286_)
);

OAI21X1 _12434_ (
    .A(_1833__bF$buf7),
    .B(_1196_),
    .C(_1286_),
    .Y(_1287_)
);

MUX2X1 _12435_ (
    .A(_1287_),
    .B(_1102_),
    .S(_1839__bF$buf4),
    .Y(_1288_)
);

NOR2X1 _12436_ (
    .A(\datapath.alu.b_3_bF$buf4 ),
    .B(_1288_),
    .Y(_1289_)
);

OAI21X1 _12437_ (
    .A(_1841__bF$buf6),
    .B(_933_),
    .C(_1824__bF$buf4),
    .Y(_1291_)
);

NAND2X1 _12438_ (
    .A(_1841__bF$buf5),
    .B(_2263_),
    .Y(_1292_)
);

AOI21X1 _12439_ (
    .A(_1292_),
    .B(\datapath.alu.b_4_bF$buf2 ),
    .C(_2039_),
    .Y(_1293_)
);

OAI21X1 _12440_ (
    .A(_1291_),
    .B(_1289_),
    .C(_1293_),
    .Y(_1294_)
);

AND2X2 _12441_ (
    .A(_1284_),
    .B(_1294_),
    .Y(_1295_)
);

NAND3X1 _12442_ (
    .A(_1271_),
    .B(_1295_),
    .C(_1266_),
    .Y(\datapath.alu.c [19])
);

INVX2 _12443_ (
    .A(_1172_),
    .Y(_1296_)
);

NAND2X1 _12444_ (
    .A(_1261_),
    .B(_1218_),
    .Y(_1297_)
);

AOI21X1 _12445_ (
    .A(_1261_),
    .B(_1238_),
    .C(_1225_),
    .Y(_1298_)
);

OAI21X1 _12446_ (
    .A(_1222_),
    .B(_1297_),
    .C(_1298_),
    .Y(_1299_)
);

INVX1 _12447_ (
    .A(_1299_),
    .Y(_1301_)
);

NOR2X1 _12448_ (
    .A(_1297_),
    .B(_1220_),
    .Y(_1302_)
);

INVX1 _12449_ (
    .A(_1302_),
    .Y(_1303_)
);

OAI21X1 _12450_ (
    .A(_1303_),
    .B(_1136_),
    .C(_1301_),
    .Y(_1304_)
);

NAND2X1 _12451_ (
    .A(_1296_),
    .B(_1304_),
    .Y(_1305_)
);

OAI21X1 _12452_ (
    .A(_1132_),
    .B(_1126_),
    .C(_1302_),
    .Y(_1306_)
);

NAND3X1 _12453_ (
    .A(_1172_),
    .B(_1301_),
    .C(_1306_),
    .Y(_1307_)
);

NAND3X1 _12454_ (
    .A(_2045_),
    .B(_1307_),
    .C(_1305_),
    .Y(_1308_)
);

OAI21X1 _12455_ (
    .A(_1267_),
    .B(_1881_),
    .C(_1879_),
    .Y(_1309_)
);

INVX1 _12456_ (
    .A(_1309_),
    .Y(_1310_)
);

OAI21X1 _12457_ (
    .A(_1300_),
    .B(_1230_),
    .C(_1310_),
    .Y(_1312_)
);

AOI21X1 _12458_ (
    .A(_1148_),
    .B(_1429_),
    .C(_1312_),
    .Y(_1313_)
);

NAND2X1 _12459_ (
    .A(_1296_),
    .B(_1313_),
    .Y(_1314_)
);

INVX1 _12460_ (
    .A(_1429_),
    .Y(_1315_)
);

INVX1 _12461_ (
    .A(_1312_),
    .Y(_1316_)
);

OAI21X1 _12462_ (
    .A(_1315_),
    .B(_1155_),
    .C(_1316_),
    .Y(_1317_)
);

AOI21X1 _12463_ (
    .A(_1317_),
    .B(_1172_),
    .C(_2134_),
    .Y(_1318_)
);

NAND2X1 _12464_ (
    .A(_1314_),
    .B(_1318_),
    .Y(_1319_)
);

NOR2X1 _12465_ (
    .A(_2285_),
    .B(_2283_),
    .Y(_1320_)
);

NAND2X1 _12466_ (
    .A(\datapath.alu.b_0_bF$buf5 ),
    .B(_1204_),
    .Y(_1321_)
);

OAI21X1 _12467_ (
    .A(\datapath.alu.b_0_bF$buf4 ),
    .B(\datapath.alu.a [20]),
    .C(_1321_),
    .Y(_1323_)
);

NAND2X1 _12468_ (
    .A(_1833__bF$buf6),
    .B(_1323_),
    .Y(_1324_)
);

OAI21X1 _12469_ (
    .A(_1833__bF$buf5),
    .B(_1248_),
    .C(_1324_),
    .Y(_1325_)
);

MUX2X1 _12470_ (
    .A(_1325_),
    .B(_1173_),
    .S(_1839__bF$buf3),
    .Y(_1326_)
);

NAND3X1 _12471_ (
    .A(\datapath.alu.b_3_bF$buf3 ),
    .B(_981_),
    .C(_982_),
    .Y(_1327_)
);

OAI21X1 _12472_ (
    .A(\datapath.alu.b_3_bF$buf2 ),
    .B(_1326_),
    .C(_1327_),
    .Y(_1328_)
);

OAI21X1 _12473_ (
    .A(_2039_),
    .B(_1328_),
    .C(_1320_),
    .Y(_1329_)
);

OAI21X1 _12474_ (
    .A(\datapath.alu.a [20]),
    .B(_2017_),
    .C(_2267__bF$buf1),
    .Y(_1330_)
);

NAND2X1 _12475_ (
    .A(\datapath.alu.b [20]),
    .B(_1330_),
    .Y(_1331_)
);

INVX1 _12476_ (
    .A(_1161_),
    .Y(_1332_)
);

AOI22X1 _12477_ (
    .A(_2197_),
    .B(_1332_),
    .C(_2553_),
    .D(_1296_),
    .Y(_1334_)
);

AOI22X1 _12478_ (
    .A(_2022_),
    .B(\datapath.alu.a [20]),
    .C(_1150_),
    .D(_2027__bF$buf3),
    .Y(_1335_)
);

NAND3X1 _12479_ (
    .A(_1334_),
    .B(_1335_),
    .C(_1331_),
    .Y(_1336_)
);

NOR2X1 _12480_ (
    .A(_1157_),
    .B(_1336_),
    .Y(_1337_)
);

OAI21X1 _12481_ (
    .A(_2313_),
    .B(_1212_),
    .C(_1337_),
    .Y(_1338_)
);

AOI21X1 _12482_ (
    .A(_1329_),
    .B(_1824__bF$buf3),
    .C(_1338_),
    .Y(_1339_)
);

NAND3X1 _12483_ (
    .A(_1339_),
    .B(_1308_),
    .C(_1319_),
    .Y(\datapath.alu.c [20])
);

AOI21X1 _12484_ (
    .A(_1304_),
    .B(_1296_),
    .C(_1332_),
    .Y(_1340_)
);

OR2X2 _12485_ (
    .A(_1340_),
    .B(_1118_),
    .Y(_1341_)
);

AOI21X1 _12486_ (
    .A(_1340_),
    .B(_1118_),
    .C(_2251__bF$buf2),
    .Y(_1342_)
);

INVX1 _12487_ (
    .A(_1118_),
    .Y(_1344_)
);

OAI21X1 _12488_ (
    .A(_1128_),
    .B(\datapath.alu.b [20]),
    .C(_1344_),
    .Y(_1345_)
);

AOI21X1 _12489_ (
    .A(_1317_),
    .B(_1172_),
    .C(_1345_),
    .Y(_1346_)
);

NOR2X1 _12490_ (
    .A(\datapath.alu.b [20]),
    .B(_1128_),
    .Y(_1347_)
);

NAND2X1 _12491_ (
    .A(_1347_),
    .B(_1118_),
    .Y(_1348_)
);

AND2X2 _12492_ (
    .A(_1348_),
    .B(_2133__bF$buf2),
    .Y(_1349_)
);

OAI21X1 _12493_ (
    .A(_1183_),
    .B(_1313_),
    .C(_1349_),
    .Y(_1350_)
);

NAND2X1 _12494_ (
    .A(\datapath.alu.b_2_bF$buf1 ),
    .B(_1197_),
    .Y(_1351_)
);

NAND2X1 _12495_ (
    .A(\datapath.alu.b_0_bF$buf3 ),
    .B(_1128_),
    .Y(_1352_)
);

OAI21X1 _12496_ (
    .A(\datapath.alu.b_0_bF$buf2 ),
    .B(\datapath.alu.a [21]),
    .C(_1352_),
    .Y(_1353_)
);

NAND2X1 _12497_ (
    .A(_1833__bF$buf4),
    .B(_1353_),
    .Y(_1355_)
);

OAI21X1 _12498_ (
    .A(_1833__bF$buf3),
    .B(_1285_),
    .C(_1355_),
    .Y(_1356_)
);

OAI21X1 _12499_ (
    .A(\datapath.alu.b_2_bF$buf0 ),
    .B(_1356_),
    .C(_1351_),
    .Y(_1357_)
);

OAI21X1 _12500_ (
    .A(_1841__bF$buf4),
    .B(_1035_),
    .C(_1824__bF$buf2),
    .Y(_1358_)
);

AOI21X1 _12501_ (
    .A(_1841__bF$buf3),
    .B(_1357_),
    .C(_1358_),
    .Y(_1359_)
);

AND2X2 _12502_ (
    .A(_2367_),
    .B(_1841__bF$buf2),
    .Y(_1360_)
);

OAI21X1 _12503_ (
    .A(_1824__bF$buf1),
    .B(_1360_),
    .C(_976_),
    .Y(_1361_)
);

AOI21X1 _12504_ (
    .A(_2197_),
    .B(\datapath.alu.b [21]),
    .C(_2022_),
    .Y(_1362_)
);

AOI21X1 _12505_ (
    .A(_2553_),
    .B(_1075_),
    .C(_2027__bF$buf2),
    .Y(_1363_)
);

OAI21X1 _12506_ (
    .A(_1086_),
    .B(_1362_),
    .C(_1363_),
    .Y(_1364_)
);

AOI21X1 _12507_ (
    .A(_1086_),
    .B(_2016__bF$buf0),
    .C(_2029_),
    .Y(_1366_)
);

OAI21X1 _12508_ (
    .A(_1096_),
    .B(_1366_),
    .C(_1158_),
    .Y(_1367_)
);

AOI21X1 _12509_ (
    .A(_1107_),
    .B(_1364_),
    .C(_1367_),
    .Y(_1368_)
);

OAI21X1 _12510_ (
    .A(_1361_),
    .B(_1359_),
    .C(_1368_),
    .Y(_1369_)
);

AOI21X1 _12511_ (
    .A(_1824__bF$buf0),
    .B(_2349_),
    .C(_1369_),
    .Y(_1370_)
);

OAI21X1 _12512_ (
    .A(_1346_),
    .B(_1350_),
    .C(_1370_),
    .Y(_1371_)
);

AOI21X1 _12513_ (
    .A(_1341_),
    .B(_1342_),
    .C(_1371_),
    .Y(_1372_)
);

INVX1 _12514_ (
    .A(_1372_),
    .Y(\datapath.alu.c [21])
);

NOR2X1 _12515_ (
    .A(_1118_),
    .B(_1172_),
    .Y(_1373_)
);

OAI21X1 _12516_ (
    .A(_1161_),
    .B(_1118_),
    .C(_1075_),
    .Y(_1374_)
);

AOI21X1 _12517_ (
    .A(_1304_),
    .B(_1373_),
    .C(_1374_),
    .Y(_1376_)
);

AOI21X1 _12518_ (
    .A(_1376_),
    .B(_1053_),
    .C(_2251__bF$buf1),
    .Y(_1377_)
);

OAI21X1 _12519_ (
    .A(_1053_),
    .B(_1376_),
    .C(_1377_),
    .Y(_1378_)
);

NOR2X1 _12520_ (
    .A(\datapath.alu.b [21]),
    .B(_1086_),
    .Y(_1379_)
);

AOI21X1 _12521_ (
    .A(_1118_),
    .B(_1347_),
    .C(_1379_),
    .Y(_1380_)
);

OAI21X1 _12522_ (
    .A(_1183_),
    .B(_1313_),
    .C(_1380_),
    .Y(_1381_)
);

NAND2X1 _12523_ (
    .A(_1053_),
    .B(_1381_),
    .Y(_1382_)
);

INVX1 _12524_ (
    .A(_1053_),
    .Y(_1383_)
);

INVX1 _12525_ (
    .A(_1183_),
    .Y(_1384_)
);

INVX1 _12526_ (
    .A(_1380_),
    .Y(_1385_)
);

AOI21X1 _12527_ (
    .A(_1317_),
    .B(_1384_),
    .C(_1385_),
    .Y(_1387_)
);

AOI21X1 _12528_ (
    .A(_1387_),
    .B(_1383_),
    .C(_2134_),
    .Y(_1388_)
);

OR2X2 _12529_ (
    .A(_2400_),
    .B(_2402_),
    .Y(_1389_)
);

OAI21X1 _12530_ (
    .A(\datapath.alu.a [22]),
    .B(_2017_),
    .C(_2267__bF$buf0),
    .Y(_1390_)
);

OAI21X1 _12531_ (
    .A(\datapath.alu.a [22]),
    .B(\datapath.alu.b [22]),
    .C(_2027__bF$buf1),
    .Y(_1391_)
);

INVX2 _12532_ (
    .A(_1042_),
    .Y(_1392_)
);

AOI22X1 _12533_ (
    .A(_2197_),
    .B(_1392_),
    .C(_2553_),
    .D(_1383_),
    .Y(_1393_)
);

NAND3X1 _12534_ (
    .A(_1391_),
    .B(_1393_),
    .C(_1158_),
    .Y(_1394_)
);

AOI21X1 _12535_ (
    .A(\datapath.alu.b [22]),
    .B(_1390_),
    .C(_1394_),
    .Y(_1395_)
);

OAI21X1 _12536_ (
    .A(_1010_),
    .B(_2118__bF$buf1),
    .C(_1395_),
    .Y(_1396_)
);

AOI21X1 _12537_ (
    .A(_1389_),
    .B(_1824__bF$buf5),
    .C(_1396_),
    .Y(_1398_)
);

MUX2X1 _12538_ (
    .A(_1086_),
    .B(_1010_),
    .S(\datapath.alu.b_0_bF$buf1 ),
    .Y(_1399_)
);

NAND2X1 _12539_ (
    .A(_1833__bF$buf2),
    .B(_1399_),
    .Y(_1400_)
);

OAI21X1 _12540_ (
    .A(_1833__bF$buf1),
    .B(_1323_),
    .C(_1400_),
    .Y(_1401_)
);

NAND2X1 _12541_ (
    .A(\datapath.alu.b_2_bF$buf7 ),
    .B(_1250_),
    .Y(_1402_)
);

OAI21X1 _12542_ (
    .A(\datapath.alu.b_2_bF$buf6 ),
    .B(_1401_),
    .C(_1402_),
    .Y(_1403_)
);

NOR2X1 _12543_ (
    .A(\datapath.alu.b_3_bF$buf1 ),
    .B(_1403_),
    .Y(_1404_)
);

OAI21X1 _12544_ (
    .A(_1841__bF$buf1),
    .B(_1063_),
    .C(_1824__bF$buf4),
    .Y(_1405_)
);

OAI21X1 _12545_ (
    .A(\datapath.alu.b_3_bF$buf0 ),
    .B(_1057_),
    .C(\datapath.alu.b_4_bF$buf1 ),
    .Y(_1406_)
);

OAI21X1 _12546_ (
    .A(_1405_),
    .B(_1404_),
    .C(_1406_),
    .Y(_1407_)
);

OAI21X1 _12547_ (
    .A(_2039_),
    .B(_1407_),
    .C(_1398_),
    .Y(_1409_)
);

AOI21X1 _12548_ (
    .A(_1388_),
    .B(_1382_),
    .C(_1409_),
    .Y(_1410_)
);

NAND2X1 _12549_ (
    .A(_1378_),
    .B(_1410_),
    .Y(\datapath.alu.c [22])
);

INVX2 _12550_ (
    .A(_1000_),
    .Y(_1411_)
);

NOR2X1 _12551_ (
    .A(_1053_),
    .B(_1376_),
    .Y(_1412_)
);

OAI21X1 _12552_ (
    .A(_1392_),
    .B(_1412_),
    .C(_1411_),
    .Y(_1413_)
);

NOR2X1 _12553_ (
    .A(_1392_),
    .B(_1412_),
    .Y(_1414_)
);

AOI21X1 _12554_ (
    .A(_1414_),
    .B(_1000_),
    .C(_2251__bF$buf0),
    .Y(_1415_)
);

NOR2X1 _12555_ (
    .A(\datapath.alu.b [22]),
    .B(_1010_),
    .Y(_1416_)
);

AOI21X1 _12556_ (
    .A(_1381_),
    .B(_1053_),
    .C(_1416_),
    .Y(_1417_)
);

AND2X2 _12557_ (
    .A(_1417_),
    .B(_1411_),
    .Y(_1419_)
);

OAI21X1 _12558_ (
    .A(_1411_),
    .B(_1417_),
    .C(_2133__bF$buf1),
    .Y(_1420_)
);

INVX1 _12559_ (
    .A(_2442_),
    .Y(_1421_)
);

MUX2X1 _12560_ (
    .A(_1010_),
    .B(_967_),
    .S(\datapath.alu.b_0_bF$buf0 ),
    .Y(_1422_)
);

NAND2X1 _12561_ (
    .A(_1833__bF$buf0),
    .B(_1422_),
    .Y(_1423_)
);

OAI21X1 _12562_ (
    .A(_1833__bF$buf7),
    .B(_1353_),
    .C(_1423_),
    .Y(_1424_)
);

MUX2X1 _12563_ (
    .A(_1287_),
    .B(_1424_),
    .S(\datapath.alu.b_2_bF$buf5 ),
    .Y(_1425_)
);

NAND2X1 _12564_ (
    .A(_1841__bF$buf0),
    .B(_1425_),
    .Y(_1426_)
);

OAI21X1 _12565_ (
    .A(_1841__bF$buf7),
    .B(_1104_),
    .C(_1426_),
    .Y(_1427_)
);

OAI21X1 _12566_ (
    .A(_2039_),
    .B(_1427_),
    .C(_1421_),
    .Y(_1428_)
);

NAND2X1 _12567_ (
    .A(_1841__bF$buf6),
    .B(_2460_),
    .Y(_1430_)
);

NOR2X1 _12568_ (
    .A(_956_),
    .B(_2014__bF$buf1),
    .Y(_1431_)
);

AOI21X1 _12569_ (
    .A(_1411_),
    .B(_2553_),
    .C(_1431_),
    .Y(_1432_)
);

AOI22X1 _12570_ (
    .A(_1888_),
    .B(_2016__bF$buf3),
    .C(\datapath.alu.b [23]),
    .D(_2029_),
    .Y(_1433_)
);

AOI21X1 _12571_ (
    .A(_989_),
    .B(_2027__bF$buf0),
    .C(_1157_),
    .Y(_1434_)
);

NAND3X1 _12572_ (
    .A(_1432_),
    .B(_1433_),
    .C(_1434_),
    .Y(_1435_)
);

AOI21X1 _12573_ (
    .A(\datapath.alu.a [23]),
    .B(_2022_),
    .C(_1435_),
    .Y(_1436_)
);

OAI21X1 _12574_ (
    .A(_1430_),
    .B(_1212_),
    .C(_1436_),
    .Y(_1437_)
);

AOI21X1 _12575_ (
    .A(_1428_),
    .B(_1824__bF$buf3),
    .C(_1437_),
    .Y(_1438_)
);

OAI21X1 _12576_ (
    .A(_1419_),
    .B(_1420_),
    .C(_1438_),
    .Y(_1439_)
);

AOI21X1 _12577_ (
    .A(_1415_),
    .B(_1413_),
    .C(_1439_),
    .Y(_1441_)
);

INVX1 _12578_ (
    .A(_1441_),
    .Y(\datapath.alu.c [23])
);

NOR2X1 _12579_ (
    .A(_1764_),
    .B(_1767_),
    .Y(_1442_)
);

OAI21X1 _12580_ (
    .A(_2480_),
    .B(_2477_),
    .C(_1135_),
    .Y(_1443_)
);

INVX1 _12581_ (
    .A(_1132_),
    .Y(_1444_)
);

NOR2X1 _12582_ (
    .A(_1000_),
    .B(_1053_),
    .Y(_1445_)
);

AND2X2 _12583_ (
    .A(_1373_),
    .B(_1445_),
    .Y(_1446_)
);

NAND2X1 _12584_ (
    .A(_1446_),
    .B(_1302_),
    .Y(_1447_)
);

AOI21X1 _12585_ (
    .A(_1444_),
    .B(_1443_),
    .C(_1447_),
    .Y(_1448_)
);

NAND2X1 _12586_ (
    .A(_1445_),
    .B(_1374_),
    .Y(_1449_)
);

OAI21X1 _12587_ (
    .A(\datapath.alu.a [23]),
    .B(\datapath.alu.b [23]),
    .C(_1392_),
    .Y(_1451_)
);

AND2X2 _12588_ (
    .A(_1451_),
    .B(_956_),
    .Y(_1452_)
);

NAND2X1 _12589_ (
    .A(_1452_),
    .B(_1449_),
    .Y(_1453_)
);

AOI21X1 _12590_ (
    .A(_1299_),
    .B(_1446_),
    .C(_1453_),
    .Y(_1454_)
);

INVX1 _12591_ (
    .A(_1454_),
    .Y(_1455_)
);

OAI21X1 _12592_ (
    .A(_1455_),
    .B(_1448_),
    .C(_1442_),
    .Y(_1456_)
);

INVX2 _12593_ (
    .A(_1442_),
    .Y(_1457_)
);

INVX1 _12594_ (
    .A(_1447_),
    .Y(_1458_)
);

OAI21X1 _12595_ (
    .A(_1132_),
    .B(_1126_),
    .C(_1458_),
    .Y(_1459_)
);

NAND3X1 _12596_ (
    .A(_1457_),
    .B(_1454_),
    .C(_1459_),
    .Y(_1460_)
);

NAND3X1 _12597_ (
    .A(_2045_),
    .B(_1460_),
    .C(_1456_),
    .Y(_1462_)
);

INVX1 _12598_ (
    .A(_1440_),
    .Y(_1463_)
);

INVX1 _12599_ (
    .A(_1886_),
    .Y(_1464_)
);

AOI21X1 _12600_ (
    .A(_1000_),
    .B(_1416_),
    .C(_1464_),
    .Y(_1465_)
);

OAI21X1 _12601_ (
    .A(_1064_),
    .B(_1380_),
    .C(_1465_),
    .Y(_1466_)
);

AOI21X1 _12602_ (
    .A(_1312_),
    .B(_1193_),
    .C(_1466_),
    .Y(_1467_)
);

INVX1 _12603_ (
    .A(_1467_),
    .Y(_1468_)
);

AOI21X1 _12604_ (
    .A(_1148_),
    .B(_1463_),
    .C(_1468_),
    .Y(_1469_)
);

NAND2X1 _12605_ (
    .A(_1442_),
    .B(_1469_),
    .Y(_1470_)
);

OAI21X1 _12606_ (
    .A(_1440_),
    .B(_1155_),
    .C(_1467_),
    .Y(_1471_)
);

OAI21X1 _12607_ (
    .A(_1764_),
    .B(_1767_),
    .C(_1471_),
    .Y(_1473_)
);

NAND3X1 _12608_ (
    .A(_2133__bF$buf0),
    .B(_1470_),
    .C(_1473_),
    .Y(_1474_)
);

NAND2X1 _12609_ (
    .A(\datapath.alu.b_0_bF$buf9 ),
    .B(_967_),
    .Y(_1475_)
);

OAI21X1 _12610_ (
    .A(\datapath.alu.b_0_bF$buf8 ),
    .B(\datapath.alu.a [24]),
    .C(_1475_),
    .Y(_1476_)
);

NAND2X1 _12611_ (
    .A(_1833__bF$buf6),
    .B(_1476_),
    .Y(_1477_)
);

OAI21X1 _12612_ (
    .A(_1833__bF$buf5),
    .B(_1399_),
    .C(_1477_),
    .Y(_1478_)
);

MUX2X1 _12613_ (
    .A(_1478_),
    .B(_1325_),
    .S(_1839__bF$buf2),
    .Y(_1479_)
);

NAND2X1 _12614_ (
    .A(\datapath.alu.b_3_bF$buf7 ),
    .B(_1175_),
    .Y(_1480_)
);

OAI21X1 _12615_ (
    .A(\datapath.alu.b_3_bF$buf6 ),
    .B(_1479_),
    .C(_1480_),
    .Y(_1481_)
);

AND2X2 _12616_ (
    .A(_2501_),
    .B(_2502_),
    .Y(_1482_)
);

INVX1 _12617_ (
    .A(_1764_),
    .Y(_1484_)
);

AOI21X1 _12618_ (
    .A(_1484_),
    .B(_2027__bF$buf3),
    .C(_1157_),
    .Y(_1485_)
);

INVX1 _12619_ (
    .A(_1767_),
    .Y(_1486_)
);

OAI22X1 _12620_ (
    .A(_1486_),
    .B(_2014__bF$buf0),
    .C(_2047__bF$buf2),
    .D(_1457_),
    .Y(_1487_)
);

AOI22X1 _12621_ (
    .A(_1893_),
    .B(_2016__bF$buf2),
    .C(\datapath.alu.b [24]),
    .D(_2029_),
    .Y(_1488_)
);

OAI21X1 _12622_ (
    .A(_1765_),
    .B(_2118__bF$buf0),
    .C(_1488_),
    .Y(_1489_)
);

NOR2X1 _12623_ (
    .A(_1489_),
    .B(_1487_),
    .Y(_1490_)
);

NAND2X1 _12624_ (
    .A(_1485_),
    .B(_1490_),
    .Y(_1491_)
);

AOI21X1 _12625_ (
    .A(_1482_),
    .B(_1211_),
    .C(_1491_),
    .Y(_1492_)
);

OAI21X1 _12626_ (
    .A(_2127_),
    .B(_1481_),
    .C(_1492_),
    .Y(_1493_)
);

AOI21X1 _12627_ (
    .A(_1824__bF$buf2),
    .B(_2495_),
    .C(_1493_),
    .Y(_1495_)
);

NAND3X1 _12628_ (
    .A(_1495_),
    .B(_1474_),
    .C(_1462_),
    .Y(\datapath.alu.c [24])
);

INVX1 _12629_ (
    .A(_1763_),
    .Y(_1496_)
);

AOI21X1 _12630_ (
    .A(_1459_),
    .B(_1454_),
    .C(_1457_),
    .Y(_1497_)
);

OAI21X1 _12631_ (
    .A(_1767_),
    .B(_1497_),
    .C(_1496_),
    .Y(_1498_)
);

OAI21X1 _12632_ (
    .A(_1447_),
    .B(_1136_),
    .C(_1454_),
    .Y(_1499_)
);

AOI21X1 _12633_ (
    .A(_1499_),
    .B(_1442_),
    .C(_1767_),
    .Y(_1500_)
);

AOI21X1 _12634_ (
    .A(_1500_),
    .B(_1763_),
    .C(_2251__bF$buf3),
    .Y(_1501_)
);

OAI21X1 _12635_ (
    .A(_1765_),
    .B(\datapath.alu.b [24]),
    .C(_1496_),
    .Y(_1502_)
);

AOI21X1 _12636_ (
    .A(_1471_),
    .B(_1457_),
    .C(_1502_),
    .Y(_1503_)
);

NOR2X1 _12637_ (
    .A(\datapath.alu.b [24]),
    .B(_1765_),
    .Y(_1505_)
);

AOI21X1 _12638_ (
    .A(_1763_),
    .B(_1505_),
    .C(_2134_),
    .Y(_1506_)
);

OAI21X1 _12639_ (
    .A(_1768_),
    .B(_1469_),
    .C(_1506_),
    .Y(_1507_)
);

OAI21X1 _12640_ (
    .A(_1841__bF$buf5),
    .B(_2130_),
    .C(_2549_),
    .Y(_1508_)
);

OAI22X1 _12641_ (
    .A(_1763_),
    .B(_2047__bF$buf1),
    .C(_1750_),
    .D(_2014__bF$buf3),
    .Y(_1509_)
);

AOI22X1 _12642_ (
    .A(_1892_),
    .B(_2016__bF$buf1),
    .C(\datapath.alu.b [25]),
    .D(_2029_),
    .Y(_1510_)
);

OAI21X1 _12643_ (
    .A(_1760_),
    .B(_2118__bF$buf3),
    .C(_1510_),
    .Y(_1511_)
);

INVX1 _12644_ (
    .A(_1762_),
    .Y(_1512_)
);

OAI21X1 _12645_ (
    .A(_1512_),
    .B(_2122_),
    .C(_1158_),
    .Y(_1513_)
);

NOR3X1 _12646_ (
    .A(_1509_),
    .B(_1511_),
    .C(_1513_),
    .Y(_1514_)
);

OAI21X1 _12647_ (
    .A(_1508_),
    .B(_1212_),
    .C(_1514_),
    .Y(_1516_)
);

NAND2X1 _12648_ (
    .A(\datapath.alu.b_0_bF$buf7 ),
    .B(_1765_),
    .Y(_1517_)
);

OAI21X1 _12649_ (
    .A(\datapath.alu.b_0_bF$buf6 ),
    .B(\datapath.alu.a [25]),
    .C(_1517_),
    .Y(_1518_)
);

NAND2X1 _12650_ (
    .A(_1833__bF$buf4),
    .B(_1518_),
    .Y(_1519_)
);

OAI21X1 _12651_ (
    .A(_1833__bF$buf3),
    .B(_1422_),
    .C(_1519_),
    .Y(_1520_)
);

NOR2X1 _12652_ (
    .A(\datapath.alu.b_2_bF$buf4 ),
    .B(_1520_),
    .Y(_1521_)
);

OAI21X1 _12653_ (
    .A(_1839__bF$buf1),
    .B(_1356_),
    .C(_1841__bF$buf4),
    .Y(_1522_)
);

NAND3X1 _12654_ (
    .A(\datapath.alu.b_3_bF$buf5 ),
    .B(_1192_),
    .C(_1198_),
    .Y(_1523_)
);

OAI21X1 _12655_ (
    .A(_1521_),
    .B(_1522_),
    .C(_1523_),
    .Y(_1524_)
);

OAI21X1 _12656_ (
    .A(_2039_),
    .B(_1524_),
    .C(_2537_),
    .Y(_1525_)
);

AOI21X1 _12657_ (
    .A(_1525_),
    .B(_1824__bF$buf1),
    .C(_1516_),
    .Y(_1527_)
);

OAI21X1 _12658_ (
    .A(_1507_),
    .B(_1503_),
    .C(_1527_),
    .Y(_1528_)
);

AOI21X1 _12659_ (
    .A(_1501_),
    .B(_1498_),
    .C(_1528_),
    .Y(_1529_)
);

INVX1 _12660_ (
    .A(_1529_),
    .Y(\datapath.alu.c [25])
);

NOR2X1 _12661_ (
    .A(_1763_),
    .B(_1457_),
    .Y(_1530_)
);

OAI21X1 _12662_ (
    .A(_1512_),
    .B(_1486_),
    .C(_1750_),
    .Y(_1531_)
);

AOI21X1 _12663_ (
    .A(_1499_),
    .B(_1530_),
    .C(_1531_),
    .Y(_1532_)
);

AOI21X1 _12664_ (
    .A(_1532_),
    .B(_1729_),
    .C(_2251__bF$buf2),
    .Y(_1533_)
);

OAI21X1 _12665_ (
    .A(_1729_),
    .B(_1532_),
    .C(_1533_),
    .Y(_1534_)
);

INVX1 _12666_ (
    .A(_1750_),
    .Y(_1535_)
);

OAI21X1 _12667_ (
    .A(_1535_),
    .B(_1512_),
    .C(_1505_),
    .Y(_1537_)
);

OAI21X1 _12668_ (
    .A(_1760_),
    .B(\datapath.alu.b [25]),
    .C(_1537_),
    .Y(_1538_)
);

INVX1 _12669_ (
    .A(_1538_),
    .Y(_1539_)
);

OAI21X1 _12670_ (
    .A(_1768_),
    .B(_1469_),
    .C(_1539_),
    .Y(_1540_)
);

AOI21X1 _12671_ (
    .A(_1540_),
    .B(_1729_),
    .C(_2134_),
    .Y(_1541_)
);

OAI21X1 _12672_ (
    .A(_1729_),
    .B(_1540_),
    .C(_1541_),
    .Y(_1542_)
);

NAND2X1 _12673_ (
    .A(\datapath.alu.b_0_bF$buf5 ),
    .B(_1760_),
    .Y(_1543_)
);

OAI21X1 _12674_ (
    .A(\datapath.alu.b_0_bF$buf4 ),
    .B(\datapath.alu.a [26]),
    .C(_1543_),
    .Y(_1544_)
);

INVX1 _12675_ (
    .A(_1544_),
    .Y(_1545_)
);

NAND2X1 _12676_ (
    .A(\datapath.alu.b_1_bF$buf2 ),
    .B(_1476_),
    .Y(_1546_)
);

OAI21X1 _12677_ (
    .A(\datapath.alu.b_1_bF$buf1 ),
    .B(_1545_),
    .C(_1546_),
    .Y(_1548_)
);

NAND2X1 _12678_ (
    .A(_1839__bF$buf0),
    .B(_1548_),
    .Y(_1549_)
);

OAI21X1 _12679_ (
    .A(_1839__bF$buf6),
    .B(_1401_),
    .C(_1549_),
    .Y(_1550_)
);

NOR2X1 _12680_ (
    .A(\datapath.alu.b_3_bF$buf4 ),
    .B(_1550_),
    .Y(_1551_)
);

NOR2X1 _12681_ (
    .A(_1841__bF$buf3),
    .B(_1252_),
    .Y(_1552_)
);

OAI21X1 _12682_ (
    .A(_1552_),
    .B(_1551_),
    .C(_2040_),
    .Y(_1553_)
);

OAI21X1 _12683_ (
    .A(_1841__bF$buf2),
    .B(_2180_),
    .C(_900_),
    .Y(_1554_)
);

OAI21X1 _12684_ (
    .A(\datapath.alu.a [26]),
    .B(_2017_),
    .C(_2267__bF$buf3),
    .Y(_1555_)
);

OAI22X1 _12685_ (
    .A(_1686_),
    .B(_2118__bF$buf2),
    .C(_1729_),
    .D(_2047__bF$buf0),
    .Y(_1556_)
);

OAI21X1 _12686_ (
    .A(\datapath.alu.a [26]),
    .B(\datapath.alu.b [26]),
    .C(_2027__bF$buf2),
    .Y(_1557_)
);

OAI21X1 _12687_ (
    .A(_1718_),
    .B(_2014__bF$buf2),
    .C(_1557_),
    .Y(_1559_)
);

NOR2X1 _12688_ (
    .A(_1556_),
    .B(_1559_),
    .Y(_1560_)
);

OAI21X1 _12689_ (
    .A(_1824__bF$buf0),
    .B(_1108_),
    .C(_1560_),
    .Y(_1561_)
);

AOI21X1 _12690_ (
    .A(\datapath.alu.b [26]),
    .B(_1555_),
    .C(_1561_),
    .Y(_1562_)
);

OAI21X1 _12691_ (
    .A(_1554_),
    .B(_1212_),
    .C(_1562_),
    .Y(_1563_)
);

AOI21X1 _12692_ (
    .A(_1824__bF$buf5),
    .B(_879_),
    .C(_1563_),
    .Y(_1564_)
);

AND2X2 _12693_ (
    .A(_1564_),
    .B(_1553_),
    .Y(_1565_)
);

NAND3X1 _12694_ (
    .A(_1542_),
    .B(_1565_),
    .C(_1534_),
    .Y(\datapath.alu.c [26])
);

NOR2X1 _12695_ (
    .A(_1676_),
    .B(_1665_),
    .Y(_1566_)
);

INVX1 _12696_ (
    .A(_1566_),
    .Y(_1567_)
);

INVX1 _12697_ (
    .A(_1718_),
    .Y(_1569_)
);

OAI21X1 _12698_ (
    .A(_1455_),
    .B(_1448_),
    .C(_1530_),
    .Y(_1570_)
);

INVX1 _12699_ (
    .A(_1531_),
    .Y(_1571_)
);

AOI21X1 _12700_ (
    .A(_1570_),
    .B(_1571_),
    .C(_1729_),
    .Y(_1572_)
);

OAI21X1 _12701_ (
    .A(_1569_),
    .B(_1572_),
    .C(_1567_),
    .Y(_1573_)
);

INVX1 _12702_ (
    .A(_1729_),
    .Y(_1574_)
);

INVX1 _12703_ (
    .A(_1530_),
    .Y(_1575_)
);

AOI21X1 _12704_ (
    .A(_1459_),
    .B(_1454_),
    .C(_1575_),
    .Y(_1576_)
);

OAI21X1 _12705_ (
    .A(_1531_),
    .B(_1576_),
    .C(_1574_),
    .Y(_1577_)
);

NAND3X1 _12706_ (
    .A(_1566_),
    .B(_1718_),
    .C(_1577_),
    .Y(_1578_)
);

AOI21X1 _12707_ (
    .A(_1573_),
    .B(_1578_),
    .C(_2251__bF$buf1),
    .Y(_1580_)
);

NOR2X1 _12708_ (
    .A(\datapath.alu.b [26]),
    .B(_1686_),
    .Y(_1581_)
);

AOI21X1 _12709_ (
    .A(_1540_),
    .B(_1729_),
    .C(_1581_),
    .Y(_1582_)
);

AND2X2 _12710_ (
    .A(_1582_),
    .B(_1566_),
    .Y(_1583_)
);

OAI21X1 _12711_ (
    .A(_1566_),
    .B(_1582_),
    .C(_2133__bF$buf3),
    .Y(_1584_)
);

NOR2X1 _12712_ (
    .A(_1841__bF$buf1),
    .B(_1288_),
    .Y(_1585_)
);

NAND2X1 _12713_ (
    .A(\datapath.alu.b_0_bF$buf3 ),
    .B(_1686_),
    .Y(_1586_)
);

OAI21X1 _12714_ (
    .A(\datapath.alu.b_0_bF$buf2 ),
    .B(\datapath.alu.a [27]),
    .C(_1586_),
    .Y(_1587_)
);

MUX2X1 _12715_ (
    .A(_1587_),
    .B(_1518_),
    .S(_1833__bF$buf2),
    .Y(_1588_)
);

MUX2X1 _12716_ (
    .A(_1588_),
    .B(_1424_),
    .S(_1839__bF$buf5),
    .Y(_1589_)
);

NOR2X1 _12717_ (
    .A(\datapath.alu.b_3_bF$buf3 ),
    .B(_1589_),
    .Y(_1591_)
);

OAI21X1 _12718_ (
    .A(_1591_),
    .B(_1585_),
    .C(_2040_),
    .Y(_1592_)
);

NAND2X1 _12719_ (
    .A(_1211_),
    .B(_936_),
    .Y(_1593_)
);

OAI21X1 _12720_ (
    .A(\datapath.alu.a [27]),
    .B(_2017_),
    .C(_2267__bF$buf2),
    .Y(_1594_)
);

AOI22X1 _12721_ (
    .A(_1665_),
    .B(_2197_),
    .C(_2553_),
    .D(_1566_),
    .Y(_1595_)
);

OAI21X1 _12722_ (
    .A(_1676_),
    .B(_2122_),
    .C(_1595_),
    .Y(_1596_)
);

OAI21X1 _12723_ (
    .A(_1643_),
    .B(_2118__bF$buf1),
    .C(_1158_),
    .Y(_1597_)
);

OR2X2 _12724_ (
    .A(_1597_),
    .B(_1596_),
    .Y(_1598_)
);

AOI21X1 _12725_ (
    .A(\datapath.alu.b [27]),
    .B(_1594_),
    .C(_1598_),
    .Y(_1599_)
);

NAND3X1 _12726_ (
    .A(_1592_),
    .B(_1593_),
    .C(_1599_),
    .Y(_1600_)
);

AOI21X1 _12727_ (
    .A(_1824__bF$buf4),
    .B(_926_),
    .C(_1600_),
    .Y(_1602_)
);

OAI21X1 _12728_ (
    .A(_1583_),
    .B(_1584_),
    .C(_1602_),
    .Y(_1603_)
);

OR2X2 _12729_ (
    .A(_1603_),
    .B(_1580_),
    .Y(\datapath.alu.c [27])
);

NOR2X1 _12730_ (
    .A(_1729_),
    .B(_1567_),
    .Y(_1604_)
);

INVX1 _12731_ (
    .A(_1604_),
    .Y(_1605_)
);

NOR2X1 _12732_ (
    .A(_1605_),
    .B(_1575_),
    .Y(_1606_)
);

AOI21X1 _12733_ (
    .A(_1566_),
    .B(_1569_),
    .C(_1665_),
    .Y(_1607_)
);

OAI21X1 _12734_ (
    .A(_1571_),
    .B(_1605_),
    .C(_1607_),
    .Y(_1608_)
);

AOI21X1 _12735_ (
    .A(_1499_),
    .B(_1606_),
    .C(_1608_),
    .Y(_1609_)
);

AOI21X1 _12736_ (
    .A(_1609_),
    .B(_1611_),
    .C(_2251__bF$buf0),
    .Y(_1610_)
);

OAI21X1 _12737_ (
    .A(_1611_),
    .B(_1609_),
    .C(_1610_),
    .Y(_1612_)
);

INVX1 _12738_ (
    .A(_1769_),
    .Y(_1613_)
);

INVX1 _12739_ (
    .A(_1740_),
    .Y(_1614_)
);

INVX1 _12740_ (
    .A(_1581_),
    .Y(_1615_)
);

OAI21X1 _12741_ (
    .A(_1897_),
    .B(_1615_),
    .C(_1895_),
    .Y(_1616_)
);

AOI21X1 _12742_ (
    .A(_1538_),
    .B(_1614_),
    .C(_1616_),
    .Y(_1617_)
);

OAI21X1 _12743_ (
    .A(_1613_),
    .B(_1469_),
    .C(_1617_),
    .Y(_1618_)
);

AOI21X1 _12744_ (
    .A(_1618_),
    .B(_1611_),
    .C(_2134_),
    .Y(_1619_)
);

OAI21X1 _12745_ (
    .A(_1611_),
    .B(_1618_),
    .C(_1619_),
    .Y(_1620_)
);

NAND2X1 _12746_ (
    .A(_992_),
    .B(_991_),
    .Y(_1621_)
);

OAI21X1 _12747_ (
    .A(\datapath.alu.a [28]),
    .B(_2017_),
    .C(_2267__bF$buf1),
    .Y(_1623_)
);

OAI21X1 _12748_ (
    .A(\datapath.alu.a [28]),
    .B(\datapath.alu.b [28]),
    .C(_2027__bF$buf1),
    .Y(_1624_)
);

INVX1 _12749_ (
    .A(_1601_),
    .Y(_1625_)
);

INVX1 _12750_ (
    .A(_1611_),
    .Y(_1626_)
);

AOI22X1 _12751_ (
    .A(_1625_),
    .B(_2197_),
    .C(_2553_),
    .D(_1626_),
    .Y(_1627_)
);

NAND3X1 _12752_ (
    .A(_1624_),
    .B(_1627_),
    .C(_1158_),
    .Y(_1628_)
);

AOI21X1 _12753_ (
    .A(\datapath.alu.b [28]),
    .B(_1623_),
    .C(_1628_),
    .Y(_1629_)
);

OAI21X1 _12754_ (
    .A(_1568_),
    .B(_2118__bF$buf0),
    .C(_1629_),
    .Y(_1630_)
);

MUX2X1 _12755_ (
    .A(_1643_),
    .B(_1568_),
    .S(\datapath.alu.b_0_bF$buf1 ),
    .Y(_1631_)
);

NAND2X1 _12756_ (
    .A(\datapath.alu.b_1_bF$buf0 ),
    .B(_1544_),
    .Y(_1632_)
);

OAI21X1 _12757_ (
    .A(\datapath.alu.b_1_bF$buf6 ),
    .B(_1631_),
    .C(_1632_),
    .Y(_1634_)
);

MUX2X1 _12758_ (
    .A(_1634_),
    .B(_1478_),
    .S(_1839__bF$buf4),
    .Y(_1635_)
);

MUX2X1 _12759_ (
    .A(_1635_),
    .B(_1326_),
    .S(_1841__bF$buf0),
    .Y(_1636_)
);

AOI22X1 _12760_ (
    .A(_2127_),
    .B(_986_),
    .C(_1824__bF$buf3),
    .D(_1636_),
    .Y(_1637_)
);

OR2X2 _12761_ (
    .A(_1630_),
    .B(_1637_),
    .Y(_1638_)
);

AOI21X1 _12762_ (
    .A(_1824__bF$buf2),
    .B(_1621_),
    .C(_1638_),
    .Y(_1639_)
);

NAND3X1 _12763_ (
    .A(_1620_),
    .B(_1639_),
    .C(_1612_),
    .Y(\datapath.alu.c [28])
);

INVX1 _12764_ (
    .A(_1606_),
    .Y(_1640_)
);

AOI21X1 _12765_ (
    .A(_1459_),
    .B(_1454_),
    .C(_1640_),
    .Y(_1641_)
);

OAI21X1 _12766_ (
    .A(_1608_),
    .B(_1641_),
    .C(_1626_),
    .Y(_1642_)
);

AOI21X1 _12767_ (
    .A(_1642_),
    .B(_1601_),
    .C(_1558_),
    .Y(_1644_)
);

INVX1 _12768_ (
    .A(_1558_),
    .Y(_1645_)
);

OAI21X1 _12769_ (
    .A(_1611_),
    .B(_1609_),
    .C(_1601_),
    .Y(_1646_)
);

OAI21X1 _12770_ (
    .A(_1645_),
    .B(_1646_),
    .C(_2045_),
    .Y(_1647_)
);

NAND2X1 _12771_ (
    .A(_1611_),
    .B(_1618_),
    .Y(_1648_)
);

NOR2X1 _12772_ (
    .A(\datapath.alu.b [28]),
    .B(_1568_),
    .Y(_1649_)
);

NOR2X1 _12773_ (
    .A(_1649_),
    .B(_1558_),
    .Y(_1650_)
);

NAND2X1 _12774_ (
    .A(_1650_),
    .B(_1648_),
    .Y(_1651_)
);

INVX1 _12775_ (
    .A(_1622_),
    .Y(_1652_)
);

NAND2X1 _12776_ (
    .A(_1649_),
    .B(_1558_),
    .Y(_1653_)
);

NAND2X1 _12777_ (
    .A(_2133__bF$buf2),
    .B(_1653_),
    .Y(_1655_)
);

AOI21X1 _12778_ (
    .A(_1618_),
    .B(_1652_),
    .C(_1655_),
    .Y(_1656_)
);

AOI22X1 _12779_ (
    .A(_1900_),
    .B(_2016__bF$buf0),
    .C(\datapath.alu.b [29]),
    .D(_2029_),
    .Y(_1657_)
);

OAI22X1 _12780_ (
    .A(_1558_),
    .B(_2047__bF$buf3),
    .C(_1515_),
    .D(_2014__bF$buf1),
    .Y(_1658_)
);

OAI21X1 _12781_ (
    .A(\datapath.alu.a [29]),
    .B(\datapath.alu.b [29]),
    .C(_2027__bF$buf0),
    .Y(_1659_)
);

OAI21X1 _12782_ (
    .A(_1526_),
    .B(_2118__bF$buf3),
    .C(_1659_),
    .Y(_1660_)
);

NOR2X1 _12783_ (
    .A(_1658_),
    .B(_1660_),
    .Y(_1661_)
);

NAND3X1 _12784_ (
    .A(_1158_),
    .B(_1657_),
    .C(_1661_),
    .Y(_1662_)
);

AOI21X1 _12785_ (
    .A(_1015_),
    .B(_1824__bF$buf1),
    .C(_1662_),
    .Y(_1663_)
);

OAI21X1 _12786_ (
    .A(\datapath.alu.b_0_bF$buf0 ),
    .B(_1526_),
    .C(_2070_),
    .Y(_1664_)
);

NAND2X1 _12787_ (
    .A(\datapath.alu.b_1_bF$buf5 ),
    .B(_1587_),
    .Y(_1666_)
);

OAI21X1 _12788_ (
    .A(\datapath.alu.b_1_bF$buf4 ),
    .B(_1664_),
    .C(_1666_),
    .Y(_1667_)
);

MUX2X1 _12789_ (
    .A(_1520_),
    .B(_1667_),
    .S(\datapath.alu.b_2_bF$buf3 ),
    .Y(_1668_)
);

NOR2X1 _12790_ (
    .A(\datapath.alu.b_3_bF$buf2 ),
    .B(_1668_),
    .Y(_1669_)
);

NOR2X1 _12791_ (
    .A(_1841__bF$buf7),
    .B(_1357_),
    .Y(_1670_)
);

OAI21X1 _12792_ (
    .A(_1670_),
    .B(_1669_),
    .C(_1824__bF$buf0),
    .Y(_1671_)
);

NAND2X1 _12793_ (
    .A(\datapath.alu.b_4_bF$buf0 ),
    .B(_1037_),
    .Y(_1672_)
);

NAND2X1 _12794_ (
    .A(_1671_),
    .B(_1672_),
    .Y(_1673_)
);

OAI21X1 _12795_ (
    .A(_2039_),
    .B(_1673_),
    .C(_1663_),
    .Y(_1674_)
);

AOI21X1 _12796_ (
    .A(_1651_),
    .B(_1656_),
    .C(_1674_),
    .Y(_1675_)
);

OAI21X1 _12797_ (
    .A(_1644_),
    .B(_1647_),
    .C(_1675_),
    .Y(\datapath.alu.c [29])
);

INVX2 _12798_ (
    .A(_1494_),
    .Y(_1677_)
);

INVX1 _12799_ (
    .A(_1515_),
    .Y(_1678_)
);

AOI21X1 _12800_ (
    .A(_1547_),
    .B(_1625_),
    .C(_1678_),
    .Y(_1679_)
);

NOR2X1 _12801_ (
    .A(_1558_),
    .B(_1611_),
    .Y(_1680_)
);

OAI21X1 _12802_ (
    .A(_1608_),
    .B(_1641_),
    .C(_1680_),
    .Y(_1681_)
);

NAND2X1 _12803_ (
    .A(_1679_),
    .B(_1681_),
    .Y(_1682_)
);

NAND2X1 _12804_ (
    .A(_1677_),
    .B(_1682_),
    .Y(_1683_)
);

AND2X2 _12805_ (
    .A(_1681_),
    .B(_1679_),
    .Y(_1684_)
);

AOI21X1 _12806_ (
    .A(_1684_),
    .B(_1494_),
    .C(_2251__bF$buf3),
    .Y(_1685_)
);

OAI21X1 _12807_ (
    .A(_1526_),
    .B(\datapath.alu.b [29]),
    .C(_1653_),
    .Y(_1687_)
);

AOI21X1 _12808_ (
    .A(_1618_),
    .B(_1652_),
    .C(_1687_),
    .Y(_1688_)
);

AND2X2 _12809_ (
    .A(_1688_),
    .B(_1677_),
    .Y(_1689_)
);

OAI21X1 _12810_ (
    .A(_1677_),
    .B(_1688_),
    .C(_2133__bF$buf1),
    .Y(_1690_)
);

OAI21X1 _12811_ (
    .A(\datapath.alu.a [30]),
    .B(_2017_),
    .C(_2267__bF$buf0),
    .Y(_1691_)
);

NAND2X1 _12812_ (
    .A(\datapath.alu.a [30]),
    .B(_2022_),
    .Y(_1692_)
);

OAI21X1 _12813_ (
    .A(_1494_),
    .B(_2047__bF$buf2),
    .C(_1692_),
    .Y(_1693_)
);

OAI21X1 _12814_ (
    .A(\datapath.alu.a [30]),
    .B(\datapath.alu.b [30]),
    .C(_2027__bF$buf3),
    .Y(_1694_)
);

OAI21X1 _12815_ (
    .A(_1483_),
    .B(_2014__bF$buf0),
    .C(_1694_),
    .Y(_1695_)
);

NOR2X1 _12816_ (
    .A(_1693_),
    .B(_1695_),
    .Y(_1696_)
);

OAI21X1 _12817_ (
    .A(_1824__bF$buf5),
    .B(_1108_),
    .C(_1696_),
    .Y(_1698_)
);

AOI21X1 _12818_ (
    .A(\datapath.alu.b [30]),
    .B(_1691_),
    .C(_1698_),
    .Y(_1699_)
);

OAI21X1 _12819_ (
    .A(\datapath.alu.b_4_bF$buf4 ),
    .B(_1074_),
    .C(_1699_),
    .Y(_1700_)
);

MUX2X1 _12820_ (
    .A(_1526_),
    .B(_1450_),
    .S(\datapath.alu.b_0_bF$buf9 ),
    .Y(_1701_)
);

MUX2X1 _12821_ (
    .A(_1701_),
    .B(_1631_),
    .S(_1833__bF$buf1),
    .Y(_1702_)
);

MUX2X1 _12822_ (
    .A(_1548_),
    .B(_1702_),
    .S(\datapath.alu.b_2_bF$buf2 ),
    .Y(_1703_)
);

NAND2X1 _12823_ (
    .A(\datapath.alu.b_3_bF$buf1 ),
    .B(_1403_),
    .Y(_1704_)
);

OAI21X1 _12824_ (
    .A(\datapath.alu.b_3_bF$buf0 ),
    .B(_1703_),
    .C(_1704_),
    .Y(_1705_)
);

AOI22X1 _12825_ (
    .A(_2127_),
    .B(_1066_),
    .C(_1824__bF$buf4),
    .D(_1705_),
    .Y(_1706_)
);

NOR2X1 _12826_ (
    .A(_1700_),
    .B(_1706_),
    .Y(_1707_)
);

OAI21X1 _12827_ (
    .A(_1689_),
    .B(_1690_),
    .C(_1707_),
    .Y(_1709_)
);

AOI21X1 _12828_ (
    .A(_1685_),
    .B(_1683_),
    .C(_1709_),
    .Y(_1710_)
);

INVX1 _12829_ (
    .A(_1710_),
    .Y(\datapath.alu.c [30])
);

INVX1 _12830_ (
    .A(_946_),
    .Y(_1711_)
);

INVX1 _12831_ (
    .A(_1483_),
    .Y(_1712_)
);

AOI21X1 _12832_ (
    .A(_1681_),
    .B(_1679_),
    .C(_1494_),
    .Y(_1713_)
);

OAI21X1 _12833_ (
    .A(_1712_),
    .B(_1713_),
    .C(_1711_),
    .Y(_1714_)
);

NAND3X1 _12834_ (
    .A(_946_),
    .B(_1483_),
    .C(_1683_),
    .Y(_1715_)
);

NAND3X1 _12835_ (
    .A(_2045_),
    .B(_1714_),
    .C(_1715_),
    .Y(_1716_)
);

NOR2X1 _12836_ (
    .A(\datapath.alu.b [30]),
    .B(_1450_),
    .Y(_1717_)
);

INVX1 _12837_ (
    .A(_1717_),
    .Y(_1719_)
);

OAI21X1 _12838_ (
    .A(_1677_),
    .B(_1688_),
    .C(_1719_),
    .Y(_1720_)
);

AOI21X1 _12839_ (
    .A(_1720_),
    .B(_946_),
    .C(_2134_),
    .Y(_1721_)
);

OAI21X1 _12840_ (
    .A(_946_),
    .B(_1720_),
    .C(_1721_),
    .Y(_1722_)
);

OAI21X1 _12841_ (
    .A(\datapath.alu.b_1_bF$buf3 ),
    .B(_2076_),
    .C(_2242_),
    .Y(_1723_)
);

AOI21X1 _12842_ (
    .A(\datapath.alu.b_1_bF$buf2 ),
    .B(_1664_),
    .C(_1723_),
    .Y(_1724_)
);

NAND2X1 _12843_ (
    .A(_1839__bF$buf3),
    .B(_1724_),
    .Y(_1725_)
);

OAI21X1 _12844_ (
    .A(_1839__bF$buf2),
    .B(_1588_),
    .C(_1725_),
    .Y(_1726_)
);

MUX2X1 _12845_ (
    .A(_1726_),
    .B(_1425_),
    .S(_1841__bF$buf6),
    .Y(_1727_)
);

INVX1 _12846_ (
    .A(_935_),
    .Y(_1728_)
);

AOI21X1 _12847_ (
    .A(_2553_),
    .B(_903_),
    .C(_2027__bF$buf2),
    .Y(_1730_)
);

OAI22X1 _12848_ (
    .A(_924_),
    .B(_2267__bF$buf3),
    .C(_903_),
    .D(_2014__bF$buf3),
    .Y(_1731_)
);

AOI21X1 _12849_ (
    .A(_1903_),
    .B(_2016__bF$buf3),
    .C(_1731_),
    .Y(_1732_)
);

OAI21X1 _12850_ (
    .A(_1728_),
    .B(_1730_),
    .C(_1732_),
    .Y(_1733_)
);

OAI21X1 _12851_ (
    .A(_2054_),
    .B(_2022_),
    .C(\datapath.alu.a [31]),
    .Y(_1734_)
);

NAND2X1 _12852_ (
    .A(_2025_),
    .B(_1975_),
    .Y(_1735_)
);

OAI21X1 _12853_ (
    .A(_1109_),
    .B(_1735_),
    .C(_1734_),
    .Y(_1736_)
);

NOR2X1 _12854_ (
    .A(_1733_),
    .B(_1736_),
    .Y(_1737_)
);

OAI21X1 _12855_ (
    .A(_1105_),
    .B(_1212_),
    .C(_1737_),
    .Y(_1738_)
);

AOI21X1 _12856_ (
    .A(_2040_),
    .B(_1727_),
    .C(_1738_),
    .Y(_1739_)
);

NAND3X1 _12857_ (
    .A(_1722_),
    .B(_1739_),
    .C(_1716_),
    .Y(\datapath.alu.c [31])
);

NOR3X1 _12858_ (
    .A(_1580_),
    .B(_1603_),
    .C(\datapath.alu.c [29]),
    .Y(_1741_)
);

NAND3X1 _12859_ (
    .A(_1378_),
    .B(_1410_),
    .C(_1529_),
    .Y(_1742_)
);

NOR3X1 _12860_ (
    .A(\datapath.alu.c [26]),
    .B(\datapath.alu.c [28]),
    .C(_1742_),
    .Y(_1743_)
);

NOR2X1 _12861_ (
    .A(\datapath.alu.c [5]),
    .B(\datapath.alu.c [8]),
    .Y(_1744_)
);

NAND3X1 _12862_ (
    .A(_2427_),
    .B(_2053_),
    .C(_1744_),
    .Y(_1745_)
);

NOR3X1 _12863_ (
    .A(\datapath.alu.c [4]),
    .B(\datapath.alu.c [2]),
    .C(\datapath.alu.c [3]),
    .Y(_1746_)
);

NAND3X1 _12864_ (
    .A(_2141_),
    .B(_2472_),
    .C(_1746_),
    .Y(_1747_)
);

NOR2X1 _12865_ (
    .A(_1745_),
    .B(_1747_),
    .Y(_1748_)
);

NAND3X1 _12866_ (
    .A(_907_),
    .B(_1003_),
    .C(_1184_),
    .Y(_1749_)
);

NOR2X1 _12867_ (
    .A(\datapath.alu.c [9]),
    .B(_1749_),
    .Y(_1751_)
);

NAND3X1 _12868_ (
    .A(_1041_),
    .B(_1751_),
    .C(_1748_),
    .Y(_1752_)
);

NOR2X1 _12869_ (
    .A(\datapath.alu.c [24]),
    .B(\datapath.alu.c [20]),
    .Y(_1753_)
);

NAND3X1 _12870_ (
    .A(_1372_),
    .B(_1753_),
    .C(_1260_),
    .Y(_1754_)
);

NOR2X1 _12871_ (
    .A(_1754_),
    .B(_1752_),
    .Y(_1755_)
);

NAND3X1 _12872_ (
    .A(_1743_),
    .B(_1741_),
    .C(_1755_),
    .Y(_1756_)
);

NAND3X1 _12873_ (
    .A(_947_),
    .B(_1088_),
    .C(_1217_),
    .Y(_1757_)
);

NOR3X1 _12874_ (
    .A(\datapath.alu.c [19]),
    .B(\datapath.alu.c [15]),
    .C(_1757_),
    .Y(_1758_)
);

NAND3X1 _12875_ (
    .A(_1441_),
    .B(_1710_),
    .C(_1758_),
    .Y(_1759_)
);

NOR3X1 _12876_ (
    .A(\datapath.alu.c [31]),
    .B(_1759_),
    .C(_1756_),
    .Y(\datapath.alu.z )
);

NAND3X1 _12877_ (
    .A(\datapath.csr.mip ),
    .B(\datapath.csr.mstatus [0]),
    .C(\datapath.csr.mie ),
    .Y(_2575_)
);

INVX1 _12878_ (
    .A(_2575_),
    .Y(\datapath.csr.csr_irq )
);

INVX2 _12879_ (
    .A(\datapath.csr.mvect [0]),
    .Y(_2576_)
);

OAI21X1 _12880_ (
    .A(_2576_),
    .B(_2575_),
    .C(\datapath.csr.mvect [2]),
    .Y(_2577_)
);

INVX1 _12881_ (
    .A(\datapath.csr.mvect [2]),
    .Y(_2578_)
);

NOR2X1 _12882_ (
    .A(_2576_),
    .B(_2575_),
    .Y(_2579_)
);

NAND2X1 _12883_ (
    .A(_2578_),
    .B(_2579_),
    .Y(_2580_)
);

AND2X2 _12884_ (
    .A(_2580_),
    .B(_2577_),
    .Y(_2581_)
);

NAND2X1 _12885_ (
    .A(\datapath.csr.mepc [0]),
    .B(\controlunit.mret_bF$buf3 ),
    .Y(_2582_)
);

OAI21X1 _12886_ (
    .A(\controlunit.mret_bF$buf2 ),
    .B(_2581_),
    .C(_2582_),
    .Y(\datapath.csr.csr_pcaddr [2])
);

INVX1 _12887_ (
    .A(\datapath.csr.mvect [3]),
    .Y(_2583_)
);

XNOR2X1 _12888_ (
    .A(_2580_),
    .B(_2583_),
    .Y(_2584_)
);

NAND2X1 _12889_ (
    .A(\controlunit.mret_bF$buf1 ),
    .B(\datapath.csr.mepc [1]),
    .Y(_2585_)
);

OAI21X1 _12890_ (
    .A(\controlunit.mret_bF$buf0 ),
    .B(_2584_),
    .C(_2585_),
    .Y(\datapath.csr.csr_pcaddr [3])
);

INVX1 _12891_ (
    .A(_2579_),
    .Y(_2586_)
);

INVX1 _12892_ (
    .A(\datapath.csr.mvect [4]),
    .Y(_2587_)
);

NOR2X1 _12893_ (
    .A(\datapath.csr.mvect [2]),
    .B(\datapath.csr.mvect [3]),
    .Y(_2588_)
);

OAI21X1 _12894_ (
    .A(_2588_),
    .B(_2586_),
    .C(_2587_),
    .Y(_2589_)
);

OAI21X1 _12895_ (
    .A(\datapath.csr.mvect [2]),
    .B(\datapath.csr.mvect [3]),
    .C(\datapath.csr.mvect [4]),
    .Y(_2590_)
);

OAI21X1 _12896_ (
    .A(_2586_),
    .B(_2590_),
    .C(_2589_),
    .Y(_2591_)
);

NAND2X1 _12897_ (
    .A(\controlunit.mret_bF$buf4 ),
    .B(\datapath.csr.mepc [2]),
    .Y(_2592_)
);

OAI21X1 _12898_ (
    .A(\controlunit.mret_bF$buf3 ),
    .B(_2591_),
    .C(_2592_),
    .Y(\datapath.csr.csr_pcaddr [4])
);

INVX2 _12899_ (
    .A(\datapath.csr.mvect [5]),
    .Y(_2593_)
);

OAI21X1 _12900_ (
    .A(_2587_),
    .B(_2588_),
    .C(_2579_),
    .Y(_2594_)
);

XNOR2X1 _12901_ (
    .A(_2594_),
    .B(_2593_),
    .Y(_2595_)
);

NAND2X1 _12902_ (
    .A(\controlunit.mret_bF$buf2 ),
    .B(\datapath.csr.mepc [3]),
    .Y(_2596_)
);

OAI21X1 _12903_ (
    .A(\controlunit.mret_bF$buf1 ),
    .B(_2595_),
    .C(_2596_),
    .Y(\datapath.csr.csr_pcaddr [5])
);

INVX8 _12904_ (
    .A(\controlunit.mret_bF$buf0 ),
    .Y(_2597_)
);

INVX1 _12905_ (
    .A(\datapath.csr.mepc [4]),
    .Y(_2598_)
);

NAND2X1 _12906_ (
    .A(_2593_),
    .B(_2590_),
    .Y(_2599_)
);

AOI21X1 _12907_ (
    .A(_2579_),
    .B(_2599_),
    .C(\datapath.csr.mvect [6]),
    .Y(_2600_)
);

INVX1 _12908_ (
    .A(\datapath.csr.mvect [6]),
    .Y(_2601_)
);

NAND2X1 _12909_ (
    .A(_2599_),
    .B(_2579_),
    .Y(_2602_)
);

OAI21X1 _12910_ (
    .A(_2601_),
    .B(_2602_),
    .C(_2597__bF$buf5),
    .Y(_2603_)
);

OAI22X1 _12911_ (
    .A(_2597__bF$buf4),
    .B(_2598_),
    .C(_2600_),
    .D(_2603_),
    .Y(\datapath.csr.csr_pcaddr [6])
);

INVX1 _12912_ (
    .A(\datapath.csr.mepc [5]),
    .Y(_2604_)
);

INVX1 _12913_ (
    .A(\datapath.csr.mvect [7]),
    .Y(_2605_)
);

OAI21X1 _12914_ (
    .A(_2601_),
    .B(_2602_),
    .C(_2605_),
    .Y(_2606_)
);

NAND2X1 _12915_ (
    .A(\datapath.csr.mvect [6]),
    .B(\datapath.csr.mvect [7]),
    .Y(_2607_)
);

INVX1 _12916_ (
    .A(_2607_),
    .Y(_2608_)
);

NAND3X1 _12917_ (
    .A(_2608_),
    .B(_2599_),
    .C(_2579_),
    .Y(_2609_)
);

NAND3X1 _12918_ (
    .A(_2597__bF$buf3),
    .B(_2609_),
    .C(_2606_),
    .Y(_2610_)
);

OAI21X1 _12919_ (
    .A(_2597__bF$buf2),
    .B(_2604_),
    .C(_2610_),
    .Y(\datapath.csr.csr_pcaddr [7])
);

INVX1 _12920_ (
    .A(\datapath.csr.mepc [6]),
    .Y(_2611_)
);

AOI21X1 _12921_ (
    .A(_2590_),
    .B(_2593_),
    .C(_2607_),
    .Y(_2612_)
);

AND2X2 _12922_ (
    .A(_2612_),
    .B(_2579_),
    .Y(_2613_)
);

NAND2X1 _12923_ (
    .A(\datapath.csr.mvect [8]),
    .B(_2613_),
    .Y(_2614_)
);

INVX1 _12924_ (
    .A(_2614_),
    .Y(_2615_)
);

OAI21X1 _12925_ (
    .A(\datapath.csr.mvect [8]),
    .B(_2613_),
    .C(_2597__bF$buf1),
    .Y(_2616_)
);

OAI22X1 _12926_ (
    .A(_2597__bF$buf0),
    .B(_2611_),
    .C(_2616_),
    .D(_2615_),
    .Y(\datapath.csr.csr_pcaddr [8])
);

INVX1 _12927_ (
    .A(\datapath.csr.mepc [7]),
    .Y(_2617_)
);

NAND2X1 _12928_ (
    .A(\datapath.csr.mvect [8]),
    .B(\datapath.csr.mvect [9]),
    .Y(_2618_)
);

INVX1 _12929_ (
    .A(_2618_),
    .Y(_2619_)
);

AOI21X1 _12930_ (
    .A(_2613_),
    .B(_2619_),
    .C(\controlunit.mret_bF$buf4 ),
    .Y(_2620_)
);

OAI21X1 _12931_ (
    .A(\datapath.csr.mvect [9]),
    .B(_2615_),
    .C(_2620_),
    .Y(_2621_)
);

OAI21X1 _12932_ (
    .A(_2597__bF$buf5),
    .B(_2617_),
    .C(_2621_),
    .Y(\datapath.csr.csr_pcaddr [9])
);

INVX1 _12933_ (
    .A(\datapath.csr.mvect [10]),
    .Y(_2622_)
);

INVX1 _12934_ (
    .A(\datapath.csr.mepc [8]),
    .Y(_2623_)
);

NAND2X1 _12935_ (
    .A(\controlunit.mret_bF$buf3 ),
    .B(_2623_),
    .Y(_2624_)
);

NAND2X1 _12936_ (
    .A(\datapath.csr.mvect [10]),
    .B(_2619_),
    .Y(_2625_)
);

INVX1 _12937_ (
    .A(_2625_),
    .Y(_2626_)
);

NAND2X1 _12938_ (
    .A(_2626_),
    .B(_2613_),
    .Y(_2627_)
);

OAI21X1 _12939_ (
    .A(\controlunit.mret_bF$buf2 ),
    .B(_2627_),
    .C(_2624_),
    .Y(_2628_)
);

AOI21X1 _12940_ (
    .A(_2622_),
    .B(_2620_),
    .C(_2628_),
    .Y(\datapath.csr.csr_pcaddr [10])
);

INVX1 _12941_ (
    .A(_2627_),
    .Y(_2629_)
);

NAND2X1 _12942_ (
    .A(\datapath.csr.mvect [10]),
    .B(\datapath.csr.mvect [11]),
    .Y(_2630_)
);

NOR2X1 _12943_ (
    .A(_2618_),
    .B(_2630_),
    .Y(_2631_)
);

NAND3X1 _12944_ (
    .A(_2579_),
    .B(_2631_),
    .C(_2612_),
    .Y(_2632_)
);

OAI21X1 _12945_ (
    .A(\datapath.csr.mvect [11]),
    .B(_2629_),
    .C(_2632_),
    .Y(_2633_)
);

NAND2X1 _12946_ (
    .A(\controlunit.mret_bF$buf1 ),
    .B(\datapath.csr.mepc [9]),
    .Y(_2634_)
);

OAI21X1 _12947_ (
    .A(\controlunit.mret_bF$buf0 ),
    .B(_2633_),
    .C(_2634_),
    .Y(\datapath.csr.csr_pcaddr [11])
);

INVX2 _12948_ (
    .A(\datapath.csr.mvect [12]),
    .Y(_2635_)
);

XNOR2X1 _12949_ (
    .A(_2632_),
    .B(_2635_),
    .Y(_2636_)
);

NAND2X1 _12950_ (
    .A(\controlunit.mret_bF$buf4 ),
    .B(\datapath.csr.mepc [10]),
    .Y(_2637_)
);

OAI21X1 _12951_ (
    .A(\controlunit.mret_bF$buf3 ),
    .B(_2636_),
    .C(_2637_),
    .Y(\datapath.csr.csr_pcaddr [12])
);

INVX1 _12952_ (
    .A(\datapath.csr.mepc [11]),
    .Y(_2638_)
);

INVX1 _12953_ (
    .A(\datapath.csr.mvect [13]),
    .Y(_2639_)
);

OAI21X1 _12954_ (
    .A(_2635_),
    .B(_2632_),
    .C(_2639_),
    .Y(_2640_)
);

INVX1 _12955_ (
    .A(_2640_),
    .Y(_2641_)
);

NAND2X1 _12956_ (
    .A(\datapath.csr.mvect [12]),
    .B(\datapath.csr.mvect [13]),
    .Y(_2642_)
);

OAI21X1 _12957_ (
    .A(_2642_),
    .B(_2632_),
    .C(_2597__bF$buf4),
    .Y(_2643_)
);

OAI22X1 _12958_ (
    .A(_2597__bF$buf3),
    .B(_2638_),
    .C(_2643_),
    .D(_2641_),
    .Y(\datapath.csr.csr_pcaddr [13])
);

INVX1 _12959_ (
    .A(\datapath.csr.mepc [12]),
    .Y(_2644_)
);

INVX1 _12960_ (
    .A(\datapath.csr.mvect [14]),
    .Y(_2645_)
);

OAI21X1 _12961_ (
    .A(_2642_),
    .B(_2632_),
    .C(_2645_),
    .Y(_2646_)
);

INVX1 _12962_ (
    .A(_2632_),
    .Y(_2647_)
);

INVX1 _12963_ (
    .A(_2642_),
    .Y(_2648_)
);

NAND3X1 _12964_ (
    .A(\datapath.csr.mvect [14]),
    .B(_2648_),
    .C(_2647_),
    .Y(_2649_)
);

NAND3X1 _12965_ (
    .A(_2597__bF$buf2),
    .B(_2646_),
    .C(_2649_),
    .Y(_2650_)
);

OAI21X1 _12966_ (
    .A(_2597__bF$buf1),
    .B(_2644_),
    .C(_2650_),
    .Y(\datapath.csr.csr_pcaddr [14])
);

INVX1 _12967_ (
    .A(\datapath.csr.mepc [13]),
    .Y(_2651_)
);

INVX1 _12968_ (
    .A(\datapath.csr.mvect [15]),
    .Y(_2652_)
);

NAND2X1 _12969_ (
    .A(_2652_),
    .B(_2649_),
    .Y(_2653_)
);

INVX1 _12970_ (
    .A(_2653_),
    .Y(_2654_)
);

NAND2X1 _12971_ (
    .A(\datapath.csr.mvect [14]),
    .B(\datapath.csr.mvect [15]),
    .Y(_2655_)
);

NOR2X1 _12972_ (
    .A(_2642_),
    .B(_2655_),
    .Y(_2656_)
);

INVX1 _12973_ (
    .A(_2656_),
    .Y(_2657_)
);

OAI21X1 _12974_ (
    .A(_2657_),
    .B(_2632_),
    .C(_2597__bF$buf0),
    .Y(_2658_)
);

OAI22X1 _12975_ (
    .A(_2597__bF$buf5),
    .B(_2651_),
    .C(_2658_),
    .D(_2654_),
    .Y(\datapath.csr.csr_pcaddr [15])
);

INVX1 _12976_ (
    .A(\datapath.csr.mepc [14]),
    .Y(_2659_)
);

NOR2X1 _12977_ (
    .A(_2657_),
    .B(_2632_),
    .Y(_2660_)
);

AOI21X1 _12978_ (
    .A(_2660_),
    .B(\datapath.csr.mvect [16]),
    .C(\controlunit.mret_bF$buf2 ),
    .Y(_2661_)
);

OAI21X1 _12979_ (
    .A(\datapath.csr.mvect [16]),
    .B(_2660_),
    .C(_2661_),
    .Y(_2662_)
);

OAI21X1 _12980_ (
    .A(_2597__bF$buf4),
    .B(_2659_),
    .C(_2662_),
    .Y(\datapath.csr.csr_pcaddr [16])
);

INVX1 _12981_ (
    .A(\datapath.csr.mepc [15]),
    .Y(_2663_)
);

AOI21X1 _12982_ (
    .A(_2660_),
    .B(\datapath.csr.mvect [16]),
    .C(\datapath.csr.mvect [17]),
    .Y(_2664_)
);

INVX1 _12983_ (
    .A(_2660_),
    .Y(_2665_)
);

AND2X2 _12984_ (
    .A(\datapath.csr.mvect [16]),
    .B(\datapath.csr.mvect [17]),
    .Y(_2666_)
);

INVX1 _12985_ (
    .A(_2666_),
    .Y(_2667_)
);

OAI21X1 _12986_ (
    .A(_2667_),
    .B(_2665_),
    .C(_2597__bF$buf3),
    .Y(_2668_)
);

OAI22X1 _12987_ (
    .A(_2597__bF$buf2),
    .B(_2663_),
    .C(_2664_),
    .D(_2668_),
    .Y(\datapath.csr.csr_pcaddr [17])
);

INVX1 _12988_ (
    .A(\datapath.csr.mepc [16]),
    .Y(_2669_)
);

AOI21X1 _12989_ (
    .A(_2660_),
    .B(_2666_),
    .C(\datapath.csr.mvect [18]),
    .Y(_2670_)
);

NAND3X1 _12990_ (
    .A(\datapath.csr.mvect [16]),
    .B(\datapath.csr.mvect [17]),
    .C(\datapath.csr.mvect [18]),
    .Y(_2671_)
);

OAI21X1 _12991_ (
    .A(_2671_),
    .B(_2665_),
    .C(_2597__bF$buf1),
    .Y(_2672_)
);

OAI22X1 _12992_ (
    .A(_2597__bF$buf0),
    .B(_2669_),
    .C(_2670_),
    .D(_2672_),
    .Y(\datapath.csr.csr_pcaddr [18])
);

INVX1 _12993_ (
    .A(\datapath.csr.mepc [17]),
    .Y(_2673_)
);

INVX1 _12994_ (
    .A(_2671_),
    .Y(_2674_)
);

AOI21X1 _12995_ (
    .A(_2660_),
    .B(_2674_),
    .C(\datapath.csr.mvect [19]),
    .Y(_2675_)
);

INVX1 _12996_ (
    .A(\datapath.csr.mvect [19]),
    .Y(_2676_)
);

NOR2X1 _12997_ (
    .A(_2676_),
    .B(_2671_),
    .Y(_2677_)
);

NAND2X1 _12998_ (
    .A(_2677_),
    .B(_2660_),
    .Y(_2678_)
);

NAND2X1 _12999_ (
    .A(_2597__bF$buf5),
    .B(_2678_),
    .Y(_2679_)
);

OAI22X1 _13000_ (
    .A(_2597__bF$buf4),
    .B(_2673_),
    .C(_2675_),
    .D(_2679_),
    .Y(\datapath.csr.csr_pcaddr [19])
);

INVX1 _13001_ (
    .A(\datapath.csr.mepc [18]),
    .Y(_2680_)
);

AOI21X1 _13002_ (
    .A(_2660_),
    .B(_2677_),
    .C(\datapath.csr.mvect [20]),
    .Y(_2681_)
);

INVX1 _13003_ (
    .A(\datapath.csr.mvect [20]),
    .Y(_2682_)
);

OAI21X1 _13004_ (
    .A(_2682_),
    .B(_2678_),
    .C(_2597__bF$buf3),
    .Y(_2683_)
);

OAI22X1 _13005_ (
    .A(_2597__bF$buf2),
    .B(_2680_),
    .C(_2681_),
    .D(_2683_),
    .Y(\datapath.csr.csr_pcaddr [20])
);

INVX1 _13006_ (
    .A(\datapath.csr.mepc [19]),
    .Y(_2684_)
);

INVX1 _13007_ (
    .A(\datapath.csr.mvect [21]),
    .Y(_2685_)
);

NAND3X1 _13008_ (
    .A(\datapath.csr.mvect [20]),
    .B(_2677_),
    .C(_2660_),
    .Y(_2686_)
);

AND2X2 _13009_ (
    .A(_2686_),
    .B(_2685_),
    .Y(_2687_)
);

AND2X2 _13010_ (
    .A(\datapath.csr.mvect [18]),
    .B(\datapath.csr.mvect [19]),
    .Y(_2688_)
);

NAND2X1 _13011_ (
    .A(\datapath.csr.mvect [20]),
    .B(\datapath.csr.mvect [21]),
    .Y(_2689_)
);

INVX1 _13012_ (
    .A(_2689_),
    .Y(_2690_)
);

NAND3X1 _13013_ (
    .A(_2666_),
    .B(_2688_),
    .C(_2690_),
    .Y(_2691_)
);

OAI21X1 _13014_ (
    .A(_2691_),
    .B(_2665_),
    .C(_2597__bF$buf1),
    .Y(_2692_)
);

OAI22X1 _13015_ (
    .A(_2597__bF$buf0),
    .B(_2684_),
    .C(_2692_),
    .D(_2687_),
    .Y(\datapath.csr.csr_pcaddr [21])
);

INVX1 _13016_ (
    .A(\datapath.csr.mepc [20]),
    .Y(_2693_)
);

NOR3X1 _13017_ (
    .A(_2676_),
    .B(_2689_),
    .C(_2671_),
    .Y(_2694_)
);

NAND3X1 _13018_ (
    .A(_2631_),
    .B(_2656_),
    .C(_2694_),
    .Y(_2695_)
);

NOR2X1 _13019_ (
    .A(_2609_),
    .B(_2695_),
    .Y(_2696_)
);

AOI21X1 _13020_ (
    .A(_2696_),
    .B(\datapath.csr.mvect [22]),
    .C(\controlunit.mret_bF$buf1 ),
    .Y(_2697_)
);

OAI21X1 _13021_ (
    .A(\datapath.csr.mvect [22]),
    .B(_2696_),
    .C(_2697_),
    .Y(_2698_)
);

OAI21X1 _13022_ (
    .A(_2597__bF$buf5),
    .B(_2693_),
    .C(_2698_),
    .Y(\datapath.csr.csr_pcaddr [22])
);

INVX1 _13023_ (
    .A(\datapath.csr.mepc [21]),
    .Y(_2699_)
);

NAND2X1 _13024_ (
    .A(\datapath.csr.mvect [22]),
    .B(_2696_),
    .Y(_2700_)
);

OR2X2 _13025_ (
    .A(_2700_),
    .B(\datapath.csr.mvect [23]),
    .Y(_2701_)
);

AOI21X1 _13026_ (
    .A(_2700_),
    .B(\datapath.csr.mvect [23]),
    .C(\controlunit.mret_bF$buf0 ),
    .Y(_2702_)
);

AOI22X1 _13027_ (
    .A(\controlunit.mret_bF$buf4 ),
    .B(_2699_),
    .C(_2702_),
    .D(_2701_),
    .Y(\datapath.csr.csr_pcaddr [23])
);

INVX1 _13028_ (
    .A(\datapath.csr.mepc [22]),
    .Y(_2703_)
);

NAND2X1 _13029_ (
    .A(\datapath.csr.mvect [22]),
    .B(\datapath.csr.mvect [23]),
    .Y(_2704_)
);

NOR3X1 _13030_ (
    .A(_2609_),
    .B(_2704_),
    .C(_2695_),
    .Y(_2705_)
);

NOR2X1 _13031_ (
    .A(\datapath.csr.mvect [24]),
    .B(_2705_),
    .Y(_2706_)
);

INVX1 _13032_ (
    .A(\datapath.csr.mvect [24]),
    .Y(_2707_)
);

NAND2X1 _13033_ (
    .A(_2631_),
    .B(_2656_),
    .Y(_2708_)
);

NOR2X1 _13034_ (
    .A(_2691_),
    .B(_2708_),
    .Y(_2709_)
);

INVX1 _13035_ (
    .A(_2704_),
    .Y(_2710_)
);

NAND3X1 _13036_ (
    .A(_2613_),
    .B(_2710_),
    .C(_2709_),
    .Y(_2711_)
);

OAI21X1 _13037_ (
    .A(_2707_),
    .B(_2711_),
    .C(_2597__bF$buf4),
    .Y(_2712_)
);

OAI22X1 _13038_ (
    .A(_2597__bF$buf3),
    .B(_2703_),
    .C(_2706_),
    .D(_2712_),
    .Y(\datapath.csr.csr_pcaddr [24])
);

INVX1 _13039_ (
    .A(\datapath.csr.mepc [23]),
    .Y(_2713_)
);

AOI21X1 _13040_ (
    .A(_2705_),
    .B(\datapath.csr.mvect [24]),
    .C(\datapath.csr.mvect [25]),
    .Y(_2714_)
);

NAND2X1 _13041_ (
    .A(\datapath.csr.mvect [24]),
    .B(\datapath.csr.mvect [25]),
    .Y(_2715_)
);

OAI21X1 _13042_ (
    .A(_2715_),
    .B(_2711_),
    .C(_2597__bF$buf2),
    .Y(_2716_)
);

OAI22X1 _13043_ (
    .A(_2597__bF$buf1),
    .B(_2713_),
    .C(_2716_),
    .D(_2714_),
    .Y(\datapath.csr.csr_pcaddr [25])
);

INVX1 _13044_ (
    .A(\datapath.csr.mepc [24]),
    .Y(_2717_)
);

INVX1 _13045_ (
    .A(\datapath.csr.mvect [26]),
    .Y(_2718_)
);

OAI21X1 _13046_ (
    .A(_2715_),
    .B(_2711_),
    .C(_2718_),
    .Y(_2719_)
);

INVX1 _13047_ (
    .A(_2715_),
    .Y(_2720_)
);

NAND3X1 _13048_ (
    .A(\datapath.csr.mvect [26]),
    .B(_2720_),
    .C(_2705_),
    .Y(_2721_)
);

NAND3X1 _13049_ (
    .A(_2597__bF$buf0),
    .B(_2721_),
    .C(_2719_),
    .Y(_2722_)
);

OAI21X1 _13050_ (
    .A(_2597__bF$buf5),
    .B(_2717_),
    .C(_2722_),
    .Y(\datapath.csr.csr_pcaddr [26])
);

INVX1 _13051_ (
    .A(\datapath.csr.mvect [27]),
    .Y(_2723_)
);

NAND3X1 _13052_ (
    .A(_2597__bF$buf4),
    .B(_2723_),
    .C(_2721_),
    .Y(_2724_)
);

INVX1 _13053_ (
    .A(\datapath.csr.mepc [25]),
    .Y(_2725_)
);

NAND2X1 _13054_ (
    .A(\datapath.csr.mvect [26]),
    .B(\datapath.csr.mvect [27]),
    .Y(_2726_)
);

NOR2X1 _13055_ (
    .A(_2715_),
    .B(_2726_),
    .Y(_2727_)
);

AND2X2 _13056_ (
    .A(_2727_),
    .B(_2597__bF$buf3),
    .Y(_2728_)
);

AOI22X1 _13057_ (
    .A(\controlunit.mret_bF$buf3 ),
    .B(_2725_),
    .C(_2728_),
    .D(_2705_),
    .Y(_2729_)
);

AND2X2 _13058_ (
    .A(_2724_),
    .B(_2729_),
    .Y(\datapath.csr.csr_pcaddr [27])
);

INVX1 _13059_ (
    .A(\datapath.csr.mepc [26]),
    .Y(_2730_)
);

NOR3X1 _13060_ (
    .A(_2704_),
    .B(_2715_),
    .C(_2726_),
    .Y(_2731_)
);

INVX1 _13061_ (
    .A(_2731_),
    .Y(_2732_)
);

NOR3X1 _13062_ (
    .A(_2609_),
    .B(_2732_),
    .C(_2695_),
    .Y(_2733_)
);

NOR2X1 _13063_ (
    .A(\datapath.csr.mvect [28]),
    .B(_2733_),
    .Y(_2734_)
);

INVX1 _13064_ (
    .A(\datapath.csr.mvect [28]),
    .Y(_2735_)
);

NAND3X1 _13065_ (
    .A(_2613_),
    .B(_2731_),
    .C(_2709_),
    .Y(_2736_)
);

OAI21X1 _13066_ (
    .A(_2735_),
    .B(_2736_),
    .C(_2597__bF$buf2),
    .Y(_2737_)
);

OAI22X1 _13067_ (
    .A(_2597__bF$buf1),
    .B(_2730_),
    .C(_2734_),
    .D(_2737_),
    .Y(\datapath.csr.csr_pcaddr [28])
);

INVX1 _13068_ (
    .A(\datapath.csr.mepc [27]),
    .Y(_2738_)
);

NAND3X1 _13069_ (
    .A(\datapath.csr.mvect [28]),
    .B(_2731_),
    .C(_2696_),
    .Y(_2739_)
);

OR2X2 _13070_ (
    .A(_2739_),
    .B(\datapath.csr.mvect [29]),
    .Y(_2740_)
);

AOI21X1 _13071_ (
    .A(_2739_),
    .B(\datapath.csr.mvect [29]),
    .C(\controlunit.mret_bF$buf2 ),
    .Y(_2741_)
);

AOI22X1 _13072_ (
    .A(\controlunit.mret_bF$buf1 ),
    .B(_2738_),
    .C(_2741_),
    .D(_2740_),
    .Y(\datapath.csr.csr_pcaddr [29])
);

NAND2X1 _13073_ (
    .A(\datapath.csr.mvect [28]),
    .B(\datapath.csr.mvect [29]),
    .Y(_2742_)
);

NOR3X1 _13074_ (
    .A(_2576_),
    .B(_2742_),
    .C(_2575_),
    .Y(_2743_)
);

NAND3X1 _13075_ (
    .A(_2612_),
    .B(_2743_),
    .C(_2731_),
    .Y(_2744_)
);

NOR2X1 _13076_ (
    .A(_2695_),
    .B(_2744_),
    .Y(_2745_)
);

XNOR2X1 _13077_ (
    .A(_2745_),
    .B(\datapath.csr.mvect [30]),
    .Y(_2746_)
);

NAND2X1 _13078_ (
    .A(\controlunit.mret_bF$buf0 ),
    .B(\datapath.csr.mepc [28]),
    .Y(_2747_)
);

OAI21X1 _13079_ (
    .A(\controlunit.mret_bF$buf4 ),
    .B(_2746_),
    .C(_2747_),
    .Y(\datapath.csr.csr_pcaddr [30])
);

INVX1 _13080_ (
    .A(\datapath.csr.mepc [29]),
    .Y(_2748_)
);

INVX1 _13081_ (
    .A(_2742_),
    .Y(_2749_)
);

NAND2X1 _13082_ (
    .A(\datapath.csr.mvect [30]),
    .B(_2749_),
    .Y(_2750_)
);

INVX1 _13083_ (
    .A(_2750_),
    .Y(_2751_)
);

NAND3X1 _13084_ (
    .A(\datapath.csr.mvect [31]),
    .B(_2751_),
    .C(_2733_),
    .Y(_2752_)
);

INVX1 _13085_ (
    .A(\datapath.csr.mvect [31]),
    .Y(_2753_)
);

OAI21X1 _13086_ (
    .A(_2750_),
    .B(_2736_),
    .C(_2753_),
    .Y(_2754_)
);

NAND3X1 _13087_ (
    .A(_2597__bF$buf0),
    .B(_2752_),
    .C(_2754_),
    .Y(_2755_)
);

OAI21X1 _13088_ (
    .A(_2597__bF$buf5),
    .B(_2748_),
    .C(_2755_),
    .Y(\datapath.csr.csr_pcaddr [31])
);

NOR2X1 _13089_ (
    .A(\datapath.idinstr [31]),
    .B(\datapath.idinstr [30]),
    .Y(_2756_)
);

NAND3X1 _13090_ (
    .A(\datapath.idinstr [29]),
    .B(\datapath.idinstr [28]),
    .C(_2756_),
    .Y(_2757_)
);

INVX1 _13091_ (
    .A(\datapath.idinstr [27]),
    .Y(_2758_)
);

NOR2X1 _13092_ (
    .A(\datapath.idinstr [25]),
    .B(\datapath.idinstr_24_bF$buf4 ),
    .Y(_2759_)
);

NAND3X1 _13093_ (
    .A(_2758_),
    .B(\datapath.idinstr [26]),
    .C(_2759_),
    .Y(_2760_)
);

NOR2X1 _13094_ (
    .A(_2757_),
    .B(_2760_),
    .Y(_2761_)
);

NOR2X1 _13095_ (
    .A(\datapath.idinstr_23_bF$buf5 ),
    .B(\datapath.idinstr_22_bF$buf40 ),
    .Y(_2762_)
);

INVX1 _13096_ (
    .A(_2762_),
    .Y(_2763_)
);

INVX1 _13097_ (
    .A(\datapath.idinstr_20_bF$buf54 ),
    .Y(_2764_)
);

NAND2X1 _13098_ (
    .A(\datapath.idinstr_21_bF$buf50 ),
    .B(_2764_),
    .Y(_2765_)
);

NOR2X1 _13099_ (
    .A(_2765_),
    .B(_2763_),
    .Y(_2766_)
);

NAND2X1 _13100_ (
    .A(_2766_),
    .B(_2761_),
    .Y(_2767_)
);

INVX2 _13101_ (
    .A(_2767__bF$buf4),
    .Y(_2768_)
);

NAND2X1 _13102_ (
    .A(\datapath.csr.mcause [0]),
    .B(_2768_),
    .Y(_2769_)
);

NOR2X1 _13103_ (
    .A(\datapath.idinstr [27]),
    .B(\datapath.idinstr [26]),
    .Y(_2770_)
);

NAND2X1 _13104_ (
    .A(_2759_),
    .B(_2770_),
    .Y(_2771_)
);

NOR2X1 _13105_ (
    .A(_2771_),
    .B(_2757_),
    .Y(_2772_)
);

OR2X2 _13106_ (
    .A(_2764_),
    .B(\datapath.idinstr_21_bF$buf49 ),
    .Y(_2773_)
);

INVX1 _13107_ (
    .A(\datapath.idinstr_23_bF$buf4 ),
    .Y(_2774_)
);

NAND2X1 _13108_ (
    .A(\datapath.idinstr_22_bF$buf39 ),
    .B(_2774_),
    .Y(_2775_)
);

NOR2X1 _13109_ (
    .A(_2775_),
    .B(_2773_),
    .Y(_2776_)
);

NAND2X1 _13110_ (
    .A(_2776_),
    .B(_2772_),
    .Y(_2777_)
);

OAI21X1 _13111_ (
    .A(_2576_),
    .B(_2777_),
    .C(_2769_),
    .Y(\datapath.csr.csr_data [0])
);

INVX1 _13112_ (
    .A(\datapath.csr.mvect [1]),
    .Y(_2778_)
);

NAND2X1 _13113_ (
    .A(\datapath.csr.mcause [1]),
    .B(_2768_),
    .Y(_2779_)
);

OAI21X1 _13114_ (
    .A(_2778_),
    .B(_2777_),
    .C(_2779_),
    .Y(\datapath.csr.csr_data [1])
);

INVX1 _13115_ (
    .A(\datapath.csr.mcause [2]),
    .Y(_2780_)
);

INVX8 _13116_ (
    .A(_2777_),
    .Y(_2781_)
);

NOR2X1 _13117_ (
    .A(_2763_),
    .B(_2773_),
    .Y(_2782_)
);

AND2X2 _13118_ (
    .A(_2761_),
    .B(_2782_),
    .Y(_2783_)
);

AOI22X1 _13119_ (
    .A(\datapath.csr.mepc [0]),
    .B(_2783__bF$buf4),
    .C(\datapath.csr.mvect [2]),
    .D(_2781__bF$buf4),
    .Y(_2784_)
);

OAI21X1 _13120_ (
    .A(_2780_),
    .B(_2767__bF$buf3),
    .C(_2784_),
    .Y(\datapath.csr.csr_data [2])
);

NOR2X1 _13121_ (
    .A(\datapath.idinstr_21_bF$buf48 ),
    .B(\datapath.idinstr_20_bF$buf53 ),
    .Y(_2785_)
);

AND2X2 _13122_ (
    .A(_2772_),
    .B(_2762_),
    .Y(_2786_)
);

AND2X2 _13123_ (
    .A(_2786_),
    .B(_2785_),
    .Y(_2787_)
);

NAND2X1 _13124_ (
    .A(\datapath.csr.mstatus [0]),
    .B(_2787_),
    .Y(_2788_)
);

NAND2X1 _13125_ (
    .A(\datapath.csr.mcause [3]),
    .B(_2768_),
    .Y(_2789_)
);

AOI22X1 _13126_ (
    .A(\datapath.csr.mepc [1]),
    .B(_2783__bF$buf3),
    .C(\datapath.csr.mvect [3]),
    .D(_2781__bF$buf3),
    .Y(_2790_)
);

NAND3X1 _13127_ (
    .A(_2789_),
    .B(_2790_),
    .C(_2788_),
    .Y(\datapath.csr.csr_data [3])
);

INVX1 _13128_ (
    .A(\datapath.csr.mcause [4]),
    .Y(_2791_)
);

AOI22X1 _13129_ (
    .A(\datapath.csr.mepc [2]),
    .B(_2783__bF$buf2),
    .C(\datapath.csr.mvect [4]),
    .D(_2781__bF$buf2),
    .Y(_2792_)
);

OAI21X1 _13130_ (
    .A(_2791_),
    .B(_2767__bF$buf2),
    .C(_2792_),
    .Y(\datapath.csr.csr_data [4])
);

INVX1 _13131_ (
    .A(\datapath.csr.mcause [5]),
    .Y(_2793_)
);

AOI22X1 _13132_ (
    .A(\datapath.csr.mepc [3]),
    .B(_2783__bF$buf1),
    .C(\datapath.csr.mvect [5]),
    .D(_2781__bF$buf1),
    .Y(_2794_)
);

OAI21X1 _13133_ (
    .A(_2793_),
    .B(_2767__bF$buf1),
    .C(_2794_),
    .Y(\datapath.csr.csr_data [5])
);

INVX1 _13134_ (
    .A(\datapath.csr.mcause [6]),
    .Y(_2795_)
);

AOI22X1 _13135_ (
    .A(\datapath.csr.mepc [4]),
    .B(_2783__bF$buf0),
    .C(\datapath.csr.mvect [6]),
    .D(_2781__bF$buf0),
    .Y(_2796_)
);

OAI21X1 _13136_ (
    .A(_2795_),
    .B(_2767__bF$buf0),
    .C(_2796_),
    .Y(\datapath.csr.csr_data [6])
);

NAND2X1 _13137_ (
    .A(\datapath.csr.mstatus [1]),
    .B(_2787_),
    .Y(_2797_)
);

NAND2X1 _13138_ (
    .A(\datapath.csr.mcause [7]),
    .B(_2768_),
    .Y(_2798_)
);

AOI22X1 _13139_ (
    .A(\datapath.csr.mepc [5]),
    .B(_2783__bF$buf4),
    .C(\datapath.csr.mvect [7]),
    .D(_2781__bF$buf4),
    .Y(_2799_)
);

NAND3X1 _13140_ (
    .A(_2798_),
    .B(_2799_),
    .C(_2797_),
    .Y(\datapath.csr.csr_data [7])
);

AOI22X1 _13141_ (
    .A(\datapath.csr.mepc [6]),
    .B(_2783__bF$buf3),
    .C(\datapath.csr.mvect [8]),
    .D(_2781__bF$buf3),
    .Y(_2800_)
);

INVX1 _13142_ (
    .A(_2773_),
    .Y(_2801_)
);

AOI22X1 _13143_ (
    .A(_2786_),
    .B(_2801_),
    .C(\datapath.csr.mcause [8]),
    .D(_2768_),
    .Y(_2802_)
);

NAND2X1 _13144_ (
    .A(_2800_),
    .B(_2802_),
    .Y(\datapath.csr.csr_data [8])
);

INVX1 _13145_ (
    .A(\datapath.csr.mcause [9]),
    .Y(_2803_)
);

AOI22X1 _13146_ (
    .A(\datapath.csr.mepc [7]),
    .B(_2783__bF$buf2),
    .C(\datapath.csr.mvect [9]),
    .D(_2781__bF$buf2),
    .Y(_2804_)
);

OAI21X1 _13147_ (
    .A(_2803_),
    .B(_2767__bF$buf4),
    .C(_2804_),
    .Y(\datapath.csr.csr_data [9])
);

INVX1 _13148_ (
    .A(\datapath.csr.mcause [10]),
    .Y(_2805_)
);

AOI22X1 _13149_ (
    .A(\datapath.csr.mepc [8]),
    .B(_2783__bF$buf1),
    .C(\datapath.csr.mvect [10]),
    .D(_2781__bF$buf1),
    .Y(_2806_)
);

OAI21X1 _13150_ (
    .A(_2805_),
    .B(_2767__bF$buf3),
    .C(_2806_),
    .Y(\datapath.csr.csr_data [10])
);

AOI21X1 _13151_ (
    .A(\datapath.csr.mepc [9]),
    .B(_2783__bF$buf0),
    .C(_2787_),
    .Y(_2807_)
);

INVX1 _13152_ (
    .A(\datapath.csr.mip ),
    .Y(_2808_)
);

INVX1 _13153_ (
    .A(\datapath.csr.mie ),
    .Y(_2809_)
);

OAI22X1 _13154_ (
    .A(_2809_),
    .B(_2771_),
    .C(_2808_),
    .D(_2760_),
    .Y(_2810_)
);

NAND3X1 _13155_ (
    .A(_2774_),
    .B(\datapath.idinstr_22_bF$buf38 ),
    .C(_2785_),
    .Y(_2811_)
);

NOR2X1 _13156_ (
    .A(_2757_),
    .B(_2811_),
    .Y(_2812_)
);

NAND2X1 _13157_ (
    .A(_2812_),
    .B(_2810_),
    .Y(_2813_)
);

AOI22X1 _13158_ (
    .A(_2781__bF$buf0),
    .B(\datapath.csr.mvect [11]),
    .C(\datapath.csr.mcause [11]),
    .D(_2768_),
    .Y(_2814_)
);

NAND3X1 _13159_ (
    .A(_2813_),
    .B(_2814_),
    .C(_2807_),
    .Y(\datapath.csr.csr_data [11])
);

AOI21X1 _13160_ (
    .A(\datapath.csr.mvect [12]),
    .B(_2781__bF$buf4),
    .C(_2787_),
    .Y(_2815_)
);

AOI22X1 _13161_ (
    .A(\datapath.csr.mepc [10]),
    .B(_2783__bF$buf4),
    .C(\datapath.csr.mcause [12]),
    .D(_2768_),
    .Y(_2816_)
);

NAND2X1 _13162_ (
    .A(_2816_),
    .B(_2815_),
    .Y(\datapath.csr.csr_data [12])
);

INVX1 _13163_ (
    .A(\datapath.csr.mcause [13]),
    .Y(_2817_)
);

AOI22X1 _13164_ (
    .A(\datapath.csr.mepc [11]),
    .B(_2783__bF$buf3),
    .C(\datapath.csr.mvect [13]),
    .D(_2781__bF$buf3),
    .Y(_2818_)
);

OAI21X1 _13165_ (
    .A(_2817_),
    .B(_2767__bF$buf2),
    .C(_2818_),
    .Y(\datapath.csr.csr_data [13])
);

INVX1 _13166_ (
    .A(\datapath.csr.mcause [14]),
    .Y(_2819_)
);

AOI22X1 _13167_ (
    .A(\datapath.csr.mepc [12]),
    .B(_2783__bF$buf2),
    .C(\datapath.csr.mvect [14]),
    .D(_2781__bF$buf2),
    .Y(_2820_)
);

OAI21X1 _13168_ (
    .A(_2819_),
    .B(_2767__bF$buf1),
    .C(_2820_),
    .Y(\datapath.csr.csr_data [14])
);

INVX1 _13169_ (
    .A(\datapath.csr.mcause [15]),
    .Y(_2821_)
);

AOI22X1 _13170_ (
    .A(\datapath.csr.mepc [13]),
    .B(_2783__bF$buf1),
    .C(\datapath.csr.mvect [15]),
    .D(_2781__bF$buf1),
    .Y(_2822_)
);

OAI21X1 _13171_ (
    .A(_2821_),
    .B(_2767__bF$buf0),
    .C(_2822_),
    .Y(\datapath.csr.csr_data [15])
);

INVX1 _13172_ (
    .A(\datapath.csr.mcause [16]),
    .Y(_2823_)
);

AOI22X1 _13173_ (
    .A(\datapath.csr.mepc [14]),
    .B(_2783__bF$buf0),
    .C(\datapath.csr.mvect [16]),
    .D(_2781__bF$buf0),
    .Y(_2824_)
);

OAI21X1 _13174_ (
    .A(_2823_),
    .B(_2767__bF$buf4),
    .C(_2824_),
    .Y(\datapath.csr.csr_data [16])
);

INVX1 _13175_ (
    .A(\datapath.csr.mcause [17]),
    .Y(_2825_)
);

AOI22X1 _13176_ (
    .A(\datapath.csr.mepc [15]),
    .B(_2783__bF$buf4),
    .C(\datapath.csr.mvect [17]),
    .D(_2781__bF$buf4),
    .Y(_2826_)
);

OAI21X1 _13177_ (
    .A(_2825_),
    .B(_2767__bF$buf3),
    .C(_2826_),
    .Y(\datapath.csr.csr_data [17])
);

INVX1 _13178_ (
    .A(\datapath.csr.mcause [18]),
    .Y(_2827_)
);

AOI22X1 _13179_ (
    .A(\datapath.csr.mepc [16]),
    .B(_2783__bF$buf3),
    .C(\datapath.csr.mvect [18]),
    .D(_2781__bF$buf3),
    .Y(_2828_)
);

OAI21X1 _13180_ (
    .A(_2827_),
    .B(_2767__bF$buf2),
    .C(_2828_),
    .Y(\datapath.csr.csr_data [18])
);

INVX1 _13181_ (
    .A(\datapath.csr.mcause [19]),
    .Y(_2829_)
);

AOI22X1 _13182_ (
    .A(\datapath.csr.mepc [17]),
    .B(_2783__bF$buf2),
    .C(\datapath.csr.mvect [19]),
    .D(_2781__bF$buf2),
    .Y(_2830_)
);

OAI21X1 _13183_ (
    .A(_2829_),
    .B(_2767__bF$buf1),
    .C(_2830_),
    .Y(\datapath.csr.csr_data [19])
);

INVX1 _13184_ (
    .A(\datapath.csr.mcause [20]),
    .Y(_2831_)
);

AOI22X1 _13185_ (
    .A(\datapath.csr.mepc [18]),
    .B(_2783__bF$buf1),
    .C(\datapath.csr.mvect [20]),
    .D(_2781__bF$buf1),
    .Y(_2832_)
);

OAI21X1 _13186_ (
    .A(_2831_),
    .B(_2767__bF$buf0),
    .C(_2832_),
    .Y(\datapath.csr.csr_data [20])
);

INVX1 _13187_ (
    .A(\datapath.csr.mcause [21]),
    .Y(_2833_)
);

AOI22X1 _13188_ (
    .A(\datapath.csr.mepc [19]),
    .B(_2783__bF$buf0),
    .C(\datapath.csr.mvect [21]),
    .D(_2781__bF$buf0),
    .Y(_2834_)
);

OAI21X1 _13189_ (
    .A(_2833_),
    .B(_2767__bF$buf4),
    .C(_2834_),
    .Y(\datapath.csr.csr_data [21])
);

INVX1 _13190_ (
    .A(\datapath.csr.mcause [22]),
    .Y(_2835_)
);

AOI22X1 _13191_ (
    .A(\datapath.csr.mepc [20]),
    .B(_2783__bF$buf4),
    .C(\datapath.csr.mvect [22]),
    .D(_2781__bF$buf4),
    .Y(_2836_)
);

OAI21X1 _13192_ (
    .A(_2835_),
    .B(_2767__bF$buf3),
    .C(_2836_),
    .Y(\datapath.csr.csr_data [22])
);

INVX1 _13193_ (
    .A(\datapath.csr.mcause [23]),
    .Y(_2837_)
);

AOI22X1 _13194_ (
    .A(\datapath.csr.mepc [21]),
    .B(_2783__bF$buf3),
    .C(\datapath.csr.mvect [23]),
    .D(_2781__bF$buf3),
    .Y(_2838_)
);

OAI21X1 _13195_ (
    .A(_2837_),
    .B(_2767__bF$buf2),
    .C(_2838_),
    .Y(\datapath.csr.csr_data [23])
);

INVX1 _13196_ (
    .A(\datapath.csr.mcause [24]),
    .Y(_2839_)
);

AOI22X1 _13197_ (
    .A(\datapath.csr.mepc [22]),
    .B(_2783__bF$buf2),
    .C(\datapath.csr.mvect [24]),
    .D(_2781__bF$buf2),
    .Y(_2840_)
);

OAI21X1 _13198_ (
    .A(_2839_),
    .B(_2767__bF$buf1),
    .C(_2840_),
    .Y(\datapath.csr.csr_data [24])
);

INVX1 _13199_ (
    .A(\datapath.csr.mcause [25]),
    .Y(_2841_)
);

AOI22X1 _13200_ (
    .A(\datapath.csr.mepc [23]),
    .B(_2783__bF$buf1),
    .C(\datapath.csr.mvect [25]),
    .D(_2781__bF$buf1),
    .Y(_2842_)
);

OAI21X1 _13201_ (
    .A(_2841_),
    .B(_2767__bF$buf0),
    .C(_2842_),
    .Y(\datapath.csr.csr_data [25])
);

INVX1 _13202_ (
    .A(\datapath.csr.mcause [26]),
    .Y(_2843_)
);

AOI22X1 _13203_ (
    .A(\datapath.csr.mepc [24]),
    .B(_2783__bF$buf0),
    .C(\datapath.csr.mvect [26]),
    .D(_2781__bF$buf0),
    .Y(_2844_)
);

OAI21X1 _13204_ (
    .A(_2843_),
    .B(_2767__bF$buf4),
    .C(_2844_),
    .Y(\datapath.csr.csr_data [26])
);

INVX1 _13205_ (
    .A(\datapath.csr.mcause [27]),
    .Y(_2845_)
);

AOI22X1 _13206_ (
    .A(\datapath.csr.mepc [25]),
    .B(_2783__bF$buf4),
    .C(\datapath.csr.mvect [27]),
    .D(_2781__bF$buf4),
    .Y(_2846_)
);

OAI21X1 _13207_ (
    .A(_2845_),
    .B(_2767__bF$buf3),
    .C(_2846_),
    .Y(\datapath.csr.csr_data [27])
);

INVX1 _13208_ (
    .A(\datapath.csr.mcause [28]),
    .Y(_2847_)
);

AOI22X1 _13209_ (
    .A(\datapath.csr.mepc [26]),
    .B(_2783__bF$buf3),
    .C(\datapath.csr.mvect [28]),
    .D(_2781__bF$buf3),
    .Y(_2848_)
);

OAI21X1 _13210_ (
    .A(_2847_),
    .B(_2767__bF$buf2),
    .C(_2848_),
    .Y(\datapath.csr.csr_data [28])
);

INVX1 _13211_ (
    .A(\datapath.csr.mcause [29]),
    .Y(_2849_)
);

AOI22X1 _13212_ (
    .A(\datapath.csr.mepc [27]),
    .B(_2783__bF$buf2),
    .C(\datapath.csr.mvect [29]),
    .D(_2781__bF$buf2),
    .Y(_2850_)
);

OAI21X1 _13213_ (
    .A(_2849_),
    .B(_2767__bF$buf1),
    .C(_2850_),
    .Y(\datapath.csr.csr_data [29])
);

AOI22X1 _13214_ (
    .A(_2801_),
    .B(_2786_),
    .C(\datapath.csr.mvect [30]),
    .D(_2781__bF$buf1),
    .Y(_2851_)
);

AOI22X1 _13215_ (
    .A(\datapath.csr.mepc [28]),
    .B(_2783__bF$buf1),
    .C(\datapath.csr.mcause [30]),
    .D(_2768_),
    .Y(_2852_)
);

NAND2X1 _13216_ (
    .A(_2851_),
    .B(_2852_),
    .Y(\datapath.csr.csr_data [30])
);

INVX1 _13217_ (
    .A(\datapath.csr.mcause [31]),
    .Y(_2853_)
);

AOI22X1 _13218_ (
    .A(\datapath.csr.mepc [29]),
    .B(_2783__bF$buf0),
    .C(\datapath.csr.mvect [31]),
    .D(_2781__bF$buf0),
    .Y(_2854_)
);

OAI21X1 _13219_ (
    .A(_2853_),
    .B(_2767__bF$buf0),
    .C(_2854_),
    .Y(\datapath.csr.csr_data [31])
);

AND2X2 _13220_ (
    .A(_2597__bF$buf4),
    .B(\datapath.allowcsrwrite ),
    .Y(_2855_)
);

NAND2X1 _13221_ (
    .A(\datapath.meminstr [20]),
    .B(_2855_),
    .Y(_2856_)
);

NOR2X1 _13222_ (
    .A(\datapath.meminstr [21]),
    .B(_2856_),
    .Y(_2857_)
);

INVX1 _13223_ (
    .A(\datapath.meminstr [23]),
    .Y(_2858_)
);

NAND2X1 _13224_ (
    .A(\datapath.meminstr [22]),
    .B(_2858_),
    .Y(_2859_)
);

NOR2X1 _13225_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf5 ),
    .B(_2859_),
    .Y(_2860_)
);

INVX1 _13226_ (
    .A(\datapath.meminstr [28]),
    .Y(_2861_)
);

NOR2X1 _13227_ (
    .A(\datapath.meminstr [31]),
    .B(_2861_),
    .Y(_2862_)
);

INVX1 _13228_ (
    .A(\datapath.meminstr [30]),
    .Y(_2863_)
);

AND2X2 _13229_ (
    .A(_2863_),
    .B(\datapath.meminstr [29]),
    .Y(_2864_)
);

NAND2X1 _13230_ (
    .A(_2862_),
    .B(_2864_),
    .Y(_2865_)
);

NOR2X1 _13231_ (
    .A(\datapath.meminstr [25]),
    .B(\datapath.meminstr [24]),
    .Y(_2866_)
);

NOR2X1 _13232_ (
    .A(\datapath.meminstr [26]),
    .B(\datapath.meminstr [27]),
    .Y(_2867_)
);

NAND2X1 _13233_ (
    .A(_2866_),
    .B(_2867_),
    .Y(_2868_)
);

NOR2X1 _13234_ (
    .A(_2868_),
    .B(_2865_),
    .Y(_2869_)
);

NAND3X1 _13235_ (
    .A(_2860_),
    .B(_2857_),
    .C(_2869_),
    .Y(_2870_)
);

NOR2X1 _13236_ (
    .A(\datapath.csr.csr_wdata [0]),
    .B(_2870__bF$buf6),
    .Y(_2871_)
);

AOI21X1 _13237_ (
    .A(_2576_),
    .B(_2870__bF$buf5),
    .C(_2871_),
    .Y(\datapath.csr._13_ [0])
);

NOR2X1 _13238_ (
    .A(\datapath.csr.csr_wdata [1]),
    .B(_2870__bF$buf4),
    .Y(_2872_)
);

AOI21X1 _13239_ (
    .A(_2778_),
    .B(_2870__bF$buf3),
    .C(_2872_),
    .Y(\datapath.csr._13_ [1])
);

NOR2X1 _13240_ (
    .A(\datapath.csr.csr_wdata [2]),
    .B(_2870__bF$buf2),
    .Y(_2873_)
);

AOI21X1 _13241_ (
    .A(_2578_),
    .B(_2870__bF$buf1),
    .C(_2873_),
    .Y(\datapath.csr._13_ [2])
);

NOR2X1 _13242_ (
    .A(\datapath.csr.csr_wdata [3]),
    .B(_2870__bF$buf0),
    .Y(_2874_)
);

AOI21X1 _13243_ (
    .A(_2583_),
    .B(_2870__bF$buf6),
    .C(_2874_),
    .Y(\datapath.csr._13_ [3])
);

NOR2X1 _13244_ (
    .A(\datapath.csr.csr_wdata [4]),
    .B(_2870__bF$buf5),
    .Y(_2875_)
);

AOI21X1 _13245_ (
    .A(_2587_),
    .B(_2870__bF$buf4),
    .C(_2875_),
    .Y(\datapath.csr._13_ [4])
);

NOR2X1 _13246_ (
    .A(\datapath.csr.csr_wdata [5]),
    .B(_2870__bF$buf3),
    .Y(_2876_)
);

AOI21X1 _13247_ (
    .A(_2593_),
    .B(_2870__bF$buf2),
    .C(_2876_),
    .Y(\datapath.csr._13_ [5])
);

NOR2X1 _13248_ (
    .A(\datapath.csr.csr_wdata [6]),
    .B(_2870__bF$buf1),
    .Y(_2877_)
);

AOI21X1 _13249_ (
    .A(_2601_),
    .B(_2870__bF$buf0),
    .C(_2877_),
    .Y(\datapath.csr._13_ [6])
);

INVX1 _13250_ (
    .A(\datapath.csr.csr_wdata [7]),
    .Y(_2878_)
);

MUX2X1 _13251_ (
    .A(_2605_),
    .B(_2878_),
    .S(_2870__bF$buf6),
    .Y(\datapath.csr._13_ [7])
);

INVX1 _13252_ (
    .A(\datapath.csr.mvect [8]),
    .Y(_2879_)
);

NOR2X1 _13253_ (
    .A(\datapath.csr.csr_wdata [8]),
    .B(_2870__bF$buf5),
    .Y(_2880_)
);

AOI21X1 _13254_ (
    .A(_2879_),
    .B(_2870__bF$buf4),
    .C(_2880_),
    .Y(\datapath.csr._13_ [8])
);

INVX1 _13255_ (
    .A(\datapath.csr.mvect [9]),
    .Y(_2881_)
);

NOR2X1 _13256_ (
    .A(\datapath.csr.csr_wdata [9]),
    .B(_2870__bF$buf3),
    .Y(_2882_)
);

AOI21X1 _13257_ (
    .A(_2881_),
    .B(_2870__bF$buf2),
    .C(_2882_),
    .Y(\datapath.csr._13_ [9])
);

NOR2X1 _13258_ (
    .A(\datapath.csr.csr_wdata [10]),
    .B(_2870__bF$buf1),
    .Y(_2883_)
);

AOI21X1 _13259_ (
    .A(_2622_),
    .B(_2870__bF$buf0),
    .C(_2883_),
    .Y(\datapath.csr._13_ [10])
);

INVX1 _13260_ (
    .A(\datapath.csr.mvect [11]),
    .Y(_2884_)
);

INVX1 _13261_ (
    .A(\datapath.csr.csr_wdata [11]),
    .Y(_2885_)
);

MUX2X1 _13262_ (
    .A(_2884_),
    .B(_2885_),
    .S(_2870__bF$buf6),
    .Y(\datapath.csr._13_ [11])
);

NOR2X1 _13263_ (
    .A(\datapath.csr.csr_wdata [12]),
    .B(_2870__bF$buf5),
    .Y(_2886_)
);

AOI21X1 _13264_ (
    .A(_2635_),
    .B(_2870__bF$buf4),
    .C(_2886_),
    .Y(\datapath.csr._13_ [12])
);

NOR2X1 _13265_ (
    .A(\datapath.csr.csr_wdata [13]),
    .B(_2870__bF$buf3),
    .Y(_2887_)
);

AOI21X1 _13266_ (
    .A(_2639_),
    .B(_2870__bF$buf2),
    .C(_2887_),
    .Y(\datapath.csr._13_ [13])
);

NOR2X1 _13267_ (
    .A(\datapath.csr.csr_wdata [14]),
    .B(_2870__bF$buf1),
    .Y(_2888_)
);

AOI21X1 _13268_ (
    .A(_2645_),
    .B(_2870__bF$buf0),
    .C(_2888_),
    .Y(\datapath.csr._13_ [14])
);

NOR2X1 _13269_ (
    .A(\datapath.csr.csr_wdata [15]),
    .B(_2870__bF$buf6),
    .Y(_2889_)
);

AOI21X1 _13270_ (
    .A(_2652_),
    .B(_2870__bF$buf5),
    .C(_2889_),
    .Y(\datapath.csr._13_ [15])
);

INVX1 _13271_ (
    .A(\datapath.csr.mvect [16]),
    .Y(_2890_)
);

NOR2X1 _13272_ (
    .A(\datapath.csr.csr_wdata [16]),
    .B(_2870__bF$buf4),
    .Y(_2891_)
);

AOI21X1 _13273_ (
    .A(_2890_),
    .B(_2870__bF$buf3),
    .C(_2891_),
    .Y(\datapath.csr._13_ [16])
);

INVX1 _13274_ (
    .A(\datapath.csr.mvect [17]),
    .Y(_2892_)
);

NOR2X1 _13275_ (
    .A(\datapath.csr.csr_wdata [17]),
    .B(_2870__bF$buf2),
    .Y(_2893_)
);

AOI21X1 _13276_ (
    .A(_2892_),
    .B(_2870__bF$buf1),
    .C(_2893_),
    .Y(\datapath.csr._13_ [17])
);

INVX1 _13277_ (
    .A(\datapath.csr.mvect [18]),
    .Y(_2894_)
);

NOR2X1 _13278_ (
    .A(\datapath.csr.csr_wdata [18]),
    .B(_2870__bF$buf0),
    .Y(_2895_)
);

AOI21X1 _13279_ (
    .A(_2894_),
    .B(_2870__bF$buf6),
    .C(_2895_),
    .Y(\datapath.csr._13_ [18])
);

NOR2X1 _13280_ (
    .A(\datapath.csr.csr_wdata [19]),
    .B(_2870__bF$buf5),
    .Y(_2896_)
);

AOI21X1 _13281_ (
    .A(_2676_),
    .B(_2870__bF$buf4),
    .C(_2896_),
    .Y(\datapath.csr._13_ [19])
);

NOR2X1 _13282_ (
    .A(\datapath.csr.csr_wdata [20]),
    .B(_2870__bF$buf3),
    .Y(_2897_)
);

AOI21X1 _13283_ (
    .A(_2682_),
    .B(_2870__bF$buf2),
    .C(_2897_),
    .Y(\datapath.csr._13_ [20])
);

NOR2X1 _13284_ (
    .A(\datapath.csr.csr_wdata [21]),
    .B(_2870__bF$buf1),
    .Y(_2898_)
);

AOI21X1 _13285_ (
    .A(_2685_),
    .B(_2870__bF$buf0),
    .C(_2898_),
    .Y(\datapath.csr._13_ [21])
);

INVX1 _13286_ (
    .A(\datapath.csr.mvect [22]),
    .Y(_2899_)
);

NOR2X1 _13287_ (
    .A(\datapath.csr.csr_wdata [22]),
    .B(_2870__bF$buf6),
    .Y(_2900_)
);

AOI21X1 _13288_ (
    .A(_2899_),
    .B(_2870__bF$buf5),
    .C(_2900_),
    .Y(\datapath.csr._13_ [22])
);

INVX1 _13289_ (
    .A(\datapath.csr.mvect [23]),
    .Y(_2901_)
);

NOR2X1 _13290_ (
    .A(\datapath.csr.csr_wdata [23]),
    .B(_2870__bF$buf4),
    .Y(_2902_)
);

AOI21X1 _13291_ (
    .A(_2901_),
    .B(_2870__bF$buf3),
    .C(_2902_),
    .Y(\datapath.csr._13_ [23])
);

NOR2X1 _13292_ (
    .A(\datapath.csr.csr_wdata [24]),
    .B(_2870__bF$buf2),
    .Y(_2903_)
);

AOI21X1 _13293_ (
    .A(_2707_),
    .B(_2870__bF$buf1),
    .C(_2903_),
    .Y(\datapath.csr._13_ [24])
);

INVX1 _13294_ (
    .A(\datapath.csr.mvect [25]),
    .Y(_2904_)
);

NOR2X1 _13295_ (
    .A(\datapath.csr.csr_wdata [25]),
    .B(_2870__bF$buf0),
    .Y(_2905_)
);

AOI21X1 _13296_ (
    .A(_2904_),
    .B(_2870__bF$buf6),
    .C(_2905_),
    .Y(\datapath.csr._13_ [25])
);

NOR2X1 _13297_ (
    .A(\datapath.csr.csr_wdata [26]),
    .B(_2870__bF$buf5),
    .Y(_2906_)
);

AOI21X1 _13298_ (
    .A(_2718_),
    .B(_2870__bF$buf4),
    .C(_2906_),
    .Y(\datapath.csr._13_ [26])
);

NOR2X1 _13299_ (
    .A(\datapath.csr.csr_wdata [27]),
    .B(_2870__bF$buf3),
    .Y(_2907_)
);

AOI21X1 _13300_ (
    .A(_2723_),
    .B(_2870__bF$buf2),
    .C(_2907_),
    .Y(\datapath.csr._13_ [27])
);

NOR2X1 _13301_ (
    .A(\datapath.csr.csr_wdata [28]),
    .B(_2870__bF$buf1),
    .Y(_2908_)
);

AOI21X1 _13302_ (
    .A(_2735_),
    .B(_2870__bF$buf0),
    .C(_2908_),
    .Y(\datapath.csr._13_ [28])
);

INVX1 _13303_ (
    .A(\datapath.csr.mvect [29]),
    .Y(_2909_)
);

NOR2X1 _13304_ (
    .A(\datapath.csr.csr_wdata [29]),
    .B(_2870__bF$buf6),
    .Y(_2910_)
);

AOI21X1 _13305_ (
    .A(_2909_),
    .B(_2870__bF$buf5),
    .C(_2910_),
    .Y(\datapath.csr._13_ [29])
);

INVX1 _13306_ (
    .A(\datapath.csr.mvect [30]),
    .Y(_2911_)
);

NOR2X1 _13307_ (
    .A(\datapath.csr.csr_wdata [30]),
    .B(_2870__bF$buf4),
    .Y(_2912_)
);

AOI21X1 _13308_ (
    .A(_2911_),
    .B(_2870__bF$buf3),
    .C(_2912_),
    .Y(\datapath.csr._13_ [30])
);

NOR2X1 _13309_ (
    .A(\datapath.csr.csr_wdata [31]),
    .B(_2870__bF$buf2),
    .Y(_2913_)
);

AOI21X1 _13310_ (
    .A(_2753_),
    .B(_2870__bF$buf1),
    .C(_2913_),
    .Y(\datapath.csr._13_ [31])
);

NAND2X1 _13311_ (
    .A(_2860_),
    .B(_2869_),
    .Y(_2914_)
);

NOR2X1 _13312_ (
    .A(\datapath.meminstr [21]),
    .B(\datapath.meminstr [20]),
    .Y(_2915_)
);

NAND2X1 _13313_ (
    .A(_2915_),
    .B(_2855_),
    .Y(_2916_)
);

NOR2X1 _13314_ (
    .A(_2916_),
    .B(_2914_),
    .Y(_2917_)
);

MUX2X1 _13315_ (
    .A(_2885_),
    .B(_2809_),
    .S(_2917_),
    .Y(\datapath.csr._20_ )
);

INVX1 _13316_ (
    .A(\datapath.meminstr [27]),
    .Y(_2918_)
);

AND2X2 _13317_ (
    .A(_2918_),
    .B(\datapath.meminstr [29]),
    .Y(_2919_)
);

NAND3X1 _13318_ (
    .A(_2863_),
    .B(_2862_),
    .C(_2919_),
    .Y(_2920_)
);

NOR2X1 _13319_ (
    .A(\datapath.meminstr [23]),
    .B(\datapath.meminstr [22]),
    .Y(_2921_)
);

NAND3X1 _13320_ (
    .A(\datapath.meminstr [26]),
    .B(_2866_),
    .C(_2921_),
    .Y(_2922_)
);

NOR2X1 _13321_ (
    .A(_2922_),
    .B(_2920_),
    .Y(_2923_)
);

NAND2X1 _13322_ (
    .A(_2857_),
    .B(_2923_),
    .Y(_2924_)
);

MUX2X1 _13323_ (
    .A(\datapath.csr.mepc [0]),
    .B(\datapath.csr.csr_wdata [2]),
    .S(_2924__bF$buf6),
    .Y(_2925_)
);

NAND2X1 _13324_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf4 ),
    .B(\datapath.csr.csr_mepc [2]),
    .Y(_2926_)
);

OAI21X1 _13325_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf3 ),
    .B(_2925_),
    .C(_2926_),
    .Y(\datapath.csr._26_ [0])
);

MUX2X1 _13326_ (
    .A(\datapath.csr.mepc [1]),
    .B(\datapath.csr.csr_wdata [3]),
    .S(_2924__bF$buf5),
    .Y(_2927_)
);

NAND2X1 _13327_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf2 ),
    .B(\datapath.csr.csr_mepc [3]),
    .Y(_2928_)
);

OAI21X1 _13328_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf1 ),
    .B(_2927_),
    .C(_2928_),
    .Y(\datapath.csr._26_ [1])
);

MUX2X1 _13329_ (
    .A(\datapath.csr.mepc [2]),
    .B(\datapath.csr.csr_wdata [4]),
    .S(_2924__bF$buf4),
    .Y(_2929_)
);

NAND2X1 _13330_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf0 ),
    .B(\datapath.csr.csr_mepc [4]),
    .Y(_2930_)
);

OAI21X1 _13331_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf7 ),
    .B(_2929_),
    .C(_2930_),
    .Y(\datapath.csr._26_ [2])
);

MUX2X1 _13332_ (
    .A(\datapath.csr.mepc [3]),
    .B(\datapath.csr.csr_wdata [5]),
    .S(_2924__bF$buf3),
    .Y(_2931_)
);

NAND2X1 _13333_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf6 ),
    .B(\datapath.csr.csr_mepc [5]),
    .Y(_2932_)
);

OAI21X1 _13334_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf5 ),
    .B(_2931_),
    .C(_2932_),
    .Y(\datapath.csr._26_ [3])
);

NAND2X1 _13335_ (
    .A(_2598_),
    .B(_2924__bF$buf2),
    .Y(_2933_)
);

OAI21X1 _13336_ (
    .A(\datapath.csr.csr_wdata [6]),
    .B(_2924__bF$buf1),
    .C(_2933_),
    .Y(_2934_)
);

NAND2X1 _13337_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf4 ),
    .B(\datapath.csr.csr_mepc [6]),
    .Y(_2935_)
);

OAI21X1 _13338_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf3 ),
    .B(_2934_),
    .C(_2935_),
    .Y(\datapath.csr._26_ [4])
);

NAND2X1 _13339_ (
    .A(_2604_),
    .B(_2924__bF$buf0),
    .Y(_2936_)
);

OAI21X1 _13340_ (
    .A(\datapath.csr.csr_wdata [7]),
    .B(_2924__bF$buf6),
    .C(_2936_),
    .Y(_2937_)
);

NAND2X1 _13341_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf2 ),
    .B(\datapath.csr.csr_mepc [7]),
    .Y(_2938_)
);

OAI21X1 _13342_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf1 ),
    .B(_2937_),
    .C(_2938_),
    .Y(\datapath.csr._26_ [5])
);

NAND2X1 _13343_ (
    .A(_2611_),
    .B(_2924__bF$buf5),
    .Y(_2939_)
);

OAI21X1 _13344_ (
    .A(\datapath.csr.csr_wdata [8]),
    .B(_2924__bF$buf4),
    .C(_2939_),
    .Y(_2940_)
);

NAND2X1 _13345_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf0 ),
    .B(\datapath.csr.csr_mepc [8]),
    .Y(_2941_)
);

OAI21X1 _13346_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf7 ),
    .B(_2940_),
    .C(_2941_),
    .Y(\datapath.csr._26_ [6])
);

NAND2X1 _13347_ (
    .A(_2617_),
    .B(_2924__bF$buf3),
    .Y(_2942_)
);

OAI21X1 _13348_ (
    .A(\datapath.csr.csr_wdata [9]),
    .B(_2924__bF$buf2),
    .C(_2942_),
    .Y(_2943_)
);

NAND2X1 _13349_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf6 ),
    .B(\datapath.csr.csr_mepc [9]),
    .Y(_2944_)
);

OAI21X1 _13350_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf5 ),
    .B(_2943_),
    .C(_2944_),
    .Y(\datapath.csr._26_ [7])
);

NAND2X1 _13351_ (
    .A(_2623_),
    .B(_2924__bF$buf1),
    .Y(_2945_)
);

OAI21X1 _13352_ (
    .A(\datapath.csr.csr_wdata [10]),
    .B(_2924__bF$buf0),
    .C(_2945_),
    .Y(_2946_)
);

NAND2X1 _13353_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf4 ),
    .B(\datapath.csr.csr_mepc [10]),
    .Y(_2947_)
);

OAI21X1 _13354_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf3 ),
    .B(_2946_),
    .C(_2947_),
    .Y(\datapath.csr._26_ [8])
);

MUX2X1 _13355_ (
    .A(\datapath.csr.mepc [9]),
    .B(\datapath.csr.csr_wdata [11]),
    .S(_2924__bF$buf6),
    .Y(_2948_)
);

NAND2X1 _13356_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf2 ),
    .B(\datapath.csr.csr_mepc [11]),
    .Y(_2949_)
);

OAI21X1 _13357_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf1 ),
    .B(_2948_),
    .C(_2949_),
    .Y(\datapath.csr._26_ [9])
);

MUX2X1 _13358_ (
    .A(\datapath.csr.mepc [10]),
    .B(\datapath.csr.csr_wdata [12]),
    .S(_2924__bF$buf5),
    .Y(_2950_)
);

NAND2X1 _13359_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf0 ),
    .B(\datapath.csr.csr_mepc [12]),
    .Y(_2951_)
);

OAI21X1 _13360_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf7 ),
    .B(_2950_),
    .C(_2951_),
    .Y(\datapath.csr._26_ [10])
);

NAND2X1 _13361_ (
    .A(_2638_),
    .B(_2924__bF$buf4),
    .Y(_2952_)
);

OAI21X1 _13362_ (
    .A(\datapath.csr.csr_wdata [13]),
    .B(_2924__bF$buf3),
    .C(_2952_),
    .Y(_2953_)
);

NAND2X1 _13363_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf6 ),
    .B(\datapath.csr.csr_mepc [13]),
    .Y(_2954_)
);

OAI21X1 _13364_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf5 ),
    .B(_2953_),
    .C(_2954_),
    .Y(\datapath.csr._26_ [11])
);

NAND2X1 _13365_ (
    .A(_2644_),
    .B(_2924__bF$buf2),
    .Y(_2955_)
);

OAI21X1 _13366_ (
    .A(\datapath.csr.csr_wdata [14]),
    .B(_2924__bF$buf1),
    .C(_2955_),
    .Y(_2956_)
);

NAND2X1 _13367_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf4 ),
    .B(\datapath.csr.csr_mepc [14]),
    .Y(_2957_)
);

OAI21X1 _13368_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf3 ),
    .B(_2956_),
    .C(_2957_),
    .Y(\datapath.csr._26_ [12])
);

NAND2X1 _13369_ (
    .A(_2651_),
    .B(_2924__bF$buf0),
    .Y(_2958_)
);

OAI21X1 _13370_ (
    .A(\datapath.csr.csr_wdata [15]),
    .B(_2924__bF$buf6),
    .C(_2958_),
    .Y(_2959_)
);

NAND2X1 _13371_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf2 ),
    .B(\datapath.csr.csr_mepc [15]),
    .Y(_2960_)
);

OAI21X1 _13372_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf1 ),
    .B(_2959_),
    .C(_2960_),
    .Y(\datapath.csr._26_ [13])
);

NAND2X1 _13373_ (
    .A(_2659_),
    .B(_2924__bF$buf5),
    .Y(_2961_)
);

OAI21X1 _13374_ (
    .A(\datapath.csr.csr_wdata [16]),
    .B(_2924__bF$buf4),
    .C(_2961_),
    .Y(_2962_)
);

NAND2X1 _13375_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf0 ),
    .B(\datapath.csr.csr_mepc [16]),
    .Y(_2963_)
);

OAI21X1 _13376_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf7 ),
    .B(_2962_),
    .C(_2963_),
    .Y(\datapath.csr._26_ [14])
);

NAND2X1 _13377_ (
    .A(_2663_),
    .B(_2924__bF$buf3),
    .Y(_2964_)
);

OAI21X1 _13378_ (
    .A(\datapath.csr.csr_wdata [17]),
    .B(_2924__bF$buf2),
    .C(_2964_),
    .Y(_2965_)
);

NAND2X1 _13379_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf6 ),
    .B(\datapath.csr.csr_mepc [17]),
    .Y(_2966_)
);

OAI21X1 _13380_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf5 ),
    .B(_2965_),
    .C(_2966_),
    .Y(\datapath.csr._26_ [15])
);

NAND2X1 _13381_ (
    .A(_2669_),
    .B(_2924__bF$buf1),
    .Y(_2967_)
);

OAI21X1 _13382_ (
    .A(\datapath.csr.csr_wdata [18]),
    .B(_2924__bF$buf0),
    .C(_2967_),
    .Y(_2968_)
);

NAND2X1 _13383_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf4 ),
    .B(\datapath.csr.csr_mepc [18]),
    .Y(_2969_)
);

OAI21X1 _13384_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf3 ),
    .B(_2968_),
    .C(_2969_),
    .Y(\datapath.csr._26_ [16])
);

NAND2X1 _13385_ (
    .A(_2673_),
    .B(_2924__bF$buf6),
    .Y(_2970_)
);

OAI21X1 _13386_ (
    .A(\datapath.csr.csr_wdata [19]),
    .B(_2924__bF$buf5),
    .C(_2970_),
    .Y(_2971_)
);

NAND2X1 _13387_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf2 ),
    .B(\datapath.csr.csr_mepc [19]),
    .Y(_2972_)
);

OAI21X1 _13388_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf1 ),
    .B(_2971_),
    .C(_2972_),
    .Y(\datapath.csr._26_ [17])
);

NAND2X1 _13389_ (
    .A(_2680_),
    .B(_2924__bF$buf4),
    .Y(_2973_)
);

OAI21X1 _13390_ (
    .A(\datapath.csr.csr_wdata [20]),
    .B(_2924__bF$buf3),
    .C(_2973_),
    .Y(_2974_)
);

NAND2X1 _13391_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf0 ),
    .B(\datapath.csr.csr_mepc [20]),
    .Y(_2975_)
);

OAI21X1 _13392_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf7 ),
    .B(_2974_),
    .C(_2975_),
    .Y(\datapath.csr._26_ [18])
);

NAND2X1 _13393_ (
    .A(_2684_),
    .B(_2924__bF$buf2),
    .Y(_2976_)
);

OAI21X1 _13394_ (
    .A(\datapath.csr.csr_wdata [21]),
    .B(_2924__bF$buf1),
    .C(_2976_),
    .Y(_2977_)
);

NAND2X1 _13395_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf6 ),
    .B(\datapath.csr.csr_mepc [21]),
    .Y(_2978_)
);

OAI21X1 _13396_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf5 ),
    .B(_2977_),
    .C(_2978_),
    .Y(\datapath.csr._26_ [19])
);

NAND2X1 _13397_ (
    .A(_2693_),
    .B(_2924__bF$buf0),
    .Y(_2979_)
);

OAI21X1 _13398_ (
    .A(\datapath.csr.csr_wdata [22]),
    .B(_2924__bF$buf6),
    .C(_2979_),
    .Y(_2980_)
);

NAND2X1 _13399_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf4 ),
    .B(\datapath.csr.csr_mepc [22]),
    .Y(_2981_)
);

OAI21X1 _13400_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf3 ),
    .B(_2980_),
    .C(_2981_),
    .Y(\datapath.csr._26_ [20])
);

NAND2X1 _13401_ (
    .A(_2699_),
    .B(_2924__bF$buf5),
    .Y(_2982_)
);

OAI21X1 _13402_ (
    .A(\datapath.csr.csr_wdata [23]),
    .B(_2924__bF$buf4),
    .C(_2982_),
    .Y(_2983_)
);

NAND2X1 _13403_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf2 ),
    .B(\datapath.csr.csr_mepc [23]),
    .Y(_2984_)
);

OAI21X1 _13404_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf1 ),
    .B(_2983_),
    .C(_2984_),
    .Y(\datapath.csr._26_ [21])
);

NAND2X1 _13405_ (
    .A(_2703_),
    .B(_2924__bF$buf3),
    .Y(_2985_)
);

OAI21X1 _13406_ (
    .A(\datapath.csr.csr_wdata [24]),
    .B(_2924__bF$buf2),
    .C(_2985_),
    .Y(_2986_)
);

NAND2X1 _13407_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf0 ),
    .B(\datapath.csr.csr_mepc [24]),
    .Y(_2987_)
);

OAI21X1 _13408_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf7 ),
    .B(_2986_),
    .C(_2987_),
    .Y(\datapath.csr._26_ [22])
);

NAND2X1 _13409_ (
    .A(_2713_),
    .B(_2924__bF$buf1),
    .Y(_2988_)
);

OAI21X1 _13410_ (
    .A(\datapath.csr.csr_wdata [25]),
    .B(_2924__bF$buf0),
    .C(_2988_),
    .Y(_2989_)
);

NAND2X1 _13411_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf6 ),
    .B(\datapath.csr.csr_mepc [25]),
    .Y(_2990_)
);

OAI21X1 _13412_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf5 ),
    .B(_2989_),
    .C(_2990_),
    .Y(\datapath.csr._26_ [23])
);

NAND2X1 _13413_ (
    .A(_2717_),
    .B(_2924__bF$buf6),
    .Y(_2991_)
);

OAI21X1 _13414_ (
    .A(\datapath.csr.csr_wdata [26]),
    .B(_2924__bF$buf5),
    .C(_2991_),
    .Y(_2992_)
);

NAND2X1 _13415_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf4 ),
    .B(\datapath.csr.csr_mepc [26]),
    .Y(_2993_)
);

OAI21X1 _13416_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf3 ),
    .B(_2992_),
    .C(_2993_),
    .Y(\datapath.csr._26_ [24])
);

NAND2X1 _13417_ (
    .A(_2725_),
    .B(_2924__bF$buf4),
    .Y(_2994_)
);

OAI21X1 _13418_ (
    .A(\datapath.csr.csr_wdata [27]),
    .B(_2924__bF$buf3),
    .C(_2994_),
    .Y(_2995_)
);

NAND2X1 _13419_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf2 ),
    .B(\datapath.csr.csr_mepc [27]),
    .Y(_2996_)
);

OAI21X1 _13420_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf1 ),
    .B(_2995_),
    .C(_2996_),
    .Y(\datapath.csr._26_ [25])
);

NAND2X1 _13421_ (
    .A(_2730_),
    .B(_2924__bF$buf2),
    .Y(_2997_)
);

OAI21X1 _13422_ (
    .A(\datapath.csr.csr_wdata [28]),
    .B(_2924__bF$buf1),
    .C(_2997_),
    .Y(_2998_)
);

NAND2X1 _13423_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf0 ),
    .B(\datapath.csr.csr_mepc [28]),
    .Y(_2999_)
);

OAI21X1 _13424_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf7 ),
    .B(_2998_),
    .C(_2999_),
    .Y(\datapath.csr._26_ [26])
);

NAND2X1 _13425_ (
    .A(_2738_),
    .B(_2924__bF$buf0),
    .Y(_3000_)
);

OAI21X1 _13426_ (
    .A(\datapath.csr.csr_wdata [29]),
    .B(_2924__bF$buf6),
    .C(_3000_),
    .Y(_3001_)
);

NAND2X1 _13427_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf6 ),
    .B(\datapath.csr.csr_mepc [29]),
    .Y(_3002_)
);

OAI21X1 _13428_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf5 ),
    .B(_3001_),
    .C(_3002_),
    .Y(\datapath.csr._26_ [27])
);

MUX2X1 _13429_ (
    .A(\datapath.csr.mepc [28]),
    .B(\datapath.csr.csr_wdata [30]),
    .S(_2924__bF$buf5),
    .Y(_3003_)
);

NAND2X1 _13430_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf4 ),
    .B(\datapath.csr.csr_mepc [30]),
    .Y(_3004_)
);

OAI21X1 _13431_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf3 ),
    .B(_3003_),
    .C(_3004_),
    .Y(\datapath.csr._26_ [28])
);

NAND2X1 _13432_ (
    .A(_2748_),
    .B(_2924__bF$buf4),
    .Y(_3005_)
);

OAI21X1 _13433_ (
    .A(\datapath.csr.csr_wdata [31]),
    .B(_2924__bF$buf3),
    .C(_3005_),
    .Y(_3006_)
);

NAND2X1 _13434_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf2 ),
    .B(\datapath.csr.csr_mepc [31]),
    .Y(_3007_)
);

OAI21X1 _13435_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf1 ),
    .B(_3006_),
    .C(_3007_),
    .Y(\datapath.csr._26_ [29])
);

NAND2X1 _13436_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf0 ),
    .B(\datapath.csr.csr_mcause [0]),
    .Y(_3008_)
);

INVX1 _13437_ (
    .A(_2921_),
    .Y(_3009_)
);

NAND3X1 _13438_ (
    .A(\datapath.meminstr [26]),
    .B(_2918_),
    .C(_2866_),
    .Y(_3010_)
);

NOR3X1 _13439_ (
    .A(_3009_),
    .B(_3010_),
    .C(_2865_),
    .Y(_3011_)
);

NAND2X1 _13440_ (
    .A(\datapath.meminstr [21]),
    .B(_2855_),
    .Y(_3012_)
);

NOR2X1 _13441_ (
    .A(\datapath.meminstr [20]),
    .B(_3012_),
    .Y(_3013_)
);

NAND2X1 _13442_ (
    .A(_3013_),
    .B(_3011_),
    .Y(_3014_)
);

INVX1 _13443_ (
    .A(_3014__bF$buf6),
    .Y(_3015_)
);

NOR2X1 _13444_ (
    .A(\datapath.csr.mcause [0]),
    .B(_3015_),
    .Y(_3016_)
);

INVX8 _13445_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf7 ),
    .Y(_3017_)
);

NAND2X1 _13446_ (
    .A(_3013_),
    .B(_2923_),
    .Y(_3018_)
);

OAI21X1 _13447_ (
    .A(\datapath.csr.csr_wdata [0]),
    .B(_3018_),
    .C(_3017__bF$buf4),
    .Y(_3019_)
);

OAI21X1 _13448_ (
    .A(_3019_),
    .B(_3016_),
    .C(_3008_),
    .Y(\datapath.csr._32_ [0])
);

NAND2X1 _13449_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf6 ),
    .B(\datapath.csr.csr_mcause [1]),
    .Y(_3020_)
);

NOR2X1 _13450_ (
    .A(\datapath.csr.mcause [1]),
    .B(_3015_),
    .Y(_3021_)
);

OAI21X1 _13451_ (
    .A(\datapath.csr.csr_wdata [1]),
    .B(_3018_),
    .C(_3017__bF$buf3),
    .Y(_3022_)
);

OAI21X1 _13452_ (
    .A(_3022_),
    .B(_3021_),
    .C(_3020_),
    .Y(\datapath.csr._32_ [1])
);

NAND2X1 _13453_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf5 ),
    .B(\datapath.csr.csr_mcause [2]),
    .Y(_3023_)
);

NAND2X1 _13454_ (
    .A(_2780_),
    .B(_3018_),
    .Y(_3024_)
);

OAI21X1 _13455_ (
    .A(\datapath.csr.csr_wdata [2]),
    .B(_3014__bF$buf5),
    .C(_3024_),
    .Y(_3025_)
);

OAI21X1 _13456_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf4 ),
    .B(_3025_),
    .C(_3023_),
    .Y(\datapath.csr._32_ [2])
);

NAND2X1 _13457_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf3 ),
    .B(\datapath.csr.csr_mcause [3]),
    .Y(_3026_)
);

NOR2X1 _13458_ (
    .A(\datapath.csr.mcause [3]),
    .B(_3015_),
    .Y(_3027_)
);

OAI21X1 _13459_ (
    .A(\datapath.csr.csr_wdata [3]),
    .B(_3018_),
    .C(_3017__bF$buf2),
    .Y(_3028_)
);

OAI21X1 _13460_ (
    .A(_3028_),
    .B(_3027_),
    .C(_3026_),
    .Y(\datapath.csr._32_ [3])
);

OAI21X1 _13461_ (
    .A(\datapath.csr.csr_wdata [4]),
    .B(_3014__bF$buf4),
    .C(_3017__bF$buf1),
    .Y(_3029_)
);

AOI21X1 _13462_ (
    .A(_2791_),
    .B(_3014__bF$buf3),
    .C(_3029_),
    .Y(\datapath.csr._32_ [4])
);

OAI21X1 _13463_ (
    .A(\datapath.csr.csr_wdata [5]),
    .B(_3014__bF$buf2),
    .C(_3017__bF$buf0),
    .Y(_3030_)
);

AOI21X1 _13464_ (
    .A(_2793_),
    .B(_3014__bF$buf1),
    .C(_3030_),
    .Y(\datapath.csr._32_ [5])
);

OAI21X1 _13465_ (
    .A(\datapath.csr.csr_wdata [6]),
    .B(_3014__bF$buf0),
    .C(_3017__bF$buf4),
    .Y(_3031_)
);

AOI21X1 _13466_ (
    .A(_2795_),
    .B(_3014__bF$buf6),
    .C(_3031_),
    .Y(\datapath.csr._32_ [6])
);

INVX1 _13467_ (
    .A(\datapath.csr.mcause [7]),
    .Y(_3032_)
);

OAI21X1 _13468_ (
    .A(\datapath.csr.csr_wdata [7]),
    .B(_3014__bF$buf5),
    .C(_3017__bF$buf3),
    .Y(_3033_)
);

AOI21X1 _13469_ (
    .A(_3032_),
    .B(_3014__bF$buf4),
    .C(_3033_),
    .Y(\datapath.csr._32_ [7])
);

INVX1 _13470_ (
    .A(\datapath.csr.mcause [8]),
    .Y(_3034_)
);

OAI21X1 _13471_ (
    .A(\datapath.csr.csr_wdata [8]),
    .B(_3014__bF$buf3),
    .C(_3017__bF$buf2),
    .Y(_3035_)
);

AOI21X1 _13472_ (
    .A(_3034_),
    .B(_3014__bF$buf2),
    .C(_3035_),
    .Y(\datapath.csr._32_ [8])
);

OAI21X1 _13473_ (
    .A(\datapath.csr.csr_wdata [9]),
    .B(_3014__bF$buf1),
    .C(_3017__bF$buf1),
    .Y(_3036_)
);

AOI21X1 _13474_ (
    .A(_2803_),
    .B(_3014__bF$buf0),
    .C(_3036_),
    .Y(\datapath.csr._32_ [9])
);

OAI21X1 _13475_ (
    .A(\datapath.csr.csr_wdata [10]),
    .B(_3014__bF$buf6),
    .C(_3017__bF$buf0),
    .Y(_3037_)
);

AOI21X1 _13476_ (
    .A(_2805_),
    .B(_3014__bF$buf5),
    .C(_3037_),
    .Y(\datapath.csr._32_ [10])
);

INVX1 _13477_ (
    .A(\datapath.csr.mcause [11]),
    .Y(_3038_)
);

OAI21X1 _13478_ (
    .A(\datapath.csr.csr_wdata [11]),
    .B(_3014__bF$buf4),
    .C(_3017__bF$buf4),
    .Y(_3039_)
);

AOI21X1 _13479_ (
    .A(_3038_),
    .B(_3014__bF$buf3),
    .C(_3039_),
    .Y(\datapath.csr._32_ [11])
);

INVX1 _13480_ (
    .A(\datapath.csr.mcause [12]),
    .Y(_3040_)
);

OAI21X1 _13481_ (
    .A(\datapath.csr.csr_wdata [12]),
    .B(_3014__bF$buf2),
    .C(_3017__bF$buf3),
    .Y(_3041_)
);

AOI21X1 _13482_ (
    .A(_3040_),
    .B(_3014__bF$buf1),
    .C(_3041_),
    .Y(\datapath.csr._32_ [12])
);

OAI21X1 _13483_ (
    .A(\datapath.csr.csr_wdata [13]),
    .B(_3014__bF$buf0),
    .C(_3017__bF$buf2),
    .Y(_3042_)
);

AOI21X1 _13484_ (
    .A(_2817_),
    .B(_3014__bF$buf6),
    .C(_3042_),
    .Y(\datapath.csr._32_ [13])
);

OAI21X1 _13485_ (
    .A(\datapath.csr.csr_wdata [14]),
    .B(_3014__bF$buf5),
    .C(_3017__bF$buf1),
    .Y(_3043_)
);

AOI21X1 _13486_ (
    .A(_2819_),
    .B(_3014__bF$buf4),
    .C(_3043_),
    .Y(\datapath.csr._32_ [14])
);

OAI21X1 _13487_ (
    .A(\datapath.csr.csr_wdata [15]),
    .B(_3014__bF$buf3),
    .C(_3017__bF$buf0),
    .Y(_3044_)
);

AOI21X1 _13488_ (
    .A(_2821_),
    .B(_3014__bF$buf2),
    .C(_3044_),
    .Y(\datapath.csr._32_ [15])
);

OAI21X1 _13489_ (
    .A(\datapath.csr.csr_wdata [16]),
    .B(_3014__bF$buf1),
    .C(_3017__bF$buf4),
    .Y(_3045_)
);

AOI21X1 _13490_ (
    .A(_2823_),
    .B(_3014__bF$buf0),
    .C(_3045_),
    .Y(\datapath.csr._32_ [16])
);

OAI21X1 _13491_ (
    .A(\datapath.csr.csr_wdata [17]),
    .B(_3014__bF$buf6),
    .C(_3017__bF$buf3),
    .Y(_3046_)
);

AOI21X1 _13492_ (
    .A(_2825_),
    .B(_3014__bF$buf5),
    .C(_3046_),
    .Y(\datapath.csr._32_ [17])
);

OAI21X1 _13493_ (
    .A(\datapath.csr.csr_wdata [18]),
    .B(_3014__bF$buf4),
    .C(_3017__bF$buf2),
    .Y(_3047_)
);

AOI21X1 _13494_ (
    .A(_2827_),
    .B(_3014__bF$buf3),
    .C(_3047_),
    .Y(\datapath.csr._32_ [18])
);

OAI21X1 _13495_ (
    .A(\datapath.csr.csr_wdata [19]),
    .B(_3014__bF$buf2),
    .C(_3017__bF$buf1),
    .Y(_3048_)
);

AOI21X1 _13496_ (
    .A(_2829_),
    .B(_3014__bF$buf1),
    .C(_3048_),
    .Y(\datapath.csr._32_ [19])
);

OAI21X1 _13497_ (
    .A(\datapath.csr.csr_wdata [20]),
    .B(_3014__bF$buf0),
    .C(_3017__bF$buf0),
    .Y(_3049_)
);

AOI21X1 _13498_ (
    .A(_2831_),
    .B(_3014__bF$buf6),
    .C(_3049_),
    .Y(\datapath.csr._32_ [20])
);

OAI21X1 _13499_ (
    .A(\datapath.csr.csr_wdata [21]),
    .B(_3014__bF$buf5),
    .C(_3017__bF$buf4),
    .Y(_3050_)
);

AOI21X1 _13500_ (
    .A(_2833_),
    .B(_3014__bF$buf4),
    .C(_3050_),
    .Y(\datapath.csr._32_ [21])
);

OAI21X1 _13501_ (
    .A(\datapath.csr.csr_wdata [22]),
    .B(_3014__bF$buf3),
    .C(_3017__bF$buf3),
    .Y(_3051_)
);

AOI21X1 _13502_ (
    .A(_2835_),
    .B(_3014__bF$buf2),
    .C(_3051_),
    .Y(\datapath.csr._32_ [22])
);

OAI21X1 _13503_ (
    .A(\datapath.csr.csr_wdata [23]),
    .B(_3014__bF$buf1),
    .C(_3017__bF$buf2),
    .Y(_3052_)
);

AOI21X1 _13504_ (
    .A(_2837_),
    .B(_3014__bF$buf0),
    .C(_3052_),
    .Y(\datapath.csr._32_ [23])
);

OAI21X1 _13505_ (
    .A(\datapath.csr.csr_wdata [24]),
    .B(_3014__bF$buf6),
    .C(_3017__bF$buf1),
    .Y(_3053_)
);

AOI21X1 _13506_ (
    .A(_2839_),
    .B(_3014__bF$buf5),
    .C(_3053_),
    .Y(\datapath.csr._32_ [24])
);

OAI21X1 _13507_ (
    .A(\datapath.csr.csr_wdata [25]),
    .B(_3014__bF$buf4),
    .C(_3017__bF$buf0),
    .Y(_3054_)
);

AOI21X1 _13508_ (
    .A(_2841_),
    .B(_3014__bF$buf3),
    .C(_3054_),
    .Y(\datapath.csr._32_ [25])
);

OAI21X1 _13509_ (
    .A(\datapath.csr.csr_wdata [26]),
    .B(_3014__bF$buf2),
    .C(_3017__bF$buf4),
    .Y(_3055_)
);

AOI21X1 _13510_ (
    .A(_2843_),
    .B(_3014__bF$buf1),
    .C(_3055_),
    .Y(\datapath.csr._32_ [26])
);

OAI21X1 _13511_ (
    .A(\datapath.csr.csr_wdata [27]),
    .B(_3014__bF$buf0),
    .C(_3017__bF$buf3),
    .Y(_3056_)
);

AOI21X1 _13512_ (
    .A(_2845_),
    .B(_3014__bF$buf6),
    .C(_3056_),
    .Y(\datapath.csr._32_ [27])
);

OAI21X1 _13513_ (
    .A(\datapath.csr.csr_wdata [28]),
    .B(_3014__bF$buf5),
    .C(_3017__bF$buf2),
    .Y(_3057_)
);

AOI21X1 _13514_ (
    .A(_2847_),
    .B(_3014__bF$buf4),
    .C(_3057_),
    .Y(\datapath.csr._32_ [28])
);

OAI21X1 _13515_ (
    .A(\datapath.csr.csr_wdata [29]),
    .B(_3014__bF$buf3),
    .C(_3017__bF$buf1),
    .Y(_3058_)
);

AOI21X1 _13516_ (
    .A(_2849_),
    .B(_3014__bF$buf2),
    .C(_3058_),
    .Y(\datapath.csr._32_ [29])
);

INVX1 _13517_ (
    .A(\datapath.csr.mcause [30]),
    .Y(_3059_)
);

OAI21X1 _13518_ (
    .A(\datapath.csr.csr_wdata [30]),
    .B(_3014__bF$buf1),
    .C(_3017__bF$buf0),
    .Y(_3060_)
);

AOI21X1 _13519_ (
    .A(_3059_),
    .B(_3014__bF$buf0),
    .C(_3060_),
    .Y(\datapath.csr._32_ [30])
);

NAND3X1 _13520_ (
    .A(\datapath.csr.mcause [31]),
    .B(_3017__bF$buf4),
    .C(_3018_),
    .Y(_3061_)
);

OAI21X1 _13521_ (
    .A(_3017__bF$buf3),
    .B(_2575_),
    .C(_3061_),
    .Y(\datapath.csr._32_ [31])
);

AND2X2 _13522_ (
    .A(_2864_),
    .B(_2862_),
    .Y(_3062_)
);

NAND2X1 _13523_ (
    .A(_2915_),
    .B(_2921_),
    .Y(_3063_)
);

NOR2X1 _13524_ (
    .A(_2868_),
    .B(_3063_),
    .Y(_3064_)
);

NAND3X1 _13525_ (
    .A(\datapath.allowcsrwrite ),
    .B(_3062_),
    .C(_3064_),
    .Y(_2568_)
);

MUX2X1 _13526_ (
    .A(\datapath.csr.mstatus [0]),
    .B(\datapath.csr.csr_wdata [3]),
    .S(_2568_),
    .Y(_2569_)
);

OAI21X1 _13527_ (
    .A(\datapath.csr.mstatus [1]),
    .B(_2597__bF$buf3),
    .C(_3017__bF$buf2),
    .Y(_2570_)
);

AOI21X1 _13528_ (
    .A(_2569_),
    .B(_2597__bF$buf2),
    .C(_2570_),
    .Y(\datapath.csr._37_ [0])
);

INVX1 _13529_ (
    .A(\datapath.csr.mstatus [0]),
    .Y(_2571_)
);

NAND2X1 _13530_ (
    .A(\datapath.csr.mstatus [1]),
    .B(_2568_),
    .Y(_2572_)
);

OAI21X1 _13531_ (
    .A(_2878_),
    .B(_2568_),
    .C(_2572_),
    .Y(_2573_)
);

OAI21X1 _13532_ (
    .A(\controlunit.mret_bF$buf3 ),
    .B(_2573_),
    .C(_3017__bF$buf1),
    .Y(_2574_)
);

OAI21X1 _13533_ (
    .A(_2571_),
    .B(_3017__bF$buf0),
    .C(_2574_),
    .Y(\datapath.csr._37_ [1])
);

DFFPOSX1 _13534_ (
    .CLK(CLK_bF$buf26),
    .D(\datapath.csr._37_ [0]),
    .Q(\datapath.csr.mstatus [0])
);

DFFPOSX1 _13535_ (
    .CLK(CLK_bF$buf25),
    .D(\datapath.csr._37_ [1]),
    .Q(\datapath.csr.mstatus [1])
);

DFFPOSX1 _13536_ (
    .CLK(CLK_bF$buf24),
    .D(\datapath.csr._32_ [0]),
    .Q(\datapath.csr.mcause [0])
);

DFFPOSX1 _13537_ (
    .CLK(CLK_bF$buf23),
    .D(\datapath.csr._32_ [1]),
    .Q(\datapath.csr.mcause [1])
);

DFFPOSX1 _13538_ (
    .CLK(CLK_bF$buf22),
    .D(\datapath.csr._32_ [2]),
    .Q(\datapath.csr.mcause [2])
);

DFFPOSX1 _13539_ (
    .CLK(CLK_bF$buf21),
    .D(\datapath.csr._32_ [3]),
    .Q(\datapath.csr.mcause [3])
);

DFFPOSX1 _13540_ (
    .CLK(CLK_bF$buf20),
    .D(\datapath.csr._32_ [4]),
    .Q(\datapath.csr.mcause [4])
);

DFFPOSX1 _13541_ (
    .CLK(CLK_bF$buf19),
    .D(\datapath.csr._32_ [5]),
    .Q(\datapath.csr.mcause [5])
);

DFFPOSX1 _13542_ (
    .CLK(CLK_bF$buf18),
    .D(\datapath.csr._32_ [6]),
    .Q(\datapath.csr.mcause [6])
);

DFFPOSX1 _13543_ (
    .CLK(CLK_bF$buf17),
    .D(\datapath.csr._32_ [7]),
    .Q(\datapath.csr.mcause [7])
);

DFFPOSX1 _13544_ (
    .CLK(CLK_bF$buf16),
    .D(\datapath.csr._32_ [8]),
    .Q(\datapath.csr.mcause [8])
);

DFFPOSX1 _13545_ (
    .CLK(CLK_bF$buf15),
    .D(\datapath.csr._32_ [9]),
    .Q(\datapath.csr.mcause [9])
);

DFFPOSX1 _13546_ (
    .CLK(CLK_bF$buf14),
    .D(\datapath.csr._32_ [10]),
    .Q(\datapath.csr.mcause [10])
);

DFFPOSX1 _13547_ (
    .CLK(CLK_bF$buf13),
    .D(\datapath.csr._32_ [11]),
    .Q(\datapath.csr.mcause [11])
);

DFFPOSX1 _13548_ (
    .CLK(CLK_bF$buf12),
    .D(\datapath.csr._32_ [12]),
    .Q(\datapath.csr.mcause [12])
);

DFFPOSX1 _13549_ (
    .CLK(CLK_bF$buf11),
    .D(\datapath.csr._32_ [13]),
    .Q(\datapath.csr.mcause [13])
);

DFFPOSX1 _13550_ (
    .CLK(CLK_bF$buf10),
    .D(\datapath.csr._32_ [14]),
    .Q(\datapath.csr.mcause [14])
);

DFFPOSX1 _13551_ (
    .CLK(CLK_bF$buf9),
    .D(\datapath.csr._32_ [15]),
    .Q(\datapath.csr.mcause [15])
);

DFFPOSX1 _13552_ (
    .CLK(CLK_bF$buf8),
    .D(\datapath.csr._32_ [16]),
    .Q(\datapath.csr.mcause [16])
);

DFFPOSX1 _13553_ (
    .CLK(CLK_bF$buf7),
    .D(\datapath.csr._32_ [17]),
    .Q(\datapath.csr.mcause [17])
);

DFFPOSX1 _13554_ (
    .CLK(CLK_bF$buf6),
    .D(\datapath.csr._32_ [18]),
    .Q(\datapath.csr.mcause [18])
);

DFFPOSX1 _13555_ (
    .CLK(CLK_bF$buf5),
    .D(\datapath.csr._32_ [19]),
    .Q(\datapath.csr.mcause [19])
);

DFFPOSX1 _13556_ (
    .CLK(CLK_bF$buf4),
    .D(\datapath.csr._32_ [20]),
    .Q(\datapath.csr.mcause [20])
);

DFFPOSX1 _13557_ (
    .CLK(CLK_bF$buf3),
    .D(\datapath.csr._32_ [21]),
    .Q(\datapath.csr.mcause [21])
);

DFFPOSX1 _13558_ (
    .CLK(CLK_bF$buf2),
    .D(\datapath.csr._32_ [22]),
    .Q(\datapath.csr.mcause [22])
);

DFFPOSX1 _13559_ (
    .CLK(CLK_bF$buf1),
    .D(\datapath.csr._32_ [23]),
    .Q(\datapath.csr.mcause [23])
);

DFFPOSX1 _13560_ (
    .CLK(CLK_bF$buf0),
    .D(\datapath.csr._32_ [24]),
    .Q(\datapath.csr.mcause [24])
);

DFFPOSX1 _13561_ (
    .CLK(CLK_bF$buf151),
    .D(\datapath.csr._32_ [25]),
    .Q(\datapath.csr.mcause [25])
);

DFFPOSX1 _13562_ (
    .CLK(CLK_bF$buf150),
    .D(\datapath.csr._32_ [26]),
    .Q(\datapath.csr.mcause [26])
);

DFFPOSX1 _13563_ (
    .CLK(CLK_bF$buf149),
    .D(\datapath.csr._32_ [27]),
    .Q(\datapath.csr.mcause [27])
);

DFFPOSX1 _13564_ (
    .CLK(CLK_bF$buf148),
    .D(\datapath.csr._32_ [28]),
    .Q(\datapath.csr.mcause [28])
);

DFFPOSX1 _13565_ (
    .CLK(CLK_bF$buf147),
    .D(\datapath.csr._32_ [29]),
    .Q(\datapath.csr.mcause [29])
);

DFFPOSX1 _13566_ (
    .CLK(CLK_bF$buf146),
    .D(\datapath.csr._32_ [30]),
    .Q(\datapath.csr.mcause [30])
);

DFFPOSX1 _13567_ (
    .CLK(CLK_bF$buf145),
    .D(\datapath.csr._32_ [31]),
    .Q(\datapath.csr.mcause [31])
);

DFFPOSX1 _13568_ (
    .CLK(CLK_bF$buf144),
    .D(\datapath.csr._26_ [0]),
    .Q(\datapath.csr.mepc [0])
);

DFFPOSX1 _13569_ (
    .CLK(CLK_bF$buf143),
    .D(\datapath.csr._26_ [1]),
    .Q(\datapath.csr.mepc [1])
);

DFFPOSX1 _13570_ (
    .CLK(CLK_bF$buf142),
    .D(\datapath.csr._26_ [2]),
    .Q(\datapath.csr.mepc [2])
);

DFFPOSX1 _13571_ (
    .CLK(CLK_bF$buf141),
    .D(\datapath.csr._26_ [3]),
    .Q(\datapath.csr.mepc [3])
);

DFFPOSX1 _13572_ (
    .CLK(CLK_bF$buf140),
    .D(\datapath.csr._26_ [4]),
    .Q(\datapath.csr.mepc [4])
);

DFFPOSX1 _13573_ (
    .CLK(CLK_bF$buf139),
    .D(\datapath.csr._26_ [5]),
    .Q(\datapath.csr.mepc [5])
);

DFFPOSX1 _13574_ (
    .CLK(CLK_bF$buf138),
    .D(\datapath.csr._26_ [6]),
    .Q(\datapath.csr.mepc [6])
);

DFFPOSX1 _13575_ (
    .CLK(CLK_bF$buf137),
    .D(\datapath.csr._26_ [7]),
    .Q(\datapath.csr.mepc [7])
);

DFFPOSX1 _13576_ (
    .CLK(CLK_bF$buf136),
    .D(\datapath.csr._26_ [8]),
    .Q(\datapath.csr.mepc [8])
);

DFFPOSX1 _13577_ (
    .CLK(CLK_bF$buf135),
    .D(\datapath.csr._26_ [9]),
    .Q(\datapath.csr.mepc [9])
);

DFFPOSX1 _13578_ (
    .CLK(CLK_bF$buf134),
    .D(\datapath.csr._26_ [10]),
    .Q(\datapath.csr.mepc [10])
);

DFFPOSX1 _13579_ (
    .CLK(CLK_bF$buf133),
    .D(\datapath.csr._26_ [11]),
    .Q(\datapath.csr.mepc [11])
);

DFFPOSX1 _13580_ (
    .CLK(CLK_bF$buf132),
    .D(\datapath.csr._26_ [12]),
    .Q(\datapath.csr.mepc [12])
);

DFFPOSX1 _13581_ (
    .CLK(CLK_bF$buf131),
    .D(\datapath.csr._26_ [13]),
    .Q(\datapath.csr.mepc [13])
);

DFFPOSX1 _13582_ (
    .CLK(CLK_bF$buf130),
    .D(\datapath.csr._26_ [14]),
    .Q(\datapath.csr.mepc [14])
);

DFFPOSX1 _13583_ (
    .CLK(CLK_bF$buf129),
    .D(\datapath.csr._26_ [15]),
    .Q(\datapath.csr.mepc [15])
);

DFFPOSX1 _13584_ (
    .CLK(CLK_bF$buf128),
    .D(\datapath.csr._26_ [16]),
    .Q(\datapath.csr.mepc [16])
);

DFFPOSX1 _13585_ (
    .CLK(CLK_bF$buf127),
    .D(\datapath.csr._26_ [17]),
    .Q(\datapath.csr.mepc [17])
);

DFFPOSX1 _13586_ (
    .CLK(CLK_bF$buf126),
    .D(\datapath.csr._26_ [18]),
    .Q(\datapath.csr.mepc [18])
);

DFFPOSX1 _13587_ (
    .CLK(CLK_bF$buf125),
    .D(\datapath.csr._26_ [19]),
    .Q(\datapath.csr.mepc [19])
);

DFFPOSX1 _13588_ (
    .CLK(CLK_bF$buf124),
    .D(\datapath.csr._26_ [20]),
    .Q(\datapath.csr.mepc [20])
);

DFFPOSX1 _13589_ (
    .CLK(CLK_bF$buf123),
    .D(\datapath.csr._26_ [21]),
    .Q(\datapath.csr.mepc [21])
);

DFFPOSX1 _13590_ (
    .CLK(CLK_bF$buf122),
    .D(\datapath.csr._26_ [22]),
    .Q(\datapath.csr.mepc [22])
);

DFFPOSX1 _13591_ (
    .CLK(CLK_bF$buf121),
    .D(\datapath.csr._26_ [23]),
    .Q(\datapath.csr.mepc [23])
);

DFFPOSX1 _13592_ (
    .CLK(CLK_bF$buf120),
    .D(\datapath.csr._26_ [24]),
    .Q(\datapath.csr.mepc [24])
);

DFFPOSX1 _13593_ (
    .CLK(CLK_bF$buf119),
    .D(\datapath.csr._26_ [25]),
    .Q(\datapath.csr.mepc [25])
);

DFFPOSX1 _13594_ (
    .CLK(CLK_bF$buf118),
    .D(\datapath.csr._26_ [26]),
    .Q(\datapath.csr.mepc [26])
);

DFFPOSX1 _13595_ (
    .CLK(CLK_bF$buf117),
    .D(\datapath.csr._26_ [27]),
    .Q(\datapath.csr.mepc [27])
);

DFFPOSX1 _13596_ (
    .CLK(CLK_bF$buf116),
    .D(\datapath.csr._26_ [28]),
    .Q(\datapath.csr.mepc [28])
);

DFFPOSX1 _13597_ (
    .CLK(CLK_bF$buf115),
    .D(\datapath.csr._26_ [29]),
    .Q(\datapath.csr.mepc [29])
);

DFFPOSX1 _13598_ (
    .CLK(CLK_bF$buf114),
    .D(IRQ),
    .Q(\datapath.csr.meta_irq )
);

DFFPOSX1 _13599_ (
    .CLK(CLK_bF$buf113),
    .D(\datapath.csr.meta_irq ),
    .Q(\datapath.csr.mip )
);

DFFPOSX1 _13600_ (
    .CLK(CLK_bF$buf112),
    .D(\datapath.csr._20_ ),
    .Q(\datapath.csr.mie )
);

DFFPOSX1 _13601_ (
    .CLK(CLK_bF$buf111),
    .D(\datapath.csr._13_ [0]),
    .Q(\datapath.csr.mvect [0])
);

DFFPOSX1 _13602_ (
    .CLK(CLK_bF$buf110),
    .D(\datapath.csr._13_ [1]),
    .Q(\datapath.csr.mvect [1])
);

DFFPOSX1 _13603_ (
    .CLK(CLK_bF$buf109),
    .D(\datapath.csr._13_ [2]),
    .Q(\datapath.csr.mvect [2])
);

DFFPOSX1 _13604_ (
    .CLK(CLK_bF$buf108),
    .D(\datapath.csr._13_ [3]),
    .Q(\datapath.csr.mvect [3])
);

DFFPOSX1 _13605_ (
    .CLK(CLK_bF$buf107),
    .D(\datapath.csr._13_ [4]),
    .Q(\datapath.csr.mvect [4])
);

DFFPOSX1 _13606_ (
    .CLK(CLK_bF$buf106),
    .D(\datapath.csr._13_ [5]),
    .Q(\datapath.csr.mvect [5])
);

DFFPOSX1 _13607_ (
    .CLK(CLK_bF$buf105),
    .D(\datapath.csr._13_ [6]),
    .Q(\datapath.csr.mvect [6])
);

DFFPOSX1 _13608_ (
    .CLK(CLK_bF$buf104),
    .D(\datapath.csr._13_ [7]),
    .Q(\datapath.csr.mvect [7])
);

DFFPOSX1 _13609_ (
    .CLK(CLK_bF$buf103),
    .D(\datapath.csr._13_ [8]),
    .Q(\datapath.csr.mvect [8])
);

DFFPOSX1 _13610_ (
    .CLK(CLK_bF$buf102),
    .D(\datapath.csr._13_ [9]),
    .Q(\datapath.csr.mvect [9])
);

DFFPOSX1 _13611_ (
    .CLK(CLK_bF$buf101),
    .D(\datapath.csr._13_ [10]),
    .Q(\datapath.csr.mvect [10])
);

DFFPOSX1 _13612_ (
    .CLK(CLK_bF$buf100),
    .D(\datapath.csr._13_ [11]),
    .Q(\datapath.csr.mvect [11])
);

DFFPOSX1 _13613_ (
    .CLK(CLK_bF$buf99),
    .D(\datapath.csr._13_ [12]),
    .Q(\datapath.csr.mvect [12])
);

DFFPOSX1 _13614_ (
    .CLK(CLK_bF$buf98),
    .D(\datapath.csr._13_ [13]),
    .Q(\datapath.csr.mvect [13])
);

DFFPOSX1 _13615_ (
    .CLK(CLK_bF$buf97),
    .D(\datapath.csr._13_ [14]),
    .Q(\datapath.csr.mvect [14])
);

DFFPOSX1 _13616_ (
    .CLK(CLK_bF$buf96),
    .D(\datapath.csr._13_ [15]),
    .Q(\datapath.csr.mvect [15])
);

DFFPOSX1 _13617_ (
    .CLK(CLK_bF$buf95),
    .D(\datapath.csr._13_ [16]),
    .Q(\datapath.csr.mvect [16])
);

DFFPOSX1 _13618_ (
    .CLK(CLK_bF$buf94),
    .D(\datapath.csr._13_ [17]),
    .Q(\datapath.csr.mvect [17])
);

DFFPOSX1 _13619_ (
    .CLK(CLK_bF$buf93),
    .D(\datapath.csr._13_ [18]),
    .Q(\datapath.csr.mvect [18])
);

DFFPOSX1 _13620_ (
    .CLK(CLK_bF$buf92),
    .D(\datapath.csr._13_ [19]),
    .Q(\datapath.csr.mvect [19])
);

DFFPOSX1 _13621_ (
    .CLK(CLK_bF$buf91),
    .D(\datapath.csr._13_ [20]),
    .Q(\datapath.csr.mvect [20])
);

DFFPOSX1 _13622_ (
    .CLK(CLK_bF$buf90),
    .D(\datapath.csr._13_ [21]),
    .Q(\datapath.csr.mvect [21])
);

DFFPOSX1 _13623_ (
    .CLK(CLK_bF$buf89),
    .D(\datapath.csr._13_ [22]),
    .Q(\datapath.csr.mvect [22])
);

DFFPOSX1 _13624_ (
    .CLK(CLK_bF$buf88),
    .D(\datapath.csr._13_ [23]),
    .Q(\datapath.csr.mvect [23])
);

DFFPOSX1 _13625_ (
    .CLK(CLK_bF$buf87),
    .D(\datapath.csr._13_ [24]),
    .Q(\datapath.csr.mvect [24])
);

DFFPOSX1 _13626_ (
    .CLK(CLK_bF$buf86),
    .D(\datapath.csr._13_ [25]),
    .Q(\datapath.csr.mvect [25])
);

DFFPOSX1 _13627_ (
    .CLK(CLK_bF$buf85),
    .D(\datapath.csr._13_ [26]),
    .Q(\datapath.csr.mvect [26])
);

DFFPOSX1 _13628_ (
    .CLK(CLK_bF$buf84),
    .D(\datapath.csr._13_ [27]),
    .Q(\datapath.csr.mvect [27])
);

DFFPOSX1 _13629_ (
    .CLK(CLK_bF$buf83),
    .D(\datapath.csr._13_ [28]),
    .Q(\datapath.csr.mvect [28])
);

DFFPOSX1 _13630_ (
    .CLK(CLK_bF$buf82),
    .D(\datapath.csr._13_ [29]),
    .Q(\datapath.csr.mvect [29])
);

DFFPOSX1 _13631_ (
    .CLK(CLK_bF$buf81),
    .D(\datapath.csr._13_ [30]),
    .Q(\datapath.csr.mvect [30])
);

DFFPOSX1 _13632_ (
    .CLK(CLK_bF$buf80),
    .D(\datapath.csr._13_ [31]),
    .Q(\datapath.csr.mvect [31])
);

INVX2 _13633_ (
    .A(\controlunit.imm_sel [2]),
    .Y(_3101_)
);

NAND3X1 _13634_ (
    .A(\controlunit.imm_sel [1]),
    .B(\controlunit.imm_sel [0]),
    .C(_3101_),
    .Y(_3102_)
);

INVX2 _13635_ (
    .A(\controlunit.imm_sel [1]),
    .Y(_3103_)
);

NAND3X1 _13636_ (
    .A(\controlunit.imm_sel [0]),
    .B(\controlunit.imm_sel [2]),
    .C(_3103_),
    .Y(_3104_)
);

AND2X2 _13637_ (
    .A(_3102_),
    .B(_3104_),
    .Y(_3105_)
);

NAND2X1 _13638_ (
    .A(\datapath.idinstr [25]),
    .B(_3105_),
    .Y(_3106_)
);

INVX1 _13639_ (
    .A(_3106_),
    .Y(\datapath.imm [5])
);

NAND2X1 _13640_ (
    .A(\datapath.idinstr [26]),
    .B(_3105_),
    .Y(_3107_)
);

INVX1 _13641_ (
    .A(_3107_),
    .Y(\datapath.imm [6])
);

NAND2X1 _13642_ (
    .A(\datapath.idinstr [27]),
    .B(_3105_),
    .Y(_3108_)
);

INVX1 _13643_ (
    .A(_3108_),
    .Y(\datapath.imm [7])
);

NAND2X1 _13644_ (
    .A(\datapath.idinstr [28]),
    .B(_3105_),
    .Y(_3109_)
);

INVX1 _13645_ (
    .A(_3109_),
    .Y(\datapath.imm [8])
);

NAND2X1 _13646_ (
    .A(\datapath.idinstr [29]),
    .B(_3105_),
    .Y(_3110_)
);

INVX1 _13647_ (
    .A(_3110_),
    .Y(\datapath.imm [9])
);

NAND2X1 _13648_ (
    .A(\datapath.idinstr [30]),
    .B(_3105_),
    .Y(_3111_)
);

INVX1 _13649_ (
    .A(_3111_),
    .Y(\datapath.imm [10])
);

NAND2X1 _13650_ (
    .A(\datapath.idinstr [31]),
    .B(_3104_),
    .Y(_3112_)
);

INVX1 _13651_ (
    .A(_3112_),
    .Y(\datapath.immediatedecoder._12_ )
);

INVX1 _13652_ (
    .A(\datapath.idinstr [31]),
    .Y(_3113_)
);

INVX2 _13653_ (
    .A(\controlunit.imm_sel [0]),
    .Y(_3114_)
);

NAND3X1 _13654_ (
    .A(\controlunit.imm_sel [1]),
    .B(_3114_),
    .C(_3101_),
    .Y(_3115_)
);

AND2X2 _13655_ (
    .A(\controlunit.imm_sel [1]),
    .B(\controlunit.imm_sel [0]),
    .Y(_3116_)
);

OAI21X1 _13656_ (
    .A(\controlunit.imm_sel [1]),
    .B(\controlunit.imm_sel [0]),
    .C(\controlunit.imm_sel [2]),
    .Y(_3117_)
);

OAI21X1 _13657_ (
    .A(\controlunit.imm_sel [2]),
    .B(_3116_),
    .C(_3117_),
    .Y(_3118_)
);

NAND3X1 _13658_ (
    .A(_3104_),
    .B(_3115_),
    .C(_3118_),
    .Y(_3119_)
);

NOR3X1 _13659_ (
    .A(\controlunit.imm_sel [0]),
    .B(\controlunit.imm_sel [2]),
    .C(_3103_),
    .Y(_3120_)
);

NOR2X1 _13660_ (
    .A(\controlunit.imm_sel [1]),
    .B(\controlunit.imm_sel [0]),
    .Y(_3121_)
);

AND2X2 _13661_ (
    .A(_3121_),
    .B(\controlunit.imm_sel [2]),
    .Y(_3122_)
);

AOI22X1 _13662_ (
    .A(\datapath.idinstr [7]),
    .B(_3120_),
    .C(\datapath.idinstr_20_bF$buf52 ),
    .D(_3122_),
    .Y(_3123_)
);

OAI21X1 _13663_ (
    .A(_3113_),
    .B(_3119_),
    .C(_3123_),
    .Y(\datapath.immediatedecoder._09_ )
);

OAI21X1 _13664_ (
    .A(\controlunit.imm_sel [2]),
    .B(_3114_),
    .C(_3103_),
    .Y(_3124_)
);

NAND3X1 _13665_ (
    .A(\datapath.idinstr [8]),
    .B(_3102_),
    .C(_3124_),
    .Y(_3125_)
);

INVX2 _13666_ (
    .A(_3104_),
    .Y(_3126_)
);

NAND2X1 _13667_ (
    .A(\datapath.idinstr_16_bF$buf50 ),
    .B(_3126_),
    .Y(_3127_)
);

NAND2X1 _13668_ (
    .A(\datapath.idinstr_21_bF$buf47 ),
    .B(_3121_),
    .Y(_3128_)
);

NAND3X1 _13669_ (
    .A(_3125_),
    .B(_3128_),
    .C(_3127_),
    .Y(\datapath.imm [1])
);

NAND3X1 _13670_ (
    .A(\datapath.idinstr [9]),
    .B(_3102_),
    .C(_3124_),
    .Y(_3129_)
);

NAND2X1 _13671_ (
    .A(\datapath.idinstr_17_bF$buf14 ),
    .B(_3126_),
    .Y(_3130_)
);

NAND2X1 _13672_ (
    .A(\datapath.idinstr_22_bF$buf37 ),
    .B(_3121_),
    .Y(_3065_)
);

NAND3X1 _13673_ (
    .A(_3129_),
    .B(_3065_),
    .C(_3130_),
    .Y(\datapath.imm [2])
);

NAND3X1 _13674_ (
    .A(\datapath.idinstr [10]),
    .B(_3102_),
    .C(_3124_),
    .Y(_3066_)
);

NAND2X1 _13675_ (
    .A(\datapath.idinstr_18_bF$buf5 ),
    .B(_3126_),
    .Y(_3067_)
);

NAND2X1 _13676_ (
    .A(\datapath.idinstr_23_bF$buf3 ),
    .B(_3121_),
    .Y(_3068_)
);

NAND3X1 _13677_ (
    .A(_3066_),
    .B(_3068_),
    .C(_3067_),
    .Y(\datapath.imm [3])
);

NAND3X1 _13678_ (
    .A(\datapath.idinstr [11]),
    .B(_3102_),
    .C(_3124_),
    .Y(_3069_)
);

NAND2X1 _13679_ (
    .A(\datapath.idinstr_19_bF$buf4 ),
    .B(_3126_),
    .Y(_3070_)
);

NAND2X1 _13680_ (
    .A(\datapath.idinstr_24_bF$buf3 ),
    .B(_3121_),
    .Y(_3071_)
);

NAND3X1 _13681_ (
    .A(_3069_),
    .B(_3071_),
    .C(_3070_),
    .Y(\datapath.imm [4])
);

NAND3X1 _13682_ (
    .A(\controlunit.imm_sel [0]),
    .B(_3103_),
    .C(_3101_),
    .Y(_3072_)
);

NAND2X1 _13683_ (
    .A(\datapath.idinstr_20_bF$buf51 ),
    .B(_3072_),
    .Y(_3073_)
);

NOR3X1 _13684_ (
    .A(\controlunit.imm_sel [1]),
    .B(\controlunit.imm_sel [2]),
    .C(_3114_),
    .Y(_3074_)
);

AOI22X1 _13685_ (
    .A(\datapath.idinstr [7]),
    .B(_3074_),
    .C(\datapath.idinstr_15_bF$buf53 ),
    .D(_3126_),
    .Y(_3075_)
);

OAI21X1 _13686_ (
    .A(_3073_),
    .B(_3119_),
    .C(_3075_),
    .Y(\datapath.immediatedecoder._06_ )
);

INVX1 _13687_ (
    .A(\datapath.idinstr_20_bF$buf50 ),
    .Y(_3076_)
);

OAI21X1 _13688_ (
    .A(_3103_),
    .B(_3101_),
    .C(_3114_),
    .Y(_3077_)
);

NAND2X1 _13689_ (
    .A(_3072_),
    .B(_3077_),
    .Y(_3078_)
);

NAND2X1 _13690_ (
    .A(\datapath.idinstr [31]),
    .B(_3078_),
    .Y(_3079_)
);

OAI21X1 _13691_ (
    .A(\controlunit.imm_sel [0]),
    .B(\controlunit.imm_sel [2]),
    .C(\controlunit.imm_sel [1]),
    .Y(_3080_)
);

OAI21X1 _13692_ (
    .A(_3076_),
    .B(_3080_),
    .C(_3079_),
    .Y(\datapath.imm [20])
);

INVX1 _13693_ (
    .A(\datapath.idinstr_21_bF$buf46 ),
    .Y(_3081_)
);

OAI21X1 _13694_ (
    .A(_3081_),
    .B(_3080_),
    .C(_3079_),
    .Y(\datapath.imm [21])
);

INVX1 _13695_ (
    .A(\datapath.idinstr_22_bF$buf36 ),
    .Y(_3082_)
);

OAI21X1 _13696_ (
    .A(_3082_),
    .B(_3080_),
    .C(_3079_),
    .Y(\datapath.imm [22])
);

INVX1 _13697_ (
    .A(\datapath.idinstr_23_bF$buf2 ),
    .Y(_3083_)
);

OAI21X1 _13698_ (
    .A(_3083_),
    .B(_3080_),
    .C(_3079_),
    .Y(\datapath.imm [23])
);

INVX1 _13699_ (
    .A(\datapath.idinstr_24_bF$buf2 ),
    .Y(_3084_)
);

OAI21X1 _13700_ (
    .A(_3084_),
    .B(_3080_),
    .C(_3079_),
    .Y(\datapath.imm [24])
);

INVX1 _13701_ (
    .A(\datapath.idinstr [25]),
    .Y(_3085_)
);

OAI21X1 _13702_ (
    .A(_3085_),
    .B(_3080_),
    .C(_3079_),
    .Y(\datapath.imm [25])
);

INVX1 _13703_ (
    .A(\datapath.idinstr [26]),
    .Y(_3086_)
);

OAI21X1 _13704_ (
    .A(_3086_),
    .B(_3080_),
    .C(_3079_),
    .Y(\datapath.imm [26])
);

INVX1 _13705_ (
    .A(\datapath.idinstr [27]),
    .Y(_3087_)
);

OAI21X1 _13706_ (
    .A(_3087_),
    .B(_3080_),
    .C(_3079_),
    .Y(\datapath.imm [27])
);

INVX1 _13707_ (
    .A(\datapath.idinstr [28]),
    .Y(_3088_)
);

OAI21X1 _13708_ (
    .A(_3088_),
    .B(_3080_),
    .C(_3079_),
    .Y(\datapath.imm [28])
);

INVX1 _13709_ (
    .A(\datapath.idinstr [29]),
    .Y(_3089_)
);

OAI21X1 _13710_ (
    .A(_3089_),
    .B(_3080_),
    .C(_3079_),
    .Y(\datapath.imm [29])
);

INVX1 _13711_ (
    .A(\datapath.idinstr [30]),
    .Y(_3090_)
);

OAI21X1 _13712_ (
    .A(_3090_),
    .B(_3080_),
    .C(_3079_),
    .Y(\datapath.imm [30])
);

NAND2X1 _13713_ (
    .A(_3103_),
    .B(_3114_),
    .Y(_3091_)
);

OAI21X1 _13714_ (
    .A(_3101_),
    .B(_3091_),
    .C(_3102_),
    .Y(_3092_)
);

NAND2X1 _13715_ (
    .A(\datapath.idinstr [12]),
    .B(_3092_),
    .Y(_3093_)
);

OAI21X1 _13716_ (
    .A(_3112_),
    .B(_3092_),
    .C(_3093_),
    .Y(\datapath.imm [12])
);

NAND2X1 _13717_ (
    .A(\datapath.idinstr [13]),
    .B(_3092_),
    .Y(_3094_)
);

OAI21X1 _13718_ (
    .A(_3112_),
    .B(_3092_),
    .C(_3094_),
    .Y(\datapath.imm [13])
);

NAND2X1 _13719_ (
    .A(\datapath.idinstr [14]),
    .B(_3092_),
    .Y(_3095_)
);

OAI21X1 _13720_ (
    .A(_3112_),
    .B(_3092_),
    .C(_3095_),
    .Y(\datapath.imm [14])
);

NAND2X1 _13721_ (
    .A(\datapath.idinstr_15_bF$buf52 ),
    .B(_3092_),
    .Y(_3096_)
);

OAI21X1 _13722_ (
    .A(_3112_),
    .B(_3092_),
    .C(_3096_),
    .Y(\datapath.imm [15])
);

NAND2X1 _13723_ (
    .A(\datapath.idinstr_16_bF$buf49 ),
    .B(_3092_),
    .Y(_3097_)
);

OAI21X1 _13724_ (
    .A(_3112_),
    .B(_3092_),
    .C(_3097_),
    .Y(\datapath.imm [16])
);

NAND2X1 _13725_ (
    .A(\datapath.idinstr_17_bF$buf13 ),
    .B(_3092_),
    .Y(_3098_)
);

OAI21X1 _13726_ (
    .A(_3112_),
    .B(_3092_),
    .C(_3098_),
    .Y(\datapath.imm [17])
);

NAND2X1 _13727_ (
    .A(\datapath.idinstr_18_bF$buf4 ),
    .B(_3092_),
    .Y(_3099_)
);

OAI21X1 _13728_ (
    .A(_3112_),
    .B(_3092_),
    .C(_3099_),
    .Y(\datapath.imm [18])
);

NAND2X1 _13729_ (
    .A(\datapath.idinstr_19_bF$buf3 ),
    .B(_3092_),
    .Y(_3100_)
);

OAI21X1 _13730_ (
    .A(_3112_),
    .B(_3092_),
    .C(_3100_),
    .Y(\datapath.imm [19])
);

INVX1 _13731_ (
    .A(\datapath.meminstr [12]),
    .Y(_3131_)
);

NAND2X1 _13732_ (
    .A(\datapath.meminstr [13]),
    .B(_3131_),
    .Y(_3132_)
);

INVX1 _13733_ (
    .A(\datapath.meminstr [13]),
    .Y(_3133_)
);

NAND2X1 _13734_ (
    .A(\datapath.meminstr [12]),
    .B(_3133_),
    .Y(_3134_)
);

NAND3X1 _13735_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [0]),
    .B(_3132__bF$buf5),
    .C(_3134__bF$buf5),
    .Y(_3135_)
);

NOR2X1 _13736_ (
    .A(\datapath.meminstr [12]),
    .B(_3133_),
    .Y(_3136_)
);

NAND2X1 _13737_ (
    .A(\datapath.memoryinterface.data_store [0]),
    .B(_3136__bF$buf7),
    .Y(_3137_)
);

NOR2X1 _13738_ (
    .A(\datapath.meminstr [13]),
    .B(_3131_),
    .Y(_3138_)
);

INVX1 _13739_ (
    .A(\datapath.memoryinterface.data_store [0]),
    .Y(_3139_)
);

NAND2X1 _13740_ (
    .A(DMEM_DATA_L[0]),
    .B(_0__1_bF$buf9),
    .Y(_3140_)
);

OAI21X1 _13741_ (
    .A(_0__1_bF$buf8),
    .B(_3139_),
    .C(_3140_),
    .Y(_3141_)
);

NAND2X1 _13742_ (
    .A(_3138__bF$buf6),
    .B(_3141_),
    .Y(_3142_)
);

NAND3X1 _13743_ (
    .A(_3137_),
    .B(_3135_),
    .C(_3142_),
    .Y(_1_[0])
);

NAND3X1 _13744_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [1]),
    .B(_3132__bF$buf4),
    .C(_3134__bF$buf4),
    .Y(_3143_)
);

NAND2X1 _13745_ (
    .A(\datapath.memoryinterface.data_store [1]),
    .B(_3136__bF$buf6),
    .Y(_3144_)
);

INVX1 _13746_ (
    .A(\datapath.memoryinterface.data_store [1]),
    .Y(_3145_)
);

NAND2X1 _13747_ (
    .A(_0__1_bF$buf7),
    .B(DMEM_DATA_L[1]),
    .Y(_3146_)
);

OAI21X1 _13748_ (
    .A(_0__1_bF$buf6),
    .B(_3145_),
    .C(_3146_),
    .Y(_3147_)
);

NAND2X1 _13749_ (
    .A(_3138__bF$buf5),
    .B(_3147_),
    .Y(_3148_)
);

NAND3X1 _13750_ (
    .A(_3144_),
    .B(_3143_),
    .C(_3148_),
    .Y(_1_[1])
);

NAND3X1 _13751_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [2]),
    .B(_3132__bF$buf3),
    .C(_3134__bF$buf3),
    .Y(_3149_)
);

NAND2X1 _13752_ (
    .A(\datapath.memoryinterface.data_store [2]),
    .B(_3136__bF$buf5),
    .Y(_3150_)
);

INVX1 _13753_ (
    .A(\datapath.memoryinterface.data_store [2]),
    .Y(_3151_)
);

NAND2X1 _13754_ (
    .A(_0__1_bF$buf5),
    .B(DMEM_DATA_L[2]),
    .Y(_3152_)
);

OAI21X1 _13755_ (
    .A(_0__1_bF$buf4),
    .B(_3151_),
    .C(_3152_),
    .Y(_3153_)
);

NAND2X1 _13756_ (
    .A(_3138__bF$buf4),
    .B(_3153_),
    .Y(_3154_)
);

NAND3X1 _13757_ (
    .A(_3150_),
    .B(_3149_),
    .C(_3154_),
    .Y(_1_[2])
);

NAND3X1 _13758_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [3]),
    .B(_3132__bF$buf2),
    .C(_3134__bF$buf2),
    .Y(_3155_)
);

NAND2X1 _13759_ (
    .A(\datapath.memoryinterface.data_store [3]),
    .B(_3136__bF$buf4),
    .Y(_3156_)
);

INVX1 _13760_ (
    .A(\datapath.memoryinterface.data_store [3]),
    .Y(_3157_)
);

NAND2X1 _13761_ (
    .A(_0__1_bF$buf3),
    .B(DMEM_DATA_L[3]),
    .Y(_3158_)
);

OAI21X1 _13762_ (
    .A(_0__1_bF$buf2),
    .B(_3157_),
    .C(_3158_),
    .Y(_3159_)
);

NAND2X1 _13763_ (
    .A(_3138__bF$buf3),
    .B(_3159_),
    .Y(_3160_)
);

NAND3X1 _13764_ (
    .A(_3156_),
    .B(_3155_),
    .C(_3160_),
    .Y(_1_[3])
);

NAND3X1 _13765_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [4]),
    .B(_3132__bF$buf1),
    .C(_3134__bF$buf1),
    .Y(_3161_)
);

NAND2X1 _13766_ (
    .A(\datapath.memoryinterface.data_store [4]),
    .B(_3136__bF$buf3),
    .Y(_3162_)
);

INVX1 _13767_ (
    .A(\datapath.memoryinterface.data_store [4]),
    .Y(_3163_)
);

NAND2X1 _13768_ (
    .A(_0__1_bF$buf1),
    .B(DMEM_DATA_L[4]),
    .Y(_3164_)
);

OAI21X1 _13769_ (
    .A(_0__1_bF$buf0),
    .B(_3163_),
    .C(_3164_),
    .Y(_3165_)
);

NAND2X1 _13770_ (
    .A(_3138__bF$buf2),
    .B(_3165_),
    .Y(_3166_)
);

NAND3X1 _13771_ (
    .A(_3162_),
    .B(_3161_),
    .C(_3166_),
    .Y(_1_[4])
);

NAND3X1 _13772_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [5]),
    .B(_3132__bF$buf0),
    .C(_3134__bF$buf0),
    .Y(_3167_)
);

NAND2X1 _13773_ (
    .A(\datapath.memoryinterface.data_store [5]),
    .B(_3136__bF$buf2),
    .Y(_3168_)
);

INVX1 _13774_ (
    .A(\datapath.memoryinterface.data_store [5]),
    .Y(_3169_)
);

NAND2X1 _13775_ (
    .A(_0__1_bF$buf10),
    .B(DMEM_DATA_L[5]),
    .Y(_3170_)
);

OAI21X1 _13776_ (
    .A(_0__1_bF$buf9),
    .B(_3169_),
    .C(_3170_),
    .Y(_3171_)
);

NAND2X1 _13777_ (
    .A(_3138__bF$buf1),
    .B(_3171_),
    .Y(_3172_)
);

NAND3X1 _13778_ (
    .A(_3168_),
    .B(_3167_),
    .C(_3172_),
    .Y(_1_[5])
);

NAND3X1 _13779_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [6]),
    .B(_3132__bF$buf5),
    .C(_3134__bF$buf5),
    .Y(_3173_)
);

NAND2X1 _13780_ (
    .A(\datapath.memoryinterface.data_store [6]),
    .B(_3136__bF$buf1),
    .Y(_3174_)
);

INVX1 _13781_ (
    .A(\datapath.memoryinterface.data_store [6]),
    .Y(_3175_)
);

NAND2X1 _13782_ (
    .A(_0__1_bF$buf8),
    .B(DMEM_DATA_L[6]),
    .Y(_3176_)
);

OAI21X1 _13783_ (
    .A(_0__1_bF$buf7),
    .B(_3175_),
    .C(_3176_),
    .Y(_3177_)
);

NAND2X1 _13784_ (
    .A(_3138__bF$buf0),
    .B(_3177_),
    .Y(_3178_)
);

NAND3X1 _13785_ (
    .A(_3174_),
    .B(_3173_),
    .C(_3178_),
    .Y(_1_[6])
);

NAND3X1 _13786_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [7]),
    .B(_3132__bF$buf4),
    .C(_3134__bF$buf4),
    .Y(_3179_)
);

NAND2X1 _13787_ (
    .A(\datapath.memoryinterface.data_store [7]),
    .B(_3136__bF$buf0),
    .Y(_3180_)
);

INVX1 _13788_ (
    .A(\datapath.memoryinterface.data_store [7]),
    .Y(_3181_)
);

NAND2X1 _13789_ (
    .A(_0__1_bF$buf6),
    .B(DMEM_DATA_L[7]),
    .Y(_3182_)
);

OAI21X1 _13790_ (
    .A(_0__1_bF$buf5),
    .B(_3181_),
    .C(_3182_),
    .Y(_3183_)
);

NAND2X1 _13791_ (
    .A(_3138__bF$buf6),
    .B(_3183_),
    .Y(_3184_)
);

NAND3X1 _13792_ (
    .A(_3180_),
    .B(_3179_),
    .C(_3184_),
    .Y(_1_[7])
);

NAND3X1 _13793_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [8]),
    .B(_3132__bF$buf3),
    .C(_3134__bF$buf3),
    .Y(_3185_)
);

NAND2X1 _13794_ (
    .A(\datapath.memoryinterface.data_store [8]),
    .B(_3136__bF$buf7),
    .Y(_3186_)
);

INVX1 _13795_ (
    .A(\datapath.memoryinterface.data_store [8]),
    .Y(_3187_)
);

NAND2X1 _13796_ (
    .A(_0__1_bF$buf4),
    .B(DMEM_DATA_L[8]),
    .Y(_3188_)
);

OAI21X1 _13797_ (
    .A(_0__1_bF$buf3),
    .B(_3187_),
    .C(_3188_),
    .Y(_3189_)
);

NAND2X1 _13798_ (
    .A(_3138__bF$buf5),
    .B(_3189_),
    .Y(_3190_)
);

NAND3X1 _13799_ (
    .A(_3186_),
    .B(_3185_),
    .C(_3190_),
    .Y(_1_[8])
);

NAND3X1 _13800_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [9]),
    .B(_3132__bF$buf2),
    .C(_3134__bF$buf2),
    .Y(_3191_)
);

NAND2X1 _13801_ (
    .A(\datapath.memoryinterface.data_store [9]),
    .B(_3136__bF$buf6),
    .Y(_3192_)
);

INVX1 _13802_ (
    .A(\datapath.memoryinterface.data_store [9]),
    .Y(_3193_)
);

NAND2X1 _13803_ (
    .A(_0__1_bF$buf2),
    .B(DMEM_DATA_L[9]),
    .Y(_3194_)
);

OAI21X1 _13804_ (
    .A(_0__1_bF$buf1),
    .B(_3193_),
    .C(_3194_),
    .Y(_3195_)
);

NAND2X1 _13805_ (
    .A(_3138__bF$buf4),
    .B(_3195_),
    .Y(_3196_)
);

NAND3X1 _13806_ (
    .A(_3192_),
    .B(_3191_),
    .C(_3196_),
    .Y(_1_[9])
);

NAND3X1 _13807_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [10]),
    .B(_3132__bF$buf1),
    .C(_3134__bF$buf1),
    .Y(_3197_)
);

NAND2X1 _13808_ (
    .A(\datapath.memoryinterface.data_store [10]),
    .B(_3136__bF$buf5),
    .Y(_3198_)
);

INVX1 _13809_ (
    .A(\datapath.memoryinterface.data_store [10]),
    .Y(_3199_)
);

NAND2X1 _13810_ (
    .A(_0__1_bF$buf0),
    .B(DMEM_DATA_L[10]),
    .Y(_3200_)
);

OAI21X1 _13811_ (
    .A(_0__1_bF$buf10),
    .B(_3199_),
    .C(_3200_),
    .Y(_3201_)
);

NAND2X1 _13812_ (
    .A(_3138__bF$buf3),
    .B(_3201_),
    .Y(_3202_)
);

NAND3X1 _13813_ (
    .A(_3198_),
    .B(_3197_),
    .C(_3202_),
    .Y(_1_[10])
);

NAND3X1 _13814_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [11]),
    .B(_3132__bF$buf0),
    .C(_3134__bF$buf0),
    .Y(_3203_)
);

NAND2X1 _13815_ (
    .A(\datapath.memoryinterface.data_store [11]),
    .B(_3136__bF$buf4),
    .Y(_3204_)
);

INVX1 _13816_ (
    .A(\datapath.memoryinterface.data_store [11]),
    .Y(_3205_)
);

NAND2X1 _13817_ (
    .A(_0__1_bF$buf9),
    .B(DMEM_DATA_L[11]),
    .Y(_3206_)
);

OAI21X1 _13818_ (
    .A(_0__1_bF$buf8),
    .B(_3205_),
    .C(_3206_),
    .Y(_3207_)
);

NAND2X1 _13819_ (
    .A(_3138__bF$buf2),
    .B(_3207_),
    .Y(_3208_)
);

NAND3X1 _13820_ (
    .A(_3204_),
    .B(_3203_),
    .C(_3208_),
    .Y(_1_[11])
);

NAND3X1 _13821_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [12]),
    .B(_3132__bF$buf5),
    .C(_3134__bF$buf5),
    .Y(_3209_)
);

NAND2X1 _13822_ (
    .A(\datapath.memoryinterface.data_store [12]),
    .B(_3136__bF$buf3),
    .Y(_3210_)
);

INVX1 _13823_ (
    .A(\datapath.memoryinterface.data_store [12]),
    .Y(_3211_)
);

NAND2X1 _13824_ (
    .A(_0__1_bF$buf7),
    .B(DMEM_DATA_L[12]),
    .Y(_3212_)
);

OAI21X1 _13825_ (
    .A(_0__1_bF$buf6),
    .B(_3211_),
    .C(_3212_),
    .Y(_3213_)
);

NAND2X1 _13826_ (
    .A(_3138__bF$buf1),
    .B(_3213_),
    .Y(_3214_)
);

NAND3X1 _13827_ (
    .A(_3210_),
    .B(_3209_),
    .C(_3214_),
    .Y(_1_[12])
);

NAND3X1 _13828_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [13]),
    .B(_3132__bF$buf4),
    .C(_3134__bF$buf4),
    .Y(_3215_)
);

NAND2X1 _13829_ (
    .A(\datapath.memoryinterface.data_store [13]),
    .B(_3136__bF$buf2),
    .Y(_3216_)
);

INVX1 _13830_ (
    .A(\datapath.memoryinterface.data_store [13]),
    .Y(_3217_)
);

NAND2X1 _13831_ (
    .A(_0__1_bF$buf5),
    .B(DMEM_DATA_L[13]),
    .Y(_3218_)
);

OAI21X1 _13832_ (
    .A(_0__1_bF$buf4),
    .B(_3217_),
    .C(_3218_),
    .Y(_3219_)
);

NAND2X1 _13833_ (
    .A(_3138__bF$buf0),
    .B(_3219_),
    .Y(_3220_)
);

NAND3X1 _13834_ (
    .A(_3216_),
    .B(_3215_),
    .C(_3220_),
    .Y(_1_[13])
);

NAND3X1 _13835_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [14]),
    .B(_3132__bF$buf3),
    .C(_3134__bF$buf3),
    .Y(_3221_)
);

NAND2X1 _13836_ (
    .A(\datapath.memoryinterface.data_store [14]),
    .B(_3136__bF$buf1),
    .Y(_3222_)
);

INVX1 _13837_ (
    .A(\datapath.memoryinterface.data_store [14]),
    .Y(_3223_)
);

NAND2X1 _13838_ (
    .A(_0__1_bF$buf3),
    .B(DMEM_DATA_L[14]),
    .Y(_3224_)
);

OAI21X1 _13839_ (
    .A(_0__1_bF$buf2),
    .B(_3223_),
    .C(_3224_),
    .Y(_3225_)
);

NAND2X1 _13840_ (
    .A(_3138__bF$buf6),
    .B(_3225_),
    .Y(_3226_)
);

NAND3X1 _13841_ (
    .A(_3222_),
    .B(_3221_),
    .C(_3226_),
    .Y(_1_[14])
);

NAND3X1 _13842_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [15]),
    .B(_3132__bF$buf2),
    .C(_3134__bF$buf2),
    .Y(_3227_)
);

NAND2X1 _13843_ (
    .A(\datapath.memoryinterface.data_store [15]),
    .B(_3136__bF$buf0),
    .Y(_3228_)
);

INVX1 _13844_ (
    .A(\datapath.memoryinterface.data_store [15]),
    .Y(_3229_)
);

NAND2X1 _13845_ (
    .A(_0__1_bF$buf1),
    .B(DMEM_DATA_L[15]),
    .Y(_3230_)
);

OAI21X1 _13846_ (
    .A(_0__1_bF$buf0),
    .B(_3229_),
    .C(_3230_),
    .Y(_3231_)
);

NAND2X1 _13847_ (
    .A(_3138__bF$buf5),
    .B(_3231_),
    .Y(_3232_)
);

NAND3X1 _13848_ (
    .A(_3228_),
    .B(_3227_),
    .C(_3232_),
    .Y(_1_[15])
);

INVX1 _13849_ (
    .A(DMEM_DATA_L[16]),
    .Y(_3233_)
);

NAND2X1 _13850_ (
    .A(\datapath.memoryinterface.data_store [0]),
    .B(_0__1_bF$buf10),
    .Y(_3234_)
);

OAI21X1 _13851_ (
    .A(_0__1_bF$buf9),
    .B(_3233_),
    .C(_3234_),
    .Y(_3235_)
);

NAND2X1 _13852_ (
    .A(_3138__bF$buf4),
    .B(_3235_),
    .Y(_3236_)
);

NAND3X1 _13853_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [16]),
    .B(_3132__bF$buf1),
    .C(_3134__bF$buf1),
    .Y(_3237_)
);

NAND2X1 _13854_ (
    .A(\datapath.memoryinterface.data_store [16]),
    .B(_3136__bF$buf7),
    .Y(_3238_)
);

NAND3X1 _13855_ (
    .A(_3238_),
    .B(_3237_),
    .C(_3236_),
    .Y(_1_[16])
);

INVX1 _13856_ (
    .A(DMEM_DATA_L[17]),
    .Y(_3239_)
);

NAND2X1 _13857_ (
    .A(_0__1_bF$buf8),
    .B(\datapath.memoryinterface.data_store [1]),
    .Y(_3240_)
);

OAI21X1 _13858_ (
    .A(_0__1_bF$buf7),
    .B(_3239_),
    .C(_3240_),
    .Y(_3241_)
);

NAND2X1 _13859_ (
    .A(_3138__bF$buf3),
    .B(_3241_),
    .Y(_3242_)
);

NAND3X1 _13860_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [17]),
    .B(_3132__bF$buf0),
    .C(_3134__bF$buf0),
    .Y(_3243_)
);

NAND2X1 _13861_ (
    .A(\datapath.memoryinterface.data_store [17]),
    .B(_3136__bF$buf6),
    .Y(_3244_)
);

NAND3X1 _13862_ (
    .A(_3244_),
    .B(_3243_),
    .C(_3242_),
    .Y(_1_[17])
);

INVX1 _13863_ (
    .A(DMEM_DATA_L[18]),
    .Y(_3245_)
);

NAND2X1 _13864_ (
    .A(_0__1_bF$buf6),
    .B(\datapath.memoryinterface.data_store [2]),
    .Y(_3246_)
);

OAI21X1 _13865_ (
    .A(_0__1_bF$buf5),
    .B(_3245_),
    .C(_3246_),
    .Y(_3247_)
);

NAND2X1 _13866_ (
    .A(_3138__bF$buf2),
    .B(_3247_),
    .Y(_3248_)
);

NAND3X1 _13867_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [18]),
    .B(_3132__bF$buf5),
    .C(_3134__bF$buf5),
    .Y(_3249_)
);

NAND2X1 _13868_ (
    .A(\datapath.memoryinterface.data_store [18]),
    .B(_3136__bF$buf5),
    .Y(_3250_)
);

NAND3X1 _13869_ (
    .A(_3250_),
    .B(_3249_),
    .C(_3248_),
    .Y(_1_[18])
);

INVX1 _13870_ (
    .A(DMEM_DATA_L[19]),
    .Y(_3251_)
);

NAND2X1 _13871_ (
    .A(_0__1_bF$buf4),
    .B(\datapath.memoryinterface.data_store [3]),
    .Y(_3252_)
);

OAI21X1 _13872_ (
    .A(_0__1_bF$buf3),
    .B(_3251_),
    .C(_3252_),
    .Y(_3253_)
);

NAND2X1 _13873_ (
    .A(_3138__bF$buf1),
    .B(_3253_),
    .Y(_3254_)
);

NAND3X1 _13874_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [19]),
    .B(_3132__bF$buf4),
    .C(_3134__bF$buf4),
    .Y(_3255_)
);

NAND2X1 _13875_ (
    .A(\datapath.memoryinterface.data_store [19]),
    .B(_3136__bF$buf4),
    .Y(_3256_)
);

NAND3X1 _13876_ (
    .A(_3256_),
    .B(_3255_),
    .C(_3254_),
    .Y(_1_[19])
);

INVX1 _13877_ (
    .A(DMEM_DATA_L[20]),
    .Y(_3257_)
);

NAND2X1 _13878_ (
    .A(_0__1_bF$buf2),
    .B(\datapath.memoryinterface.data_store [4]),
    .Y(_3258_)
);

OAI21X1 _13879_ (
    .A(_0__1_bF$buf1),
    .B(_3257_),
    .C(_3258_),
    .Y(_3259_)
);

NAND2X1 _13880_ (
    .A(_3138__bF$buf0),
    .B(_3259_),
    .Y(_3260_)
);

NAND3X1 _13881_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [20]),
    .B(_3132__bF$buf3),
    .C(_3134__bF$buf3),
    .Y(_3261_)
);

NAND2X1 _13882_ (
    .A(\datapath.memoryinterface.data_store [20]),
    .B(_3136__bF$buf3),
    .Y(_3262_)
);

NAND3X1 _13883_ (
    .A(_3262_),
    .B(_3261_),
    .C(_3260_),
    .Y(_1_[20])
);

INVX1 _13884_ (
    .A(DMEM_DATA_L[21]),
    .Y(_3263_)
);

NAND2X1 _13885_ (
    .A(_0__1_bF$buf0),
    .B(\datapath.memoryinterface.data_store [5]),
    .Y(_3264_)
);

OAI21X1 _13886_ (
    .A(_0__1_bF$buf10),
    .B(_3263_),
    .C(_3264_),
    .Y(_3265_)
);

NAND2X1 _13887_ (
    .A(_3138__bF$buf6),
    .B(_3265_),
    .Y(_3266_)
);

NAND3X1 _13888_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [21]),
    .B(_3132__bF$buf2),
    .C(_3134__bF$buf2),
    .Y(_3267_)
);

NAND2X1 _13889_ (
    .A(\datapath.memoryinterface.data_store [21]),
    .B(_3136__bF$buf2),
    .Y(_3268_)
);

NAND3X1 _13890_ (
    .A(_3268_),
    .B(_3267_),
    .C(_3266_),
    .Y(_1_[21])
);

INVX1 _13891_ (
    .A(DMEM_DATA_L[22]),
    .Y(_3269_)
);

NAND2X1 _13892_ (
    .A(_0__1_bF$buf9),
    .B(\datapath.memoryinterface.data_store [6]),
    .Y(_3270_)
);

OAI21X1 _13893_ (
    .A(_0__1_bF$buf8),
    .B(_3269_),
    .C(_3270_),
    .Y(_3271_)
);

NAND2X1 _13894_ (
    .A(_3138__bF$buf5),
    .B(_3271_),
    .Y(_3272_)
);

NAND3X1 _13895_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [22]),
    .B(_3132__bF$buf1),
    .C(_3134__bF$buf1),
    .Y(_3273_)
);

NAND2X1 _13896_ (
    .A(\datapath.memoryinterface.data_store [22]),
    .B(_3136__bF$buf1),
    .Y(_3274_)
);

NAND3X1 _13897_ (
    .A(_3274_),
    .B(_3273_),
    .C(_3272_),
    .Y(_1_[22])
);

INVX1 _13898_ (
    .A(DMEM_DATA_L[23]),
    .Y(_3275_)
);

NAND2X1 _13899_ (
    .A(_0__1_bF$buf7),
    .B(\datapath.memoryinterface.data_store [7]),
    .Y(_3276_)
);

OAI21X1 _13900_ (
    .A(_0__1_bF$buf6),
    .B(_3275_),
    .C(_3276_),
    .Y(_3277_)
);

NAND2X1 _13901_ (
    .A(_3138__bF$buf4),
    .B(_3277_),
    .Y(_3278_)
);

NAND3X1 _13902_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [23]),
    .B(_3132__bF$buf0),
    .C(_3134__bF$buf0),
    .Y(_3279_)
);

NAND2X1 _13903_ (
    .A(\datapath.memoryinterface.data_store [23]),
    .B(_3136__bF$buf0),
    .Y(_3280_)
);

NAND3X1 _13904_ (
    .A(_3280_),
    .B(_3279_),
    .C(_3278_),
    .Y(_1_[23])
);

INVX1 _13905_ (
    .A(DMEM_DATA_L[24]),
    .Y(_3281_)
);

NAND2X1 _13906_ (
    .A(_0__1_bF$buf5),
    .B(\datapath.memoryinterface.data_store [8]),
    .Y(_3282_)
);

OAI21X1 _13907_ (
    .A(_0__1_bF$buf4),
    .B(_3281_),
    .C(_3282_),
    .Y(_3283_)
);

NAND2X1 _13908_ (
    .A(_3138__bF$buf3),
    .B(_3283_),
    .Y(_3284_)
);

NAND3X1 _13909_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [24]),
    .B(_3132__bF$buf5),
    .C(_3134__bF$buf5),
    .Y(_3285_)
);

NAND2X1 _13910_ (
    .A(\datapath.memoryinterface.data_store [24]),
    .B(_3136__bF$buf7),
    .Y(_3286_)
);

NAND3X1 _13911_ (
    .A(_3286_),
    .B(_3285_),
    .C(_3284_),
    .Y(_1_[24])
);

INVX1 _13912_ (
    .A(DMEM_DATA_L[25]),
    .Y(_3287_)
);

NAND2X1 _13913_ (
    .A(_0__1_bF$buf3),
    .B(\datapath.memoryinterface.data_store [9]),
    .Y(_3288_)
);

OAI21X1 _13914_ (
    .A(_0__1_bF$buf2),
    .B(_3287_),
    .C(_3288_),
    .Y(_3289_)
);

NAND2X1 _13915_ (
    .A(_3138__bF$buf2),
    .B(_3289_),
    .Y(_3290_)
);

NAND3X1 _13916_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [25]),
    .B(_3132__bF$buf4),
    .C(_3134__bF$buf4),
    .Y(_3291_)
);

NAND2X1 _13917_ (
    .A(\datapath.memoryinterface.data_store [25]),
    .B(_3136__bF$buf6),
    .Y(_3292_)
);

NAND3X1 _13918_ (
    .A(_3292_),
    .B(_3291_),
    .C(_3290_),
    .Y(_1_[25])
);

INVX1 _13919_ (
    .A(DMEM_DATA_L[26]),
    .Y(_3293_)
);

NAND2X1 _13920_ (
    .A(_0__1_bF$buf1),
    .B(\datapath.memoryinterface.data_store [10]),
    .Y(_3294_)
);

OAI21X1 _13921_ (
    .A(_0__1_bF$buf0),
    .B(_3293_),
    .C(_3294_),
    .Y(_3295_)
);

NAND2X1 _13922_ (
    .A(_3138__bF$buf1),
    .B(_3295_),
    .Y(_3296_)
);

NAND3X1 _13923_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [26]),
    .B(_3132__bF$buf3),
    .C(_3134__bF$buf3),
    .Y(_3297_)
);

NAND2X1 _13924_ (
    .A(\datapath.memoryinterface.data_store [26]),
    .B(_3136__bF$buf5),
    .Y(_3298_)
);

NAND3X1 _13925_ (
    .A(_3298_),
    .B(_3297_),
    .C(_3296_),
    .Y(_1_[26])
);

INVX1 _13926_ (
    .A(DMEM_DATA_L[27]),
    .Y(_3299_)
);

NAND2X1 _13927_ (
    .A(_0__1_bF$buf10),
    .B(\datapath.memoryinterface.data_store [11]),
    .Y(_3300_)
);

OAI21X1 _13928_ (
    .A(_0__1_bF$buf9),
    .B(_3299_),
    .C(_3300_),
    .Y(_3301_)
);

NAND2X1 _13929_ (
    .A(_3138__bF$buf0),
    .B(_3301_),
    .Y(_3302_)
);

NAND3X1 _13930_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [27]),
    .B(_3132__bF$buf2),
    .C(_3134__bF$buf2),
    .Y(_3303_)
);

NAND2X1 _13931_ (
    .A(\datapath.memoryinterface.data_store [27]),
    .B(_3136__bF$buf4),
    .Y(_3304_)
);

NAND3X1 _13932_ (
    .A(_3304_),
    .B(_3303_),
    .C(_3302_),
    .Y(_1_[27])
);

INVX1 _13933_ (
    .A(DMEM_DATA_L[28]),
    .Y(_3305_)
);

NAND2X1 _13934_ (
    .A(_0__1_bF$buf8),
    .B(\datapath.memoryinterface.data_store [12]),
    .Y(_3306_)
);

OAI21X1 _13935_ (
    .A(_0__1_bF$buf7),
    .B(_3305_),
    .C(_3306_),
    .Y(_3307_)
);

NAND2X1 _13936_ (
    .A(_3138__bF$buf6),
    .B(_3307_),
    .Y(_3308_)
);

NAND3X1 _13937_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [28]),
    .B(_3132__bF$buf1),
    .C(_3134__bF$buf1),
    .Y(_3309_)
);

NAND2X1 _13938_ (
    .A(\datapath.memoryinterface.data_store [28]),
    .B(_3136__bF$buf3),
    .Y(_3310_)
);

NAND3X1 _13939_ (
    .A(_3310_),
    .B(_3309_),
    .C(_3308_),
    .Y(_1_[28])
);

INVX1 _13940_ (
    .A(DMEM_DATA_L[29]),
    .Y(_3311_)
);

NAND2X1 _13941_ (
    .A(_0__1_bF$buf6),
    .B(\datapath.memoryinterface.data_store [13]),
    .Y(_3312_)
);

OAI21X1 _13942_ (
    .A(_0__1_bF$buf5),
    .B(_3311_),
    .C(_3312_),
    .Y(_3313_)
);

NAND2X1 _13943_ (
    .A(_3138__bF$buf5),
    .B(_3313_),
    .Y(_3314_)
);

NAND3X1 _13944_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [29]),
    .B(_3132__bF$buf0),
    .C(_3134__bF$buf0),
    .Y(_3315_)
);

NAND2X1 _13945_ (
    .A(\datapath.memoryinterface.data_store [29]),
    .B(_3136__bF$buf2),
    .Y(_3316_)
);

NAND3X1 _13946_ (
    .A(_3316_),
    .B(_3315_),
    .C(_3314_),
    .Y(_1_[29])
);

INVX1 _13947_ (
    .A(DMEM_DATA_L[30]),
    .Y(_3317_)
);

NAND2X1 _13948_ (
    .A(_0__1_bF$buf4),
    .B(\datapath.memoryinterface.data_store [14]),
    .Y(_3318_)
);

OAI21X1 _13949_ (
    .A(_0__1_bF$buf3),
    .B(_3317_),
    .C(_3318_),
    .Y(_3319_)
);

NAND2X1 _13950_ (
    .A(_3138__bF$buf4),
    .B(_3319_),
    .Y(_3320_)
);

NAND3X1 _13951_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [30]),
    .B(_3132__bF$buf5),
    .C(_3134__bF$buf5),
    .Y(_3321_)
);

NAND2X1 _13952_ (
    .A(\datapath.memoryinterface.data_store [30]),
    .B(_3136__bF$buf1),
    .Y(_3322_)
);

NAND3X1 _13953_ (
    .A(_3322_),
    .B(_3321_),
    .C(_3320_),
    .Y(_1_[30])
);

INVX1 _13954_ (
    .A(DMEM_DATA_L[31]),
    .Y(_3323_)
);

NAND2X1 _13955_ (
    .A(_0__1_bF$buf2),
    .B(\datapath.memoryinterface.data_store [15]),
    .Y(_3324_)
);

OAI21X1 _13956_ (
    .A(_0__1_bF$buf1),
    .B(_3323_),
    .C(_3324_),
    .Y(_3325_)
);

NAND2X1 _13957_ (
    .A(_3138__bF$buf3),
    .B(_3325_),
    .Y(_3326_)
);

NAND3X1 _13958_ (
    .A(\datapath.memoryinterface.byte_size_store.storebyte [31]),
    .B(_3132__bF$buf4),
    .C(_3134__bF$buf4),
    .Y(_3327_)
);

NAND2X1 _13959_ (
    .A(\datapath.memoryinterface.data_store [31]),
    .B(_3136__bF$buf0),
    .Y(_3328_)
);

NAND3X1 _13960_ (
    .A(_3328_),
    .B(_3327_),
    .C(_3326_),
    .Y(_1_[31])
);

NOR2X1 _13961_ (
    .A(_0__1_bF$buf0),
    .B(_0__0_bF$buf3),
    .Y(_3329_)
);

INVX4 _13962_ (
    .A(_3329_),
    .Y(_3330_)
);

OAI21X1 _13963_ (
    .A(_0__1_bF$buf10),
    .B(_0__0_bF$buf2),
    .C(DMEM_DATA_L[0]),
    .Y(_3331_)
);

OAI21X1 _13964_ (
    .A(_3139_),
    .B(_3330_),
    .C(_3331_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [0])
);

OAI21X1 _13965_ (
    .A(_0__1_bF$buf9),
    .B(_0__0_bF$buf1),
    .C(DMEM_DATA_L[1]),
    .Y(_3332_)
);

OAI21X1 _13966_ (
    .A(_3145_),
    .B(_3330_),
    .C(_3332_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [1])
);

OAI21X1 _13967_ (
    .A(_0__1_bF$buf8),
    .B(_0__0_bF$buf0),
    .C(DMEM_DATA_L[2]),
    .Y(_3333_)
);

OAI21X1 _13968_ (
    .A(_3151_),
    .B(_3330_),
    .C(_3333_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [2])
);

OAI21X1 _13969_ (
    .A(_0__1_bF$buf7),
    .B(_0__0_bF$buf4),
    .C(DMEM_DATA_L[3]),
    .Y(_3334_)
);

OAI21X1 _13970_ (
    .A(_3157_),
    .B(_3330_),
    .C(_3334_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [3])
);

OAI21X1 _13971_ (
    .A(_0__1_bF$buf6),
    .B(_0__0_bF$buf3),
    .C(DMEM_DATA_L[4]),
    .Y(_3335_)
);

OAI21X1 _13972_ (
    .A(_3163_),
    .B(_3330_),
    .C(_3335_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [4])
);

OAI21X1 _13973_ (
    .A(_0__1_bF$buf5),
    .B(_0__0_bF$buf2),
    .C(DMEM_DATA_L[5]),
    .Y(_3336_)
);

OAI21X1 _13974_ (
    .A(_3169_),
    .B(_3330_),
    .C(_3336_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [5])
);

OAI21X1 _13975_ (
    .A(_0__1_bF$buf4),
    .B(_0__0_bF$buf1),
    .C(DMEM_DATA_L[6]),
    .Y(_3337_)
);

OAI21X1 _13976_ (
    .A(_3175_),
    .B(_3330_),
    .C(_3337_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [6])
);

OAI21X1 _13977_ (
    .A(_0__1_bF$buf3),
    .B(_0__0_bF$buf0),
    .C(DMEM_DATA_L[7]),
    .Y(_3338_)
);

OAI21X1 _13978_ (
    .A(_3181_),
    .B(_3330_),
    .C(_3338_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [7])
);

INVX1 _13979_ (
    .A(DMEM_DATA_L[8]),
    .Y(_3339_)
);

INVX1 _13980_ (
    .A(_0__0_bF$buf4),
    .Y(_3340_)
);

NOR2X1 _13981_ (
    .A(_0__1_bF$buf2),
    .B(_3340_),
    .Y(_3341_)
);

MUX2X1 _13982_ (
    .A(_3139_),
    .B(_3339_),
    .S(_3341_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [8])
);

INVX1 _13983_ (
    .A(DMEM_DATA_L[9]),
    .Y(_3342_)
);

MUX2X1 _13984_ (
    .A(_3145_),
    .B(_3342_),
    .S(_3341_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [9])
);

INVX1 _13985_ (
    .A(DMEM_DATA_L[10]),
    .Y(_3343_)
);

MUX2X1 _13986_ (
    .A(_3151_),
    .B(_3343_),
    .S(_3341_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [10])
);

INVX1 _13987_ (
    .A(DMEM_DATA_L[11]),
    .Y(_3344_)
);

MUX2X1 _13988_ (
    .A(_3157_),
    .B(_3344_),
    .S(_3341_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [11])
);

INVX1 _13989_ (
    .A(DMEM_DATA_L[12]),
    .Y(_3345_)
);

MUX2X1 _13990_ (
    .A(_3163_),
    .B(_3345_),
    .S(_3341_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [12])
);

INVX1 _13991_ (
    .A(DMEM_DATA_L[13]),
    .Y(_3346_)
);

MUX2X1 _13992_ (
    .A(_3169_),
    .B(_3346_),
    .S(_3341_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [13])
);

INVX1 _13993_ (
    .A(DMEM_DATA_L[14]),
    .Y(_3347_)
);

MUX2X1 _13994_ (
    .A(_3175_),
    .B(_3347_),
    .S(_3341_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [14])
);

INVX1 _13995_ (
    .A(DMEM_DATA_L[15]),
    .Y(_3348_)
);

MUX2X1 _13996_ (
    .A(_3181_),
    .B(_3348_),
    .S(_3341_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [15])
);

INVX1 _13997_ (
    .A(_0__1_bF$buf1),
    .Y(_3349_)
);

NOR2X1 _13998_ (
    .A(_0__0_bF$buf3),
    .B(_3349_),
    .Y(_3350_)
);

OAI22X1 _13999_ (
    .A(_0__0_bF$buf2),
    .B(_3234_),
    .C(_3233_),
    .D(_3350_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [16])
);

OAI22X1 _14000_ (
    .A(_0__0_bF$buf1),
    .B(_3240_),
    .C(_3239_),
    .D(_3350_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [17])
);

OAI22X1 _14001_ (
    .A(_0__0_bF$buf0),
    .B(_3246_),
    .C(_3245_),
    .D(_3350_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [18])
);

OAI22X1 _14002_ (
    .A(_0__0_bF$buf4),
    .B(_3252_),
    .C(_3251_),
    .D(_3350_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [19])
);

OAI22X1 _14003_ (
    .A(_0__0_bF$buf3),
    .B(_3258_),
    .C(_3257_),
    .D(_3350_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [20])
);

OAI22X1 _14004_ (
    .A(_0__0_bF$buf2),
    .B(_3264_),
    .C(_3263_),
    .D(_3350_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [21])
);

OAI22X1 _14005_ (
    .A(_0__0_bF$buf1),
    .B(_3270_),
    .C(_3269_),
    .D(_3350_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [22])
);

OAI22X1 _14006_ (
    .A(_0__0_bF$buf0),
    .B(_3276_),
    .C(_3275_),
    .D(_3350_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [23])
);

NOR2X1 _14007_ (
    .A(_3349_),
    .B(_3340_),
    .Y(_3351_)
);

NAND2X1 _14008_ (
    .A(\datapath.memoryinterface.data_store [0]),
    .B(_3351_),
    .Y(_3352_)
);

OAI21X1 _14009_ (
    .A(_3281_),
    .B(_3351_),
    .C(_3352_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [24])
);

NAND2X1 _14010_ (
    .A(\datapath.memoryinterface.data_store [1]),
    .B(_3351_),
    .Y(_3353_)
);

OAI21X1 _14011_ (
    .A(_3287_),
    .B(_3351_),
    .C(_3353_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [25])
);

NAND2X1 _14012_ (
    .A(\datapath.memoryinterface.data_store [2]),
    .B(_3351_),
    .Y(_3354_)
);

OAI21X1 _14013_ (
    .A(_3293_),
    .B(_3351_),
    .C(_3354_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [26])
);

NAND2X1 _14014_ (
    .A(\datapath.memoryinterface.data_store [3]),
    .B(_3351_),
    .Y(_3355_)
);

OAI21X1 _14015_ (
    .A(_3299_),
    .B(_3351_),
    .C(_3355_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [27])
);

NAND2X1 _14016_ (
    .A(\datapath.memoryinterface.data_store [4]),
    .B(_3351_),
    .Y(_3356_)
);

OAI21X1 _14017_ (
    .A(_3305_),
    .B(_3351_),
    .C(_3356_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [28])
);

NAND2X1 _14018_ (
    .A(\datapath.memoryinterface.data_store [5]),
    .B(_3351_),
    .Y(_3357_)
);

OAI21X1 _14019_ (
    .A(_3311_),
    .B(_3351_),
    .C(_3357_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [29])
);

NAND2X1 _14020_ (
    .A(\datapath.memoryinterface.data_store [6]),
    .B(_3351_),
    .Y(_3358_)
);

OAI21X1 _14021_ (
    .A(_3317_),
    .B(_3351_),
    .C(_3358_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [30])
);

NAND2X1 _14022_ (
    .A(\datapath.memoryinterface.data_store [7]),
    .B(_3351_),
    .Y(_3359_)
);

OAI21X1 _14023_ (
    .A(_3323_),
    .B(_3351_),
    .C(_3359_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [31])
);

NAND3X1 _14024_ (
    .A(\datapath.memoryinterface.byte_size_load.byteval [0]),
    .B(_3132__bF$buf3),
    .C(_3134__bF$buf3),
    .Y(_3360_)
);

NAND2X1 _14025_ (
    .A(DMEM_DATA_L[0]),
    .B(_3136__bF$buf7),
    .Y(_3361_)
);

INVX1 _14026_ (
    .A(DMEM_DATA_L[0]),
    .Y(_3362_)
);

NAND2X1 _14027_ (
    .A(_0__1_bF$buf0),
    .B(DMEM_DATA_L[16]),
    .Y(_3363_)
);

OAI21X1 _14028_ (
    .A(_0__1_bF$buf10),
    .B(_3362_),
    .C(_3363_),
    .Y(_3364_)
);

NAND2X1 _14029_ (
    .A(_3138__bF$buf2),
    .B(_3364_),
    .Y(_3365_)
);

NAND3X1 _14030_ (
    .A(_3361_),
    .B(_3360_),
    .C(_3365_),
    .Y(\datapath.memdataload [0])
);

NAND3X1 _14031_ (
    .A(\datapath.memoryinterface.byte_size_load.byteval [1]),
    .B(_3132__bF$buf2),
    .C(_3134__bF$buf2),
    .Y(_3366_)
);

NAND2X1 _14032_ (
    .A(DMEM_DATA_L[1]),
    .B(_3136__bF$buf6),
    .Y(_3367_)
);

INVX1 _14033_ (
    .A(DMEM_DATA_L[1]),
    .Y(_3368_)
);

NAND2X1 _14034_ (
    .A(_0__1_bF$buf9),
    .B(DMEM_DATA_L[17]),
    .Y(_3369_)
);

OAI21X1 _14035_ (
    .A(_0__1_bF$buf8),
    .B(_3368_),
    .C(_3369_),
    .Y(_3370_)
);

NAND2X1 _14036_ (
    .A(_3138__bF$buf1),
    .B(_3370_),
    .Y(_3371_)
);

NAND3X1 _14037_ (
    .A(_3367_),
    .B(_3366_),
    .C(_3371_),
    .Y(\datapath.memdataload [1])
);

NAND3X1 _14038_ (
    .A(\datapath.memoryinterface.byte_size_load.byteval [2]),
    .B(_3132__bF$buf1),
    .C(_3134__bF$buf1),
    .Y(_3372_)
);

NAND2X1 _14039_ (
    .A(DMEM_DATA_L[2]),
    .B(_3136__bF$buf5),
    .Y(_3373_)
);

INVX1 _14040_ (
    .A(DMEM_DATA_L[2]),
    .Y(_3374_)
);

NAND2X1 _14041_ (
    .A(_0__1_bF$buf7),
    .B(DMEM_DATA_L[18]),
    .Y(_3375_)
);

OAI21X1 _14042_ (
    .A(_0__1_bF$buf6),
    .B(_3374_),
    .C(_3375_),
    .Y(_3376_)
);

NAND2X1 _14043_ (
    .A(_3138__bF$buf0),
    .B(_3376_),
    .Y(_3377_)
);

NAND3X1 _14044_ (
    .A(_3373_),
    .B(_3372_),
    .C(_3377_),
    .Y(\datapath.memdataload [2])
);

NAND3X1 _14045_ (
    .A(\datapath.memoryinterface.byte_size_load.byteval [3]),
    .B(_3132__bF$buf0),
    .C(_3134__bF$buf0),
    .Y(_3378_)
);

NAND2X1 _14046_ (
    .A(DMEM_DATA_L[3]),
    .B(_3136__bF$buf4),
    .Y(_3379_)
);

INVX1 _14047_ (
    .A(DMEM_DATA_L[3]),
    .Y(_3380_)
);

NAND2X1 _14048_ (
    .A(_0__1_bF$buf5),
    .B(DMEM_DATA_L[19]),
    .Y(_3381_)
);

OAI21X1 _14049_ (
    .A(_0__1_bF$buf4),
    .B(_3380_),
    .C(_3381_),
    .Y(_3382_)
);

NAND2X1 _14050_ (
    .A(_3138__bF$buf6),
    .B(_3382_),
    .Y(_3383_)
);

NAND3X1 _14051_ (
    .A(_3379_),
    .B(_3378_),
    .C(_3383_),
    .Y(\datapath.memdataload [3])
);

NAND3X1 _14052_ (
    .A(\datapath.memoryinterface.byte_size_load.byteval [4]),
    .B(_3132__bF$buf5),
    .C(_3134__bF$buf5),
    .Y(_3384_)
);

NAND2X1 _14053_ (
    .A(DMEM_DATA_L[4]),
    .B(_3136__bF$buf3),
    .Y(_3385_)
);

INVX1 _14054_ (
    .A(DMEM_DATA_L[4]),
    .Y(_3386_)
);

NAND2X1 _14055_ (
    .A(_0__1_bF$buf3),
    .B(DMEM_DATA_L[20]),
    .Y(_3387_)
);

OAI21X1 _14056_ (
    .A(_0__1_bF$buf2),
    .B(_3386_),
    .C(_3387_),
    .Y(_3388_)
);

NAND2X1 _14057_ (
    .A(_3138__bF$buf5),
    .B(_3388_),
    .Y(_3389_)
);

NAND3X1 _14058_ (
    .A(_3385_),
    .B(_3384_),
    .C(_3389_),
    .Y(\datapath.memdataload [4])
);

NAND3X1 _14059_ (
    .A(\datapath.memoryinterface.byte_size_load.byteval [5]),
    .B(_3132__bF$buf4),
    .C(_3134__bF$buf4),
    .Y(_3390_)
);

NAND2X1 _14060_ (
    .A(DMEM_DATA_L[5]),
    .B(_3136__bF$buf2),
    .Y(_3391_)
);

INVX1 _14061_ (
    .A(DMEM_DATA_L[5]),
    .Y(_3392_)
);

NAND2X1 _14062_ (
    .A(_0__1_bF$buf1),
    .B(DMEM_DATA_L[21]),
    .Y(_3393_)
);

OAI21X1 _14063_ (
    .A(_0__1_bF$buf0),
    .B(_3392_),
    .C(_3393_),
    .Y(_3394_)
);

NAND2X1 _14064_ (
    .A(_3138__bF$buf4),
    .B(_3394_),
    .Y(_3395_)
);

NAND3X1 _14065_ (
    .A(_3391_),
    .B(_3390_),
    .C(_3395_),
    .Y(\datapath.memdataload [5])
);

NAND3X1 _14066_ (
    .A(\datapath.memoryinterface.byte_size_load.byteval [6]),
    .B(_3132__bF$buf3),
    .C(_3134__bF$buf3),
    .Y(_3396_)
);

NAND2X1 _14067_ (
    .A(DMEM_DATA_L[6]),
    .B(_3136__bF$buf1),
    .Y(_3397_)
);

INVX1 _14068_ (
    .A(DMEM_DATA_L[6]),
    .Y(_3398_)
);

NAND2X1 _14069_ (
    .A(_0__1_bF$buf10),
    .B(DMEM_DATA_L[22]),
    .Y(_3399_)
);

OAI21X1 _14070_ (
    .A(_0__1_bF$buf9),
    .B(_3398_),
    .C(_3399_),
    .Y(_3400_)
);

NAND2X1 _14071_ (
    .A(_3138__bF$buf3),
    .B(_3400_),
    .Y(_3401_)
);

NAND3X1 _14072_ (
    .A(_3397_),
    .B(_3396_),
    .C(_3401_),
    .Y(\datapath.memdataload [6])
);

NAND3X1 _14073_ (
    .A(\datapath.memoryinterface.byte_size_load.byteval [7]),
    .B(_3132__bF$buf2),
    .C(_3134__bF$buf2),
    .Y(_3402_)
);

NAND2X1 _14074_ (
    .A(DMEM_DATA_L[7]),
    .B(_3136__bF$buf0),
    .Y(_3403_)
);

INVX1 _14075_ (
    .A(DMEM_DATA_L[7]),
    .Y(_3404_)
);

NAND2X1 _14076_ (
    .A(_0__1_bF$buf8),
    .B(DMEM_DATA_L[23]),
    .Y(_3405_)
);

OAI21X1 _14077_ (
    .A(_0__1_bF$buf7),
    .B(_3404_),
    .C(_3405_),
    .Y(_3406_)
);

NAND2X1 _14078_ (
    .A(_3138__bF$buf2),
    .B(_3406_),
    .Y(_3407_)
);

NAND3X1 _14079_ (
    .A(_3403_),
    .B(_3402_),
    .C(_3407_),
    .Y(\datapath.memdataload [7])
);

INVX1 _14080_ (
    .A(\datapath.memoryinterface.byte_size_load.byteval [7]),
    .Y(_3408_)
);

NOR2X1 _14081_ (
    .A(\datapath.meminstr [14]),
    .B(_3408_),
    .Y(_3409_)
);

NAND3X1 _14082_ (
    .A(_3132__bF$buf1),
    .B(_3134__bF$buf1),
    .C(_3409_),
    .Y(_3410_)
);

NAND2X1 _14083_ (
    .A(DMEM_DATA_L[8]),
    .B(_3136__bF$buf7),
    .Y(_3411_)
);

NAND2X1 _14084_ (
    .A(_0__1_bF$buf6),
    .B(DMEM_DATA_L[24]),
    .Y(_3412_)
);

OAI21X1 _14085_ (
    .A(_0__1_bF$buf5),
    .B(_3339_),
    .C(_3412_),
    .Y(_3413_)
);

NAND2X1 _14086_ (
    .A(_3138__bF$buf1),
    .B(_3413_),
    .Y(_3414_)
);

NAND3X1 _14087_ (
    .A(_3411_),
    .B(_3414_),
    .C(_3410__bF$buf3),
    .Y(\datapath.memdataload [8])
);

NAND2X1 _14088_ (
    .A(DMEM_DATA_L[9]),
    .B(_3136__bF$buf6),
    .Y(_3415_)
);

NAND2X1 _14089_ (
    .A(_0__1_bF$buf4),
    .B(DMEM_DATA_L[25]),
    .Y(_3416_)
);

OAI21X1 _14090_ (
    .A(_0__1_bF$buf3),
    .B(_3342_),
    .C(_3416_),
    .Y(_3417_)
);

NAND2X1 _14091_ (
    .A(_3138__bF$buf0),
    .B(_3417_),
    .Y(_3418_)
);

NAND3X1 _14092_ (
    .A(_3415_),
    .B(_3418_),
    .C(_3410__bF$buf2),
    .Y(\datapath.memdataload [9])
);

NAND2X1 _14093_ (
    .A(DMEM_DATA_L[10]),
    .B(_3136__bF$buf5),
    .Y(_3419_)
);

NAND2X1 _14094_ (
    .A(_0__1_bF$buf2),
    .B(DMEM_DATA_L[26]),
    .Y(_3420_)
);

OAI21X1 _14095_ (
    .A(_0__1_bF$buf1),
    .B(_3343_),
    .C(_3420_),
    .Y(_3421_)
);

NAND2X1 _14096_ (
    .A(_3138__bF$buf6),
    .B(_3421_),
    .Y(_3422_)
);

NAND3X1 _14097_ (
    .A(_3419_),
    .B(_3422_),
    .C(_3410__bF$buf1),
    .Y(\datapath.memdataload [10])
);

NAND2X1 _14098_ (
    .A(DMEM_DATA_L[11]),
    .B(_3136__bF$buf4),
    .Y(_3423_)
);

NAND2X1 _14099_ (
    .A(_0__1_bF$buf0),
    .B(DMEM_DATA_L[27]),
    .Y(_3424_)
);

OAI21X1 _14100_ (
    .A(_0__1_bF$buf10),
    .B(_3344_),
    .C(_3424_),
    .Y(_3425_)
);

NAND2X1 _14101_ (
    .A(_3138__bF$buf5),
    .B(_3425_),
    .Y(_3426_)
);

NAND3X1 _14102_ (
    .A(_3423_),
    .B(_3426_),
    .C(_3410__bF$buf0),
    .Y(\datapath.memdataload [11])
);

NAND2X1 _14103_ (
    .A(DMEM_DATA_L[12]),
    .B(_3136__bF$buf3),
    .Y(_3427_)
);

NAND2X1 _14104_ (
    .A(_0__1_bF$buf9),
    .B(DMEM_DATA_L[28]),
    .Y(_3428_)
);

OAI21X1 _14105_ (
    .A(_0__1_bF$buf8),
    .B(_3345_),
    .C(_3428_),
    .Y(_3429_)
);

NAND2X1 _14106_ (
    .A(_3138__bF$buf4),
    .B(_3429_),
    .Y(_3430_)
);

NAND3X1 _14107_ (
    .A(_3427_),
    .B(_3430_),
    .C(_3410__bF$buf3),
    .Y(\datapath.memdataload [12])
);

NAND2X1 _14108_ (
    .A(DMEM_DATA_L[13]),
    .B(_3136__bF$buf2),
    .Y(_3431_)
);

NAND2X1 _14109_ (
    .A(_0__1_bF$buf7),
    .B(DMEM_DATA_L[29]),
    .Y(_3432_)
);

OAI21X1 _14110_ (
    .A(_0__1_bF$buf6),
    .B(_3346_),
    .C(_3432_),
    .Y(_3433_)
);

NAND2X1 _14111_ (
    .A(_3138__bF$buf3),
    .B(_3433_),
    .Y(_3434_)
);

NAND3X1 _14112_ (
    .A(_3431_),
    .B(_3434_),
    .C(_3410__bF$buf2),
    .Y(\datapath.memdataload [13])
);

NAND2X1 _14113_ (
    .A(DMEM_DATA_L[14]),
    .B(_3136__bF$buf1),
    .Y(_3435_)
);

NAND2X1 _14114_ (
    .A(_0__1_bF$buf5),
    .B(DMEM_DATA_L[30]),
    .Y(_3436_)
);

OAI21X1 _14115_ (
    .A(_0__1_bF$buf4),
    .B(_3347_),
    .C(_3436_),
    .Y(_3437_)
);

NAND2X1 _14116_ (
    .A(_3138__bF$buf2),
    .B(_3437_),
    .Y(_3438_)
);

NAND3X1 _14117_ (
    .A(_3435_),
    .B(_3438_),
    .C(_3410__bF$buf1),
    .Y(\datapath.memdataload [14])
);

NAND2X1 _14118_ (
    .A(_0__1_bF$buf3),
    .B(DMEM_DATA_L[31]),
    .Y(_3439_)
);

OAI21X1 _14119_ (
    .A(_0__1_bF$buf2),
    .B(_3348_),
    .C(_3439_),
    .Y(_3440_)
);

NAND2X1 _14120_ (
    .A(_3138__bF$buf1),
    .B(_3440_),
    .Y(_3441_)
);

NAND2X1 _14121_ (
    .A(DMEM_DATA_L[15]),
    .B(_3136__bF$buf0),
    .Y(_3442_)
);

NAND3X1 _14122_ (
    .A(_3442_),
    .B(_3441_),
    .C(_3410__bF$buf0),
    .Y(\datapath.memdataload [15])
);

NAND2X1 _14123_ (
    .A(DMEM_DATA_L[16]),
    .B(_3136__bF$buf7),
    .Y(_3443_)
);

INVX1 _14124_ (
    .A(\datapath.meminstr [14]),
    .Y(_3444_)
);

NAND3X1 _14125_ (
    .A(_3444_),
    .B(_3138__bF$buf0),
    .C(_3440_),
    .Y(_3445_)
);

NAND3X1 _14126_ (
    .A(_3443_),
    .B(_3410__bF$buf3),
    .C(_3445_),
    .Y(\datapath.memdataload [16])
);

NAND2X1 _14127_ (
    .A(DMEM_DATA_L[17]),
    .B(_3136__bF$buf6),
    .Y(_3446_)
);

NAND3X1 _14128_ (
    .A(_3446_),
    .B(_3410__bF$buf2),
    .C(_3445_),
    .Y(\datapath.memdataload [17])
);

NAND2X1 _14129_ (
    .A(DMEM_DATA_L[18]),
    .B(_3136__bF$buf5),
    .Y(_3447_)
);

NAND3X1 _14130_ (
    .A(_3447_),
    .B(_3410__bF$buf1),
    .C(_3445_),
    .Y(\datapath.memdataload [18])
);

NAND2X1 _14131_ (
    .A(DMEM_DATA_L[19]),
    .B(_3136__bF$buf4),
    .Y(_3448_)
);

NAND3X1 _14132_ (
    .A(_3448_),
    .B(_3410__bF$buf0),
    .C(_3445_),
    .Y(\datapath.memdataload [19])
);

NAND2X1 _14133_ (
    .A(DMEM_DATA_L[20]),
    .B(_3136__bF$buf3),
    .Y(_3449_)
);

NAND3X1 _14134_ (
    .A(_3449_),
    .B(_3410__bF$buf3),
    .C(_3445_),
    .Y(\datapath.memdataload [20])
);

NAND2X1 _14135_ (
    .A(DMEM_DATA_L[21]),
    .B(_3136__bF$buf2),
    .Y(_3450_)
);

NAND3X1 _14136_ (
    .A(_3450_),
    .B(_3410__bF$buf2),
    .C(_3445_),
    .Y(\datapath.memdataload [21])
);

NAND2X1 _14137_ (
    .A(DMEM_DATA_L[22]),
    .B(_3136__bF$buf1),
    .Y(_3451_)
);

NAND3X1 _14138_ (
    .A(_3451_),
    .B(_3410__bF$buf1),
    .C(_3445_),
    .Y(\datapath.memdataload [22])
);

NAND2X1 _14139_ (
    .A(DMEM_DATA_L[23]),
    .B(_3136__bF$buf0),
    .Y(_3452_)
);

NAND3X1 _14140_ (
    .A(_3452_),
    .B(_3410__bF$buf0),
    .C(_3445_),
    .Y(\datapath.memdataload [23])
);

NAND2X1 _14141_ (
    .A(DMEM_DATA_L[24]),
    .B(_3136__bF$buf7),
    .Y(_3453_)
);

NAND3X1 _14142_ (
    .A(_3453_),
    .B(_3410__bF$buf3),
    .C(_3445_),
    .Y(\datapath.memdataload [24])
);

NAND2X1 _14143_ (
    .A(DMEM_DATA_L[25]),
    .B(_3136__bF$buf6),
    .Y(_3454_)
);

NAND3X1 _14144_ (
    .A(_3454_),
    .B(_3410__bF$buf2),
    .C(_3445_),
    .Y(\datapath.memdataload [25])
);

NAND2X1 _14145_ (
    .A(DMEM_DATA_L[26]),
    .B(_3136__bF$buf5),
    .Y(_3455_)
);

NAND3X1 _14146_ (
    .A(_3455_),
    .B(_3410__bF$buf1),
    .C(_3445_),
    .Y(\datapath.memdataload [26])
);

NAND2X1 _14147_ (
    .A(DMEM_DATA_L[27]),
    .B(_3136__bF$buf4),
    .Y(_3456_)
);

NAND3X1 _14148_ (
    .A(_3456_),
    .B(_3410__bF$buf0),
    .C(_3445_),
    .Y(\datapath.memdataload [27])
);

NAND2X1 _14149_ (
    .A(DMEM_DATA_L[28]),
    .B(_3136__bF$buf3),
    .Y(_3457_)
);

NAND3X1 _14150_ (
    .A(_3457_),
    .B(_3410__bF$buf3),
    .C(_3445_),
    .Y(\datapath.memdataload [28])
);

NAND2X1 _14151_ (
    .A(DMEM_DATA_L[29]),
    .B(_3136__bF$buf2),
    .Y(_3458_)
);

NAND3X1 _14152_ (
    .A(_3458_),
    .B(_3410__bF$buf2),
    .C(_3445_),
    .Y(\datapath.memdataload [29])
);

NAND2X1 _14153_ (
    .A(DMEM_DATA_L[30]),
    .B(_3136__bF$buf1),
    .Y(_3459_)
);

NAND3X1 _14154_ (
    .A(_3459_),
    .B(_3410__bF$buf1),
    .C(_3445_),
    .Y(\datapath.memdataload [30])
);

NAND2X1 _14155_ (
    .A(DMEM_DATA_L[31]),
    .B(_3136__bF$buf0),
    .Y(_3460_)
);

NAND3X1 _14156_ (
    .A(_3460_),
    .B(_3410__bF$buf0),
    .C(_3445_),
    .Y(\datapath.memdataload [31])
);

NAND3X1 _14157_ (
    .A(_0__1_bF$buf1),
    .B(DMEM_DATA_L[24]),
    .C(_0__0_bF$buf4),
    .Y(_3461_)
);

INVX1 _14158_ (
    .A(_3461_),
    .Y(_3462_)
);

AOI21X1 _14159_ (
    .A(_3350_),
    .B(DMEM_DATA_L[16]),
    .C(_3462_),
    .Y(_3463_)
);

AOI22X1 _14160_ (
    .A(DMEM_DATA_L[0]),
    .B(_3329_),
    .C(DMEM_DATA_L[8]),
    .D(_3341_),
    .Y(_3464_)
);

NAND2X1 _14161_ (
    .A(_3464_),
    .B(_3463_),
    .Y(\datapath.memoryinterface.byte_size_load.byteval [0])
);

NAND3X1 _14162_ (
    .A(_0__1_bF$buf0),
    .B(DMEM_DATA_L[25]),
    .C(_0__0_bF$buf3),
    .Y(_3465_)
);

INVX1 _14163_ (
    .A(_3465_),
    .Y(_3466_)
);

AOI21X1 _14164_ (
    .A(_3350_),
    .B(DMEM_DATA_L[17]),
    .C(_3466_),
    .Y(_3467_)
);

AOI22X1 _14165_ (
    .A(DMEM_DATA_L[1]),
    .B(_3329_),
    .C(DMEM_DATA_L[9]),
    .D(_3341_),
    .Y(_3468_)
);

NAND2X1 _14166_ (
    .A(_3468_),
    .B(_3467_),
    .Y(\datapath.memoryinterface.byte_size_load.byteval [1])
);

NAND3X1 _14167_ (
    .A(_0__1_bF$buf10),
    .B(DMEM_DATA_L[26]),
    .C(_0__0_bF$buf2),
    .Y(_3469_)
);

INVX1 _14168_ (
    .A(_3469_),
    .Y(_3470_)
);

AOI21X1 _14169_ (
    .A(_3350_),
    .B(DMEM_DATA_L[18]),
    .C(_3470_),
    .Y(_3471_)
);

AOI22X1 _14170_ (
    .A(DMEM_DATA_L[2]),
    .B(_3329_),
    .C(DMEM_DATA_L[10]),
    .D(_3341_),
    .Y(_3472_)
);

NAND2X1 _14171_ (
    .A(_3472_),
    .B(_3471_),
    .Y(\datapath.memoryinterface.byte_size_load.byteval [2])
);

NAND3X1 _14172_ (
    .A(_0__1_bF$buf9),
    .B(DMEM_DATA_L[27]),
    .C(_0__0_bF$buf1),
    .Y(_3473_)
);

INVX1 _14173_ (
    .A(_3473_),
    .Y(_3474_)
);

AOI21X1 _14174_ (
    .A(_3350_),
    .B(DMEM_DATA_L[19]),
    .C(_3474_),
    .Y(_3475_)
);

AOI22X1 _14175_ (
    .A(DMEM_DATA_L[3]),
    .B(_3329_),
    .C(DMEM_DATA_L[11]),
    .D(_3341_),
    .Y(_3476_)
);

NAND2X1 _14176_ (
    .A(_3476_),
    .B(_3475_),
    .Y(\datapath.memoryinterface.byte_size_load.byteval [3])
);

NAND3X1 _14177_ (
    .A(_0__1_bF$buf8),
    .B(DMEM_DATA_L[28]),
    .C(_0__0_bF$buf0),
    .Y(_3477_)
);

INVX1 _14178_ (
    .A(_3477_),
    .Y(_3478_)
);

AOI21X1 _14179_ (
    .A(_3350_),
    .B(DMEM_DATA_L[20]),
    .C(_3478_),
    .Y(_3479_)
);

AOI22X1 _14180_ (
    .A(DMEM_DATA_L[4]),
    .B(_3329_),
    .C(DMEM_DATA_L[12]),
    .D(_3341_),
    .Y(_3480_)
);

NAND2X1 _14181_ (
    .A(_3480_),
    .B(_3479_),
    .Y(\datapath.memoryinterface.byte_size_load.byteval [4])
);

NAND3X1 _14182_ (
    .A(_0__1_bF$buf7),
    .B(DMEM_DATA_L[29]),
    .C(_0__0_bF$buf4),
    .Y(_3481_)
);

INVX1 _14183_ (
    .A(_3481_),
    .Y(_3482_)
);

AOI21X1 _14184_ (
    .A(_3350_),
    .B(DMEM_DATA_L[21]),
    .C(_3482_),
    .Y(_3483_)
);

AOI22X1 _14185_ (
    .A(DMEM_DATA_L[5]),
    .B(_3329_),
    .C(DMEM_DATA_L[13]),
    .D(_3341_),
    .Y(_3484_)
);

NAND2X1 _14186_ (
    .A(_3484_),
    .B(_3483_),
    .Y(\datapath.memoryinterface.byte_size_load.byteval [5])
);

NAND3X1 _14187_ (
    .A(_0__1_bF$buf6),
    .B(DMEM_DATA_L[30]),
    .C(_0__0_bF$buf3),
    .Y(_3485_)
);

INVX1 _14188_ (
    .A(_3485_),
    .Y(_3486_)
);

AOI21X1 _14189_ (
    .A(_3350_),
    .B(DMEM_DATA_L[22]),
    .C(_3486_),
    .Y(_3487_)
);

AOI22X1 _14190_ (
    .A(DMEM_DATA_L[6]),
    .B(_3329_),
    .C(DMEM_DATA_L[14]),
    .D(_3341_),
    .Y(_3488_)
);

NAND2X1 _14191_ (
    .A(_3488_),
    .B(_3487_),
    .Y(\datapath.memoryinterface.byte_size_load.byteval [6])
);

AOI22X1 _14192_ (
    .A(DMEM_DATA_L[7]),
    .B(_3329_),
    .C(DMEM_DATA_L[23]),
    .D(_3350_),
    .Y(_3489_)
);

NAND3X1 _14193_ (
    .A(_0__1_bF$buf5),
    .B(DMEM_DATA_L[31]),
    .C(_0__0_bF$buf2),
    .Y(_3490_)
);

INVX1 _14194_ (
    .A(_3490_),
    .Y(_3491_)
);

AOI21X1 _14195_ (
    .A(_3341_),
    .B(DMEM_DATA_L[15]),
    .C(_3491_),
    .Y(_3492_)
);

NAND2X1 _14196_ (
    .A(_3489_),
    .B(_3492_),
    .Y(\datapath.memoryinterface.byte_size_load.byteval [7])
);

INVX1 _14197_ (
    .A(\datapath.programcounter.pc_mux [0]),
    .Y(_3493_)
);

NAND2X1 _14198_ (
    .A(\datapath.programcounter.pc [0]),
    .B(1'h0),
    .Y(_3494_)
);

OAI21X1 _14199_ (
    .A(1'h0),
    .B(_3493_),
    .C(_3494_),
    .Y(\datapath.programcounter._1_ [0])
);

INVX1 _14200_ (
    .A(\datapath.programcounter.pc_mux [1]),
    .Y(_3495_)
);

NAND2X1 _14201_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc [1]),
    .Y(_3496_)
);

OAI21X1 _14202_ (
    .A(1'h0),
    .B(_3495_),
    .C(_3496_),
    .Y(\datapath.programcounter._1_ [1])
);

INVX2 _14203_ (
    .A(\datapath.programcounter.pc [2]),
    .Y(\datapath.nextpc [2])
);

NOR2X1 _14204_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [2]),
    .Y(_3497_)
);

AOI21X1 _14205_ (
    .A(1'h0),
    .B(\datapath.nextpc [2]),
    .C(_3497_),
    .Y(\datapath.programcounter._1_ [2])
);

INVX1 _14206_ (
    .A(\datapath.programcounter.pc [3]),
    .Y(_3498_)
);

NOR2X1 _14207_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [3]),
    .Y(_3499_)
);

AOI21X1 _14208_ (
    .A(1'h0),
    .B(_3498_),
    .C(_3499_),
    .Y(\datapath.programcounter._1_ [3])
);

INVX1 _14209_ (
    .A(\datapath.programcounter.pc [4]),
    .Y(_3500_)
);

NOR2X1 _14210_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [4]),
    .Y(_3501_)
);

AOI21X1 _14211_ (
    .A(1'h0),
    .B(_3500_),
    .C(_3501_),
    .Y(\datapath.programcounter._1_ [4])
);

INVX1 _14212_ (
    .A(\datapath.programcounter.pc [5]),
    .Y(_3502_)
);

NOR2X1 _14213_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [5]),
    .Y(_3503_)
);

AOI21X1 _14214_ (
    .A(1'h0),
    .B(_3502_),
    .C(_3503_),
    .Y(\datapath.programcounter._1_ [5])
);

INVX1 _14215_ (
    .A(\datapath.programcounter.pc [6]),
    .Y(_3504_)
);

NOR2X1 _14216_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [6]),
    .Y(_3505_)
);

AOI21X1 _14217_ (
    .A(1'h0),
    .B(_3504_),
    .C(_3505_),
    .Y(\datapath.programcounter._1_ [6])
);

INVX1 _14218_ (
    .A(\datapath.programcounter.pc [7]),
    .Y(_3506_)
);

NOR2X1 _14219_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [7]),
    .Y(_3507_)
);

AOI21X1 _14220_ (
    .A(1'h0),
    .B(_3506_),
    .C(_3507_),
    .Y(\datapath.programcounter._1_ [7])
);

INVX1 _14221_ (
    .A(\datapath.programcounter.pc [8]),
    .Y(_3508_)
);

NOR2X1 _14222_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [8]),
    .Y(_3509_)
);

AOI21X1 _14223_ (
    .A(1'h0),
    .B(_3508_),
    .C(_3509_),
    .Y(\datapath.programcounter._1_ [8])
);

INVX1 _14224_ (
    .A(\datapath.programcounter.pc [9]),
    .Y(_3510_)
);

NOR2X1 _14225_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [9]),
    .Y(_3511_)
);

AOI21X1 _14226_ (
    .A(1'h0),
    .B(_3510_),
    .C(_3511_),
    .Y(\datapath.programcounter._1_ [9])
);

INVX1 _14227_ (
    .A(\datapath.programcounter.pc [10]),
    .Y(_3512_)
);

NOR2X1 _14228_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [10]),
    .Y(_3513_)
);

AOI21X1 _14229_ (
    .A(1'h0),
    .B(_3512_),
    .C(_3513_),
    .Y(\datapath.programcounter._1_ [10])
);

INVX1 _14230_ (
    .A(\datapath.programcounter.pc [11]),
    .Y(_3514_)
);

NOR2X1 _14231_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [11]),
    .Y(_3515_)
);

AOI21X1 _14232_ (
    .A(1'h0),
    .B(_3514_),
    .C(_3515_),
    .Y(\datapath.programcounter._1_ [11])
);

INVX1 _14233_ (
    .A(\datapath.programcounter.pc [12]),
    .Y(_3516_)
);

NOR2X1 _14234_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [12]),
    .Y(_3517_)
);

AOI21X1 _14235_ (
    .A(1'h0),
    .B(_3516_),
    .C(_3517_),
    .Y(\datapath.programcounter._1_ [12])
);

INVX1 _14236_ (
    .A(\datapath.programcounter.pc [13]),
    .Y(_3518_)
);

NOR2X1 _14237_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [13]),
    .Y(_3519_)
);

AOI21X1 _14238_ (
    .A(1'h0),
    .B(_3518_),
    .C(_3519_),
    .Y(\datapath.programcounter._1_ [13])
);

INVX1 _14239_ (
    .A(\datapath.programcounter.pc [14]),
    .Y(_3520_)
);

NOR2X1 _14240_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [14]),
    .Y(_3521_)
);

AOI21X1 _14241_ (
    .A(1'h0),
    .B(_3520_),
    .C(_3521_),
    .Y(\datapath.programcounter._1_ [14])
);

INVX1 _14242_ (
    .A(\datapath.programcounter.pc [15]),
    .Y(_3522_)
);

NOR2X1 _14243_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [15]),
    .Y(_3523_)
);

AOI21X1 _14244_ (
    .A(1'h0),
    .B(_3522_),
    .C(_3523_),
    .Y(\datapath.programcounter._1_ [15])
);

INVX1 _14245_ (
    .A(\datapath.programcounter.pc [16]),
    .Y(_3524_)
);

NOR2X1 _14246_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [16]),
    .Y(_3525_)
);

AOI21X1 _14247_ (
    .A(1'h0),
    .B(_3524_),
    .C(_3525_),
    .Y(\datapath.programcounter._1_ [16])
);

INVX1 _14248_ (
    .A(\datapath.programcounter.pc [17]),
    .Y(_3526_)
);

NOR2X1 _14249_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [17]),
    .Y(_3527_)
);

AOI21X1 _14250_ (
    .A(1'h0),
    .B(_3526_),
    .C(_3527_),
    .Y(\datapath.programcounter._1_ [17])
);

INVX2 _14251_ (
    .A(\datapath.programcounter.pc [18]),
    .Y(_3528_)
);

NOR2X1 _14252_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [18]),
    .Y(_3529_)
);

AOI21X1 _14253_ (
    .A(1'h0),
    .B(_3528_),
    .C(_3529_),
    .Y(\datapath.programcounter._1_ [18])
);

INVX1 _14254_ (
    .A(\datapath.programcounter.pc [19]),
    .Y(_3530_)
);

NOR2X1 _14255_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [19]),
    .Y(_3531_)
);

AOI21X1 _14256_ (
    .A(1'h0),
    .B(_3530_),
    .C(_3531_),
    .Y(\datapath.programcounter._1_ [19])
);

INVX1 _14257_ (
    .A(\datapath.programcounter.pc [20]),
    .Y(_3532_)
);

NOR2X1 _14258_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [20]),
    .Y(_3533_)
);

AOI21X1 _14259_ (
    .A(1'h0),
    .B(_3532_),
    .C(_3533_),
    .Y(\datapath.programcounter._1_ [20])
);

INVX1 _14260_ (
    .A(\datapath.programcounter.pc [21]),
    .Y(_3534_)
);

NOR2X1 _14261_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [21]),
    .Y(_3535_)
);

AOI21X1 _14262_ (
    .A(1'h0),
    .B(_3534_),
    .C(_3535_),
    .Y(\datapath.programcounter._1_ [21])
);

INVX2 _14263_ (
    .A(\datapath.programcounter.pc [22]),
    .Y(_3536_)
);

NOR2X1 _14264_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [22]),
    .Y(_3537_)
);

AOI21X1 _14265_ (
    .A(1'h0),
    .B(_3536_),
    .C(_3537_),
    .Y(\datapath.programcounter._1_ [22])
);

INVX1 _14266_ (
    .A(\datapath.programcounter.pc [23]),
    .Y(_3538_)
);

NOR2X1 _14267_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [23]),
    .Y(_3539_)
);

AOI21X1 _14268_ (
    .A(1'h0),
    .B(_3538_),
    .C(_3539_),
    .Y(\datapath.programcounter._1_ [23])
);

INVX1 _14269_ (
    .A(\datapath.programcounter.pc [24]),
    .Y(_3540_)
);

NOR2X1 _14270_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [24]),
    .Y(_3541_)
);

AOI21X1 _14271_ (
    .A(1'h0),
    .B(_3540_),
    .C(_3541_),
    .Y(\datapath.programcounter._1_ [24])
);

INVX1 _14272_ (
    .A(\datapath.programcounter.pc [25]),
    .Y(_3542_)
);

NOR2X1 _14273_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [25]),
    .Y(_3543_)
);

AOI21X1 _14274_ (
    .A(1'h0),
    .B(_3542_),
    .C(_3543_),
    .Y(\datapath.programcounter._1_ [25])
);

INVX1 _14275_ (
    .A(\datapath.programcounter.pc [26]),
    .Y(_3544_)
);

NOR2X1 _14276_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [26]),
    .Y(_3545_)
);

AOI21X1 _14277_ (
    .A(1'h0),
    .B(_3544_),
    .C(_3545_),
    .Y(\datapath.programcounter._1_ [26])
);

INVX1 _14278_ (
    .A(\datapath.programcounter.pc [27]),
    .Y(_3546_)
);

NOR2X1 _14279_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [27]),
    .Y(_3547_)
);

AOI21X1 _14280_ (
    .A(1'h0),
    .B(_3546_),
    .C(_3547_),
    .Y(\datapath.programcounter._1_ [27])
);

INVX2 _14281_ (
    .A(\datapath.programcounter.pc [28]),
    .Y(_3548_)
);

NOR2X1 _14282_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [28]),
    .Y(_3549_)
);

AOI21X1 _14283_ (
    .A(1'h0),
    .B(_3548_),
    .C(_3549_),
    .Y(\datapath.programcounter._1_ [28])
);

INVX1 _14284_ (
    .A(\datapath.programcounter.pc [29]),
    .Y(_3550_)
);

NOR2X1 _14285_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [29]),
    .Y(_3551_)
);

AOI21X1 _14286_ (
    .A(1'h0),
    .B(_3550_),
    .C(_3551_),
    .Y(\datapath.programcounter._1_ [29])
);

INVX1 _14287_ (
    .A(\datapath.programcounter.pc [30]),
    .Y(_3552_)
);

NOR2X1 _14288_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [30]),
    .Y(_3553_)
);

AOI21X1 _14289_ (
    .A(1'h0),
    .B(_3552_),
    .C(_3553_),
    .Y(\datapath.programcounter._1_ [30])
);

INVX1 _14290_ (
    .A(\datapath.programcounter.pc [31]),
    .Y(_3554_)
);

NOR2X1 _14291_ (
    .A(1'h0),
    .B(\datapath.programcounter.pc_mux [31]),
    .Y(_3555_)
);

AOI21X1 _14292_ (
    .A(1'h0),
    .B(_3554_),
    .C(_3555_),
    .Y(\datapath.programcounter._1_ [31])
);

INVX1 _14293_ (
    .A(\datapath._36_ ),
    .Y(_3556_)
);

NOR2X1 _14294_ (
    .A(\datapath._34_ ),
    .B(_3556_),
    .Y(_3557_)
);

NOR2X1 _14295_ (
    .A(\datapath._34_ ),
    .B(\datapath._36_ ),
    .Y(_3558_)
);

AOI22X1 _14296_ (
    .A(\datapath.programcounter.pc [0]),
    .B(_3558__bF$buf4),
    .C(1'h0),
    .D(_3557__bF$buf4),
    .Y(_3559_)
);

INVX1 _14297_ (
    .A(\datapath._34_ ),
    .Y(_3560_)
);

NOR2X1 _14298_ (
    .A(\datapath._36_ ),
    .B(_3560_),
    .Y(_3561_)
);

NAND2X1 _14299_ (
    .A(\datapath.programcounter.jumps [0]),
    .B(_3561__bF$buf4),
    .Y(_3562_)
);

NOR2X1 _14300_ (
    .A(_3560_),
    .B(_3556_),
    .Y(_3563_)
);

NAND2X1 _14301_ (
    .A(1'h0),
    .B(_3563__bF$buf4),
    .Y(_3564_)
);

NAND3X1 _14302_ (
    .A(_3562_),
    .B(_3564_),
    .C(_3559_),
    .Y(\datapath.programcounter.pc_mux [0])
);

AOI22X1 _14303_ (
    .A(\datapath.programcounter.pc [1]),
    .B(_3558__bF$buf3),
    .C(_0__1_bF$buf4),
    .D(_3557__bF$buf3),
    .Y(_3565_)
);

NAND2X1 _14304_ (
    .A(\datapath.programcounter.jumps [1]),
    .B(_3561__bF$buf3),
    .Y(_3566_)
);

NAND2X1 _14305_ (
    .A(1'h0),
    .B(_3563__bF$buf3),
    .Y(_3567_)
);

NAND3X1 _14306_ (
    .A(_3566_),
    .B(_3567_),
    .C(_3565_),
    .Y(\datapath.programcounter.pc_mux [1])
);

AOI22X1 _14307_ (
    .A(\datapath.nextpc [2]),
    .B(_3558__bF$buf2),
    .C(_0_[2]),
    .D(_3557__bF$buf2),
    .Y(_3568_)
);

NAND2X1 _14308_ (
    .A(\datapath.programcounter.jumps [2]),
    .B(_3561__bF$buf2),
    .Y(_3569_)
);

NAND2X1 _14309_ (
    .A(\datapath.csr.csr_pcaddr [2]),
    .B(_3563__bF$buf2),
    .Y(_3570_)
);

NAND3X1 _14310_ (
    .A(_3569_),
    .B(_3570_),
    .C(_3568_),
    .Y(\datapath.programcounter.pc_mux [2])
);

NOR2X1 _14311_ (
    .A(\datapath.nextpc [2]),
    .B(_3498_),
    .Y(_3571_)
);

NOR2X1 _14312_ (
    .A(\datapath.programcounter.pc [2]),
    .B(\datapath.programcounter.pc [3]),
    .Y(_3572_)
);

NOR2X1 _14313_ (
    .A(_3572_),
    .B(_3571_),
    .Y(\datapath.nextpc [3])
);

NAND2X1 _14314_ (
    .A(_3558__bF$buf1),
    .B(\datapath.nextpc [3]),
    .Y(_3573_)
);

NAND2X1 _14315_ (
    .A(\datapath.programcounter.jumps [3]),
    .B(_3561__bF$buf1),
    .Y(_3574_)
);

AOI22X1 _14316_ (
    .A(_3557__bF$buf1),
    .B(_0_[3]),
    .C(\datapath.csr.csr_pcaddr [3]),
    .D(_3563__bF$buf1),
    .Y(_3575_)
);

NAND3X1 _14317_ (
    .A(_3574_),
    .B(_3575_),
    .C(_3573_),
    .Y(\datapath.programcounter.pc_mux [3])
);

NAND3X1 _14318_ (
    .A(\datapath.programcounter.pc [2]),
    .B(\datapath.programcounter.pc [3]),
    .C(\datapath.programcounter.pc [4]),
    .Y(_3576_)
);

INVX1 _14319_ (
    .A(_3576_),
    .Y(_3577_)
);

NOR2X1 _14320_ (
    .A(\datapath.programcounter.pc [4]),
    .B(_3571_),
    .Y(_3578_)
);

NOR2X1 _14321_ (
    .A(_3577_),
    .B(_3578_),
    .Y(\datapath.nextpc [4])
);

NAND2X1 _14322_ (
    .A(_3558__bF$buf0),
    .B(\datapath.nextpc [4]),
    .Y(_3579_)
);

NAND2X1 _14323_ (
    .A(\datapath.programcounter.jumps [4]),
    .B(_3561__bF$buf0),
    .Y(_3580_)
);

AOI22X1 _14324_ (
    .A(_3557__bF$buf0),
    .B(_0_[4]),
    .C(\datapath.csr.csr_pcaddr [4]),
    .D(_3563__bF$buf0),
    .Y(_3581_)
);

NAND3X1 _14325_ (
    .A(_3580_),
    .B(_3581_),
    .C(_3579_),
    .Y(\datapath.programcounter.pc_mux [4])
);

XNOR2X1 _14326_ (
    .A(_3576_),
    .B(\datapath.programcounter.pc [5]),
    .Y(\datapath.nextpc [5])
);

NAND2X1 _14327_ (
    .A(_3558__bF$buf4),
    .B(\datapath.nextpc [5]),
    .Y(_3582_)
);

NAND2X1 _14328_ (
    .A(\datapath.programcounter.jumps [5]),
    .B(_3561__bF$buf4),
    .Y(_3583_)
);

AOI22X1 _14329_ (
    .A(_3557__bF$buf4),
    .B(_0_[5]),
    .C(\datapath.csr.csr_pcaddr [5]),
    .D(_3563__bF$buf4),
    .Y(_3584_)
);

NAND3X1 _14330_ (
    .A(_3583_),
    .B(_3584_),
    .C(_3582_),
    .Y(\datapath.programcounter.pc_mux [5])
);

NAND2X1 _14331_ (
    .A(\datapath.programcounter.pc [5]),
    .B(\datapath.programcounter.pc [6]),
    .Y(_3585_)
);

OR2X2 _14332_ (
    .A(_3576_),
    .B(_3585_),
    .Y(_3586_)
);

OAI21X1 _14333_ (
    .A(_3502_),
    .B(_3576_),
    .C(_3504_),
    .Y(_3587_)
);

AND2X2 _14334_ (
    .A(_3586_),
    .B(_3587_),
    .Y(\datapath.nextpc [6])
);

NAND2X1 _14335_ (
    .A(_3558__bF$buf3),
    .B(\datapath.nextpc [6]),
    .Y(_3588_)
);

NAND2X1 _14336_ (
    .A(\datapath.programcounter.jumps [6]),
    .B(_3561__bF$buf3),
    .Y(_3589_)
);

AOI22X1 _14337_ (
    .A(_3557__bF$buf3),
    .B(_0_[6]),
    .C(\datapath.csr.csr_pcaddr [6]),
    .D(_3563__bF$buf3),
    .Y(_3590_)
);

NAND3X1 _14338_ (
    .A(_3589_),
    .B(_3590_),
    .C(_3588_),
    .Y(\datapath.programcounter.pc_mux [6])
);

XNOR2X1 _14339_ (
    .A(_3586_),
    .B(\datapath.programcounter.pc [7]),
    .Y(\datapath.nextpc [7])
);

NAND2X1 _14340_ (
    .A(\datapath.programcounter.jumps [7]),
    .B(_3561__bF$buf2),
    .Y(_3591_)
);

NAND2X1 _14341_ (
    .A(\datapath.csr.csr_pcaddr [7]),
    .B(_3563__bF$buf2),
    .Y(_3592_)
);

AOI22X1 _14342_ (
    .A(_0_[7]),
    .B(_3557__bF$buf2),
    .C(_3558__bF$buf2),
    .D(\datapath.nextpc [7]),
    .Y(_3593_)
);

NAND3X1 _14343_ (
    .A(_3591_),
    .B(_3592_),
    .C(_3593_),
    .Y(\datapath.programcounter.pc_mux [7])
);

NAND3X1 _14344_ (
    .A(\datapath.programcounter.pc [5]),
    .B(\datapath.programcounter.pc [6]),
    .C(\datapath.programcounter.pc [7]),
    .Y(_3594_)
);

OAI21X1 _14345_ (
    .A(_3576_),
    .B(_3594_),
    .C(_3508_),
    .Y(_3595_)
);

NOR2X1 _14346_ (
    .A(_3576_),
    .B(_3594_),
    .Y(_3596_)
);

NAND2X1 _14347_ (
    .A(\datapath.programcounter.pc [8]),
    .B(_3596_),
    .Y(_3597_)
);

AND2X2 _14348_ (
    .A(_3597_),
    .B(_3595_),
    .Y(\datapath.nextpc [8])
);

NAND2X1 _14349_ (
    .A(\datapath.programcounter.jumps [8]),
    .B(_3561__bF$buf1),
    .Y(_3598_)
);

NAND2X1 _14350_ (
    .A(\datapath.csr.csr_pcaddr [8]),
    .B(_3563__bF$buf1),
    .Y(_3599_)
);

AOI22X1 _14351_ (
    .A(_0_[8]),
    .B(_3557__bF$buf1),
    .C(_3558__bF$buf1),
    .D(\datapath.nextpc [8]),
    .Y(_3600_)
);

NAND3X1 _14352_ (
    .A(_3598_),
    .B(_3599_),
    .C(_3600_),
    .Y(\datapath.programcounter.pc_mux [8])
);

XNOR2X1 _14353_ (
    .A(_3597_),
    .B(\datapath.programcounter.pc [9]),
    .Y(\datapath.nextpc [9])
);

NAND2X1 _14354_ (
    .A(\datapath.programcounter.jumps [9]),
    .B(_3561__bF$buf0),
    .Y(_3601_)
);

NAND2X1 _14355_ (
    .A(\datapath.csr.csr_pcaddr [9]),
    .B(_3563__bF$buf0),
    .Y(_3602_)
);

AOI22X1 _14356_ (
    .A(_0_[9]),
    .B(_3557__bF$buf0),
    .C(_3558__bF$buf0),
    .D(\datapath.nextpc [9]),
    .Y(_3603_)
);

NAND3X1 _14357_ (
    .A(_3601_),
    .B(_3602_),
    .C(_3603_),
    .Y(\datapath.programcounter.pc_mux [9])
);

OAI21X1 _14358_ (
    .A(_3510_),
    .B(_3597_),
    .C(_3512_),
    .Y(_3604_)
);

NOR2X1 _14359_ (
    .A(_3506_),
    .B(_3586_),
    .Y(_3605_)
);

NAND2X1 _14360_ (
    .A(\datapath.programcounter.pc [8]),
    .B(\datapath.programcounter.pc [9]),
    .Y(_3606_)
);

INVX1 _14361_ (
    .A(_3606_),
    .Y(_3607_)
);

NAND3X1 _14362_ (
    .A(\datapath.programcounter.pc [10]),
    .B(_3607_),
    .C(_3605_),
    .Y(_3608_)
);

AND2X2 _14363_ (
    .A(_3608_),
    .B(_3604_),
    .Y(\datapath.nextpc [10])
);

NAND2X1 _14364_ (
    .A(\datapath.programcounter.jumps [10]),
    .B(_3561__bF$buf4),
    .Y(_3609_)
);

NAND2X1 _14365_ (
    .A(\datapath.csr.csr_pcaddr [10]),
    .B(_3563__bF$buf4),
    .Y(_3610_)
);

AOI22X1 _14366_ (
    .A(_0_[10]),
    .B(_3557__bF$buf4),
    .C(_3558__bF$buf4),
    .D(\datapath.nextpc [10]),
    .Y(_3611_)
);

NAND3X1 _14367_ (
    .A(_3609_),
    .B(_3610_),
    .C(_3611_),
    .Y(\datapath.programcounter.pc_mux [10])
);

NAND2X1 _14368_ (
    .A(_3514_),
    .B(_3608_),
    .Y(_3612_)
);

OR2X2 _14369_ (
    .A(_3608_),
    .B(_3514_),
    .Y(_3613_)
);

AND2X2 _14370_ (
    .A(_3613_),
    .B(_3612_),
    .Y(\datapath.nextpc [11])
);

NAND3X1 _14371_ (
    .A(_3558__bF$buf3),
    .B(_3612_),
    .C(_3613_),
    .Y(_3614_)
);

NAND2X1 _14372_ (
    .A(\datapath.programcounter.jumps [11]),
    .B(_3561__bF$buf3),
    .Y(_3615_)
);

AOI22X1 _14373_ (
    .A(_3557__bF$buf3),
    .B(_0_[11]),
    .C(\datapath.csr.csr_pcaddr [11]),
    .D(_3563__bF$buf3),
    .Y(_3616_)
);

NAND3X1 _14374_ (
    .A(_3615_),
    .B(_3616_),
    .C(_3614_),
    .Y(\datapath.programcounter.pc_mux [11])
);

NAND2X1 _14375_ (
    .A(\datapath.programcounter.pc [4]),
    .B(\datapath.programcounter.pc [5]),
    .Y(_3617_)
);

NAND2X1 _14376_ (
    .A(\datapath.programcounter.pc [6]),
    .B(\datapath.programcounter.pc [7]),
    .Y(_3618_)
);

NOR2X1 _14377_ (
    .A(_3617_),
    .B(_3618_),
    .Y(_3619_)
);

NAND2X1 _14378_ (
    .A(\datapath.programcounter.pc [10]),
    .B(\datapath.programcounter.pc [11]),
    .Y(_3620_)
);

NOR2X1 _14379_ (
    .A(_3606_),
    .B(_3620_),
    .Y(_3621_)
);

NAND3X1 _14380_ (
    .A(_3571_),
    .B(_3619_),
    .C(_3621_),
    .Y(_3622_)
);

XNOR2X1 _14381_ (
    .A(_3622_),
    .B(\datapath.programcounter.pc [12]),
    .Y(\datapath.nextpc [12])
);

NAND2X1 _14382_ (
    .A(\datapath.programcounter.jumps [12]),
    .B(_3561__bF$buf2),
    .Y(_3623_)
);

NAND2X1 _14383_ (
    .A(\datapath.csr.csr_pcaddr [12]),
    .B(_3563__bF$buf2),
    .Y(_3624_)
);

AOI22X1 _14384_ (
    .A(_0_[12]),
    .B(_3557__bF$buf2),
    .C(_3558__bF$buf2),
    .D(\datapath.nextpc [12]),
    .Y(_3625_)
);

NAND3X1 _14385_ (
    .A(_3623_),
    .B(_3624_),
    .C(_3625_),
    .Y(\datapath.programcounter.pc_mux [12])
);

NAND3X1 _14386_ (
    .A(\datapath.programcounter.pc [12]),
    .B(_3621_),
    .C(_3596_),
    .Y(_3626_)
);

AND2X2 _14387_ (
    .A(_3626_),
    .B(\datapath.programcounter.pc [13]),
    .Y(_3627_)
);

NOR2X1 _14388_ (
    .A(\datapath.programcounter.pc [13]),
    .B(_3626_),
    .Y(_3628_)
);

OR2X2 _14389_ (
    .A(_3627_),
    .B(_3628_),
    .Y(\datapath.nextpc [13])
);

OAI21X1 _14390_ (
    .A(_3628_),
    .B(_3627_),
    .C(_3558__bF$buf1),
    .Y(_3629_)
);

NAND2X1 _14391_ (
    .A(\datapath.programcounter.jumps [13]),
    .B(_3561__bF$buf1),
    .Y(_3630_)
);

AOI22X1 _14392_ (
    .A(_3557__bF$buf1),
    .B(_0_[13]),
    .C(\datapath.csr.csr_pcaddr [13]),
    .D(_3563__bF$buf1),
    .Y(_3631_)
);

NAND3X1 _14393_ (
    .A(_3630_),
    .B(_3631_),
    .C(_3629_),
    .Y(\datapath.programcounter.pc_mux [13])
);

OAI21X1 _14394_ (
    .A(_3518_),
    .B(_3626_),
    .C(_3520_),
    .Y(_3632_)
);

NOR2X1 _14395_ (
    .A(_3518_),
    .B(_3626_),
    .Y(_3633_)
);

NAND2X1 _14396_ (
    .A(\datapath.programcounter.pc [14]),
    .B(_3633_),
    .Y(_3634_)
);

AND2X2 _14397_ (
    .A(_3634_),
    .B(_3632_),
    .Y(\datapath.nextpc [14])
);

NAND2X1 _14398_ (
    .A(_3558__bF$buf0),
    .B(\datapath.nextpc [14]),
    .Y(_3635_)
);

NAND2X1 _14399_ (
    .A(\datapath.programcounter.jumps [14]),
    .B(_3561__bF$buf0),
    .Y(_3636_)
);

AOI22X1 _14400_ (
    .A(_3557__bF$buf0),
    .B(_0_[14]),
    .C(\datapath.csr.csr_pcaddr [14]),
    .D(_3563__bF$buf0),
    .Y(_3637_)
);

NAND3X1 _14401_ (
    .A(_3636_),
    .B(_3637_),
    .C(_3635_),
    .Y(\datapath.programcounter.pc_mux [14])
);

NAND2X1 _14402_ (
    .A(\datapath.programcounter.pc [12]),
    .B(\datapath.programcounter.pc [13]),
    .Y(_3638_)
);

NOR2X1 _14403_ (
    .A(_3638_),
    .B(_3622_),
    .Y(_3639_)
);

AOI21X1 _14404_ (
    .A(_3639_),
    .B(\datapath.programcounter.pc [14]),
    .C(_3522_),
    .Y(_3640_)
);

NAND2X1 _14405_ (
    .A(\datapath.programcounter.pc [14]),
    .B(_3639_),
    .Y(_3641_)
);

NOR2X1 _14406_ (
    .A(\datapath.programcounter.pc [15]),
    .B(_3641_),
    .Y(_3642_)
);

OR2X2 _14407_ (
    .A(_3642_),
    .B(_3640_),
    .Y(\datapath.nextpc [15])
);

OAI21X1 _14408_ (
    .A(_3640_),
    .B(_3642_),
    .C(_3558__bF$buf4),
    .Y(_3643_)
);

NAND2X1 _14409_ (
    .A(\datapath.csr.csr_pcaddr [15]),
    .B(_3563__bF$buf4),
    .Y(_3644_)
);

AOI22X1 _14410_ (
    .A(_3557__bF$buf4),
    .B(_0_[15]),
    .C(\datapath.programcounter.jumps [15]),
    .D(_3561__bF$buf4),
    .Y(_3645_)
);

NAND3X1 _14411_ (
    .A(_3644_),
    .B(_3645_),
    .C(_3643_),
    .Y(\datapath.programcounter.pc_mux [15])
);

OR2X2 _14412_ (
    .A(_3576_),
    .B(_3594_),
    .Y(_3646_)
);

NAND2X1 _14413_ (
    .A(\datapath.programcounter.pc [14]),
    .B(\datapath.programcounter.pc [15]),
    .Y(_3647_)
);

NOR2X1 _14414_ (
    .A(_3638_),
    .B(_3647_),
    .Y(_3648_)
);

NAND2X1 _14415_ (
    .A(_3621_),
    .B(_3648_),
    .Y(_3649_)
);

OAI21X1 _14416_ (
    .A(_3646_),
    .B(_3649_),
    .C(_3524_),
    .Y(_3650_)
);

NOR2X1 _14417_ (
    .A(_3646_),
    .B(_3649_),
    .Y(_3651_)
);

NAND2X1 _14418_ (
    .A(\datapath.programcounter.pc [16]),
    .B(_3651_),
    .Y(_3652_)
);

AND2X2 _14419_ (
    .A(_3652_),
    .B(_3650_),
    .Y(\datapath.nextpc [16])
);

NAND2X1 _14420_ (
    .A(\datapath.programcounter.jumps [16]),
    .B(_3561__bF$buf3),
    .Y(_3653_)
);

NAND2X1 _14421_ (
    .A(\datapath.csr.csr_pcaddr [16]),
    .B(_3563__bF$buf3),
    .Y(_3654_)
);

AOI22X1 _14422_ (
    .A(_0_[16]),
    .B(_3557__bF$buf3),
    .C(_3558__bF$buf3),
    .D(\datapath.nextpc [16]),
    .Y(_3655_)
);

NAND3X1 _14423_ (
    .A(_3653_),
    .B(_3654_),
    .C(_3655_),
    .Y(\datapath.programcounter.pc_mux [16])
);

AOI21X1 _14424_ (
    .A(_3651_),
    .B(\datapath.programcounter.pc [16]),
    .C(_3526_),
    .Y(_3656_)
);

NOR2X1 _14425_ (
    .A(\datapath.programcounter.pc [17]),
    .B(_3652_),
    .Y(_3657_)
);

OR2X2 _14426_ (
    .A(_3657_),
    .B(_3656_),
    .Y(\datapath.nextpc [17])
);

OAI21X1 _14427_ (
    .A(_3656_),
    .B(_3657_),
    .C(_3558__bF$buf2),
    .Y(_3658_)
);

NAND2X1 _14428_ (
    .A(\datapath.programcounter.jumps [17]),
    .B(_3561__bF$buf2),
    .Y(_3659_)
);

AOI22X1 _14429_ (
    .A(_3557__bF$buf2),
    .B(_0_[17]),
    .C(\datapath.csr.csr_pcaddr [17]),
    .D(_3563__bF$buf2),
    .Y(_3660_)
);

NAND3X1 _14430_ (
    .A(_3659_),
    .B(_3660_),
    .C(_3658_),
    .Y(\datapath.programcounter.pc_mux [17])
);

NAND3X1 _14431_ (
    .A(\datapath.programcounter.pc [7]),
    .B(\datapath.programcounter.pc [14]),
    .C(\datapath.programcounter.pc [15]),
    .Y(_3661_)
);

NOR3X1 _14432_ (
    .A(_3585_),
    .B(_3638_),
    .C(_3661_),
    .Y(_3662_)
);

NOR3X1 _14433_ (
    .A(_3606_),
    .B(_3620_),
    .C(_3576_),
    .Y(_3663_)
);

NAND2X1 _14434_ (
    .A(_3662_),
    .B(_3663_),
    .Y(_3664_)
);

NAND2X1 _14435_ (
    .A(\datapath.programcounter.pc [16]),
    .B(\datapath.programcounter.pc [17]),
    .Y(_3665_)
);

OAI21X1 _14436_ (
    .A(_3665_),
    .B(_3664_),
    .C(_3528_),
    .Y(_3666_)
);

INVX1 _14437_ (
    .A(_3665_),
    .Y(_3667_)
);

NAND3X1 _14438_ (
    .A(_3667_),
    .B(_3662_),
    .C(_3663_),
    .Y(_3668_)
);

NOR2X1 _14439_ (
    .A(_3528_),
    .B(_3668_),
    .Y(_3669_)
);

INVX1 _14440_ (
    .A(_3669_),
    .Y(_3670_)
);

AND2X2 _14441_ (
    .A(_3670_),
    .B(_3666_),
    .Y(\datapath.nextpc [18])
);

NAND2X1 _14442_ (
    .A(_3558__bF$buf1),
    .B(\datapath.nextpc [18]),
    .Y(_3671_)
);

NAND2X1 _14443_ (
    .A(\datapath.programcounter.jumps [18]),
    .B(_3561__bF$buf1),
    .Y(_3672_)
);

AOI22X1 _14444_ (
    .A(_3557__bF$buf1),
    .B(_0_[18]),
    .C(\datapath.csr.csr_pcaddr [18]),
    .D(_3563__bF$buf1),
    .Y(_3673_)
);

NAND3X1 _14445_ (
    .A(_3672_),
    .B(_3673_),
    .C(_3671_),
    .Y(\datapath.programcounter.pc_mux [18])
);

OAI21X1 _14446_ (
    .A(_3528_),
    .B(_3668_),
    .C(_3530_),
    .Y(_3674_)
);

NAND2X1 _14447_ (
    .A(\datapath.programcounter.pc [19]),
    .B(_3669_),
    .Y(_3675_)
);

AND2X2 _14448_ (
    .A(_3675_),
    .B(_3674_),
    .Y(\datapath.nextpc [19])
);

NAND3X1 _14449_ (
    .A(_3558__bF$buf0),
    .B(_3674_),
    .C(_3675_),
    .Y(_3676_)
);

NAND2X1 _14450_ (
    .A(\datapath.programcounter.jumps [19]),
    .B(_3561__bF$buf0),
    .Y(_3677_)
);

AOI22X1 _14451_ (
    .A(_3557__bF$buf0),
    .B(_0_[19]),
    .C(\datapath.csr.csr_pcaddr [19]),
    .D(_3563__bF$buf0),
    .Y(_3678_)
);

NAND3X1 _14452_ (
    .A(_3677_),
    .B(_3678_),
    .C(_3676_),
    .Y(\datapath.programcounter.pc_mux [19])
);

NAND2X1 _14453_ (
    .A(\datapath.programcounter.pc [18]),
    .B(\datapath.programcounter.pc [19]),
    .Y(_3679_)
);

NOR2X1 _14454_ (
    .A(_3665_),
    .B(_3679_),
    .Y(_3680_)
);

NAND3X1 _14455_ (
    .A(_3680_),
    .B(_3662_),
    .C(_3663_),
    .Y(_3681_)
);

XNOR2X1 _14456_ (
    .A(_3681_),
    .B(\datapath.programcounter.pc [20]),
    .Y(\datapath.nextpc [20])
);

NAND2X1 _14457_ (
    .A(\datapath.programcounter.jumps [20]),
    .B(_3561__bF$buf4),
    .Y(_3682_)
);

NAND2X1 _14458_ (
    .A(\datapath.csr.csr_pcaddr [20]),
    .B(_3563__bF$buf4),
    .Y(_3683_)
);

AOI22X1 _14459_ (
    .A(_0_[20]),
    .B(_3557__bF$buf4),
    .C(_3558__bF$buf4),
    .D(\datapath.nextpc [20]),
    .Y(_3684_)
);

NAND3X1 _14460_ (
    .A(_3682_),
    .B(_3683_),
    .C(_3684_),
    .Y(\datapath.programcounter.pc_mux [20])
);

OAI21X1 _14461_ (
    .A(_3532_),
    .B(_3681_),
    .C(_3534_),
    .Y(_3685_)
);

NAND2X1 _14462_ (
    .A(\datapath.programcounter.pc [20]),
    .B(\datapath.programcounter.pc [21]),
    .Y(_3686_)
);

OR2X2 _14463_ (
    .A(_3681_),
    .B(_3686_),
    .Y(_3687_)
);

AND2X2 _14464_ (
    .A(_3687_),
    .B(_3685_),
    .Y(\datapath.nextpc [21])
);

NAND2X1 _14465_ (
    .A(\datapath.programcounter.jumps [21]),
    .B(_3561__bF$buf3),
    .Y(_3688_)
);

NAND2X1 _14466_ (
    .A(\datapath.csr.csr_pcaddr [21]),
    .B(_3563__bF$buf3),
    .Y(_3689_)
);

AOI22X1 _14467_ (
    .A(_0_[21]),
    .B(_3557__bF$buf3),
    .C(_3558__bF$buf3),
    .D(\datapath.nextpc [21]),
    .Y(_3690_)
);

NAND3X1 _14468_ (
    .A(_3688_),
    .B(_3689_),
    .C(_3690_),
    .Y(\datapath.programcounter.pc_mux [21])
);

NOR2X1 _14469_ (
    .A(_3686_),
    .B(_3681_),
    .Y(_3691_)
);

XNOR2X1 _14470_ (
    .A(_3691_),
    .B(_3536_),
    .Y(\datapath.nextpc [22])
);

NAND2X1 _14471_ (
    .A(_3558__bF$buf2),
    .B(\datapath.nextpc [22]),
    .Y(_3692_)
);

NAND2X1 _14472_ (
    .A(\datapath.programcounter.jumps [22]),
    .B(_3561__bF$buf2),
    .Y(_3693_)
);

NAND2X1 _14473_ (
    .A(\datapath.csr.csr_pcaddr [22]),
    .B(_3563__bF$buf2),
    .Y(_3694_)
);

NAND2X1 _14474_ (
    .A(_0_[22]),
    .B(_3557__bF$buf2),
    .Y(_3695_)
);

AND2X2 _14475_ (
    .A(_3694_),
    .B(_3695_),
    .Y(_3696_)
);

NAND3X1 _14476_ (
    .A(_3693_),
    .B(_3696_),
    .C(_3692_),
    .Y(\datapath.programcounter.pc_mux [22])
);

OAI21X1 _14477_ (
    .A(_3536_),
    .B(_3687_),
    .C(_3538_),
    .Y(_3697_)
);

NAND3X1 _14478_ (
    .A(\datapath.programcounter.pc [22]),
    .B(\datapath.programcounter.pc [23]),
    .C(_3691_),
    .Y(_3698_)
);

AND2X2 _14479_ (
    .A(_3697_),
    .B(_3698_),
    .Y(\datapath.nextpc [23])
);

NAND3X1 _14480_ (
    .A(_3558__bF$buf1),
    .B(_3698_),
    .C(_3697_),
    .Y(_3699_)
);

NAND2X1 _14481_ (
    .A(_0_[23]),
    .B(_3557__bF$buf1),
    .Y(_3700_)
);

AOI22X1 _14482_ (
    .A(_3561__bF$buf1),
    .B(\datapath.programcounter.jumps [23]),
    .C(\datapath.csr.csr_pcaddr [23]),
    .D(_3563__bF$buf1),
    .Y(_3701_)
);

NAND3X1 _14483_ (
    .A(_3700_),
    .B(_3701_),
    .C(_3699_),
    .Y(\datapath.programcounter.pc_mux [23])
);

NAND2X1 _14484_ (
    .A(\datapath.programcounter.pc [22]),
    .B(\datapath.programcounter.pc [23]),
    .Y(_3702_)
);

NOR2X1 _14485_ (
    .A(_3686_),
    .B(_3702_),
    .Y(_3703_)
);

AND2X2 _14486_ (
    .A(_3680_),
    .B(_3703_),
    .Y(_3704_)
);

NAND3X1 _14487_ (
    .A(_3662_),
    .B(_3663_),
    .C(_3704_),
    .Y(_3705_)
);

XNOR2X1 _14488_ (
    .A(_3705_),
    .B(\datapath.programcounter.pc [24]),
    .Y(\datapath.nextpc [24])
);

NAND2X1 _14489_ (
    .A(\datapath.programcounter.jumps [24]),
    .B(_3561__bF$buf0),
    .Y(_3706_)
);

NAND2X1 _14490_ (
    .A(\datapath.csr.csr_pcaddr [24]),
    .B(_3563__bF$buf0),
    .Y(_3707_)
);

AOI22X1 _14491_ (
    .A(_0_[24]),
    .B(_3557__bF$buf0),
    .C(_3558__bF$buf0),
    .D(\datapath.nextpc [24]),
    .Y(_3708_)
);

NAND3X1 _14492_ (
    .A(_3706_),
    .B(_3707_),
    .C(_3708_),
    .Y(\datapath.programcounter.pc_mux [24])
);

OAI21X1 _14493_ (
    .A(_3540_),
    .B(_3705_),
    .C(_3542_),
    .Y(_3709_)
);

NAND2X1 _14494_ (
    .A(_3680_),
    .B(_3703_),
    .Y(_3710_)
);

NOR2X1 _14495_ (
    .A(_3710_),
    .B(_3664_),
    .Y(_3711_)
);

NAND3X1 _14496_ (
    .A(\datapath.programcounter.pc [24]),
    .B(\datapath.programcounter.pc [25]),
    .C(_3711_),
    .Y(_3712_)
);

AND2X2 _14497_ (
    .A(_3712_),
    .B(_3709_),
    .Y(\datapath.nextpc [25])
);

NAND2X1 _14498_ (
    .A(_3558__bF$buf4),
    .B(\datapath.nextpc [25]),
    .Y(_3713_)
);

NAND2X1 _14499_ (
    .A(\datapath.programcounter.jumps [25]),
    .B(_3561__bF$buf4),
    .Y(_3714_)
);

AOI22X1 _14500_ (
    .A(_3557__bF$buf4),
    .B(_0_[25]),
    .C(\datapath.csr.csr_pcaddr [25]),
    .D(_3563__bF$buf4),
    .Y(_3715_)
);

NAND3X1 _14501_ (
    .A(_3714_),
    .B(_3715_),
    .C(_3713_),
    .Y(\datapath.programcounter.pc_mux [25])
);

NAND2X1 _14502_ (
    .A(\datapath.programcounter.pc [24]),
    .B(\datapath.programcounter.pc [25]),
    .Y(_3716_)
);

OAI21X1 _14503_ (
    .A(_3716_),
    .B(_3705_),
    .C(_3544_),
    .Y(_3717_)
);

NOR2X1 _14504_ (
    .A(_3716_),
    .B(_3705_),
    .Y(_3718_)
);

NAND2X1 _14505_ (
    .A(\datapath.programcounter.pc [26]),
    .B(_3718_),
    .Y(_3719_)
);

AND2X2 _14506_ (
    .A(_3719_),
    .B(_3717_),
    .Y(\datapath.nextpc [26])
);

NAND3X1 _14507_ (
    .A(_3558__bF$buf3),
    .B(_3717_),
    .C(_3719_),
    .Y(_3720_)
);

NAND2X1 _14508_ (
    .A(\datapath.programcounter.jumps [26]),
    .B(_3561__bF$buf3),
    .Y(_3721_)
);

AOI22X1 _14509_ (
    .A(_3557__bF$buf3),
    .B(_0_[26]),
    .C(\datapath.csr.csr_pcaddr [26]),
    .D(_3563__bF$buf3),
    .Y(_3722_)
);

NAND3X1 _14510_ (
    .A(_3721_),
    .B(_3722_),
    .C(_3720_),
    .Y(\datapath.programcounter.pc_mux [26])
);

INVX1 _14511_ (
    .A(_3716_),
    .Y(_3723_)
);

NAND2X1 _14512_ (
    .A(_3723_),
    .B(_3711_),
    .Y(_3724_)
);

OAI21X1 _14513_ (
    .A(_3544_),
    .B(_3724_),
    .C(_3546_),
    .Y(_3725_)
);

NAND3X1 _14514_ (
    .A(\datapath.programcounter.pc [26]),
    .B(\datapath.programcounter.pc [27]),
    .C(_3718_),
    .Y(_3726_)
);

AND2X2 _14515_ (
    .A(_3725_),
    .B(_3726_),
    .Y(\datapath.nextpc [27])
);

NAND3X1 _14516_ (
    .A(_3558__bF$buf2),
    .B(_3726_),
    .C(_3725_),
    .Y(_3727_)
);

NAND2X1 _14517_ (
    .A(_0_[27]),
    .B(_3557__bF$buf2),
    .Y(_3728_)
);

AOI22X1 _14518_ (
    .A(_3561__bF$buf2),
    .B(\datapath.programcounter.jumps [27]),
    .C(\datapath.csr.csr_pcaddr [27]),
    .D(_3563__bF$buf2),
    .Y(_3729_)
);

NAND3X1 _14519_ (
    .A(_3728_),
    .B(_3729_),
    .C(_3727_),
    .Y(\datapath.programcounter.pc_mux [27])
);

NAND2X1 _14520_ (
    .A(\datapath.programcounter.pc [26]),
    .B(\datapath.programcounter.pc [27]),
    .Y(_3730_)
);

NOR2X1 _14521_ (
    .A(_3716_),
    .B(_3730_),
    .Y(_3731_)
);

INVX1 _14522_ (
    .A(_3731_),
    .Y(_3732_)
);

NOR3X1 _14523_ (
    .A(_3710_),
    .B(_3732_),
    .C(_3664_),
    .Y(_3733_)
);

XNOR2X1 _14524_ (
    .A(_3733_),
    .B(_3548_),
    .Y(\datapath.nextpc [28])
);

NAND2X1 _14525_ (
    .A(_3558__bF$buf1),
    .B(\datapath.nextpc [28]),
    .Y(_3734_)
);

NAND2X1 _14526_ (
    .A(\datapath.programcounter.jumps [28]),
    .B(_3561__bF$buf1),
    .Y(_3735_)
);

NAND2X1 _14527_ (
    .A(\datapath.csr.csr_pcaddr [28]),
    .B(_3563__bF$buf1),
    .Y(_3736_)
);

NAND2X1 _14528_ (
    .A(_0_[28]),
    .B(_3557__bF$buf1),
    .Y(_3737_)
);

NAND3X1 _14529_ (
    .A(_3735_),
    .B(_3737_),
    .C(_3736_),
    .Y(_3738_)
);

INVX1 _14530_ (
    .A(_3738_),
    .Y(_3739_)
);

NAND2X1 _14531_ (
    .A(_3739_),
    .B(_3734_),
    .Y(\datapath.programcounter.pc_mux [28])
);

NAND2X1 _14532_ (
    .A(_3731_),
    .B(_3711_),
    .Y(_3740_)
);

OAI21X1 _14533_ (
    .A(_3548_),
    .B(_3740_),
    .C(_3550_),
    .Y(_3741_)
);

NAND3X1 _14534_ (
    .A(\datapath.programcounter.pc [28]),
    .B(\datapath.programcounter.pc [29]),
    .C(_3733_),
    .Y(_3742_)
);

AND2X2 _14535_ (
    .A(_3741_),
    .B(_3742_),
    .Y(\datapath.nextpc [29])
);

NAND3X1 _14536_ (
    .A(_3558__bF$buf0),
    .B(_3742_),
    .C(_3741_),
    .Y(_3743_)
);

NAND2X1 _14537_ (
    .A(\datapath.csr.csr_pcaddr [29]),
    .B(_3563__bF$buf0),
    .Y(_3744_)
);

AOI22X1 _14538_ (
    .A(_3557__bF$buf0),
    .B(_0_[29]),
    .C(\datapath.programcounter.jumps [29]),
    .D(_3561__bF$buf0),
    .Y(_3745_)
);

NAND3X1 _14539_ (
    .A(_3744_),
    .B(_3745_),
    .C(_3743_),
    .Y(\datapath.programcounter.pc_mux [29])
);

NAND2X1 _14540_ (
    .A(\datapath.programcounter.pc [28]),
    .B(\datapath.programcounter.pc [29]),
    .Y(_3746_)
);

OAI21X1 _14541_ (
    .A(_3746_),
    .B(_3740_),
    .C(_3552_),
    .Y(_3747_)
);

INVX1 _14542_ (
    .A(_3746_),
    .Y(_3748_)
);

NAND3X1 _14543_ (
    .A(\datapath.programcounter.pc [30]),
    .B(_3748_),
    .C(_3733_),
    .Y(_3749_)
);

AND2X2 _14544_ (
    .A(_3747_),
    .B(_3749_),
    .Y(\datapath.nextpc [30])
);

NAND3X1 _14545_ (
    .A(_3558__bF$buf4),
    .B(_3749_),
    .C(_3747_),
    .Y(_3750_)
);

NAND2X1 _14546_ (
    .A(\datapath.csr.csr_pcaddr [30]),
    .B(_3563__bF$buf4),
    .Y(_3751_)
);

AOI22X1 _14547_ (
    .A(_3557__bF$buf4),
    .B(_0_[30]),
    .C(\datapath.programcounter.jumps [30]),
    .D(_3561__bF$buf4),
    .Y(_3752_)
);

NAND3X1 _14548_ (
    .A(_3751_),
    .B(_3752_),
    .C(_3750_),
    .Y(\datapath.programcounter.pc_mux [30])
);

NAND2X1 _14549_ (
    .A(_3554_),
    .B(_3749_),
    .Y(_3753_)
);

NOR3X1 _14550_ (
    .A(_3732_),
    .B(_3746_),
    .C(_3705_),
    .Y(_3754_)
);

NAND3X1 _14551_ (
    .A(\datapath.programcounter.pc [30]),
    .B(\datapath.programcounter.pc [31]),
    .C(_3754_),
    .Y(_3755_)
);

AND2X2 _14552_ (
    .A(_3753_),
    .B(_3755_),
    .Y(\datapath.nextpc [31])
);

NAND3X1 _14553_ (
    .A(_3558__bF$buf3),
    .B(_3755_),
    .C(_3753_),
    .Y(_3756_)
);

NAND2X1 _14554_ (
    .A(_0_[31]),
    .B(_3557__bF$buf3),
    .Y(_3757_)
);

NAND2X1 _14555_ (
    .A(\datapath.programcounter.jumps [31]),
    .B(_3561__bF$buf3),
    .Y(_3758_)
);

NAND2X1 _14556_ (
    .A(\datapath.csr.csr_pcaddr [31]),
    .B(_3563__bF$buf3),
    .Y(_3759_)
);

NAND3X1 _14557_ (
    .A(_3757_),
    .B(_3758_),
    .C(_3759_),
    .Y(_3760_)
);

INVX1 _14558_ (
    .A(_3760_),
    .Y(_3761_)
);

NAND2X1 _14559_ (
    .A(_3761_),
    .B(_3756_),
    .Y(\datapath.programcounter.pc_mux [31])
);

DFFPOSX1 _14560_ (
    .CLK(CLK_bF$buf79),
    .D(\datapath.programcounter._1_ [0]),
    .Q(\datapath.programcounter.pc [0])
);

DFFPOSX1 _14561_ (
    .CLK(CLK_bF$buf78),
    .D(\datapath.programcounter._1_ [1]),
    .Q(\datapath.programcounter.pc [1])
);

DFFPOSX1 _14562_ (
    .CLK(CLK_bF$buf77),
    .D(\datapath.programcounter._1_ [2]),
    .Q(\datapath.programcounter.pc [2])
);

DFFPOSX1 _14563_ (
    .CLK(CLK_bF$buf76),
    .D(\datapath.programcounter._1_ [3]),
    .Q(\datapath.programcounter.pc [3])
);

DFFPOSX1 _14564_ (
    .CLK(CLK_bF$buf75),
    .D(\datapath.programcounter._1_ [4]),
    .Q(\datapath.programcounter.pc [4])
);

DFFPOSX1 _14565_ (
    .CLK(CLK_bF$buf74),
    .D(\datapath.programcounter._1_ [5]),
    .Q(\datapath.programcounter.pc [5])
);

DFFPOSX1 _14566_ (
    .CLK(CLK_bF$buf73),
    .D(\datapath.programcounter._1_ [6]),
    .Q(\datapath.programcounter.pc [6])
);

DFFPOSX1 _14567_ (
    .CLK(CLK_bF$buf72),
    .D(\datapath.programcounter._1_ [7]),
    .Q(\datapath.programcounter.pc [7])
);

DFFPOSX1 _14568_ (
    .CLK(CLK_bF$buf71),
    .D(\datapath.programcounter._1_ [8]),
    .Q(\datapath.programcounter.pc [8])
);

DFFPOSX1 _14569_ (
    .CLK(CLK_bF$buf70),
    .D(\datapath.programcounter._1_ [9]),
    .Q(\datapath.programcounter.pc [9])
);

DFFPOSX1 _14570_ (
    .CLK(CLK_bF$buf69),
    .D(\datapath.programcounter._1_ [10]),
    .Q(\datapath.programcounter.pc [10])
);

DFFPOSX1 _14571_ (
    .CLK(CLK_bF$buf68),
    .D(\datapath.programcounter._1_ [11]),
    .Q(\datapath.programcounter.pc [11])
);

DFFPOSX1 _14572_ (
    .CLK(CLK_bF$buf67),
    .D(\datapath.programcounter._1_ [12]),
    .Q(\datapath.programcounter.pc [12])
);

DFFPOSX1 _14573_ (
    .CLK(CLK_bF$buf66),
    .D(\datapath.programcounter._1_ [13]),
    .Q(\datapath.programcounter.pc [13])
);

DFFPOSX1 _14574_ (
    .CLK(CLK_bF$buf65),
    .D(\datapath.programcounter._1_ [14]),
    .Q(\datapath.programcounter.pc [14])
);

DFFPOSX1 _14575_ (
    .CLK(CLK_bF$buf64),
    .D(\datapath.programcounter._1_ [15]),
    .Q(\datapath.programcounter.pc [15])
);

DFFPOSX1 _14576_ (
    .CLK(CLK_bF$buf63),
    .D(\datapath.programcounter._1_ [16]),
    .Q(\datapath.programcounter.pc [16])
);

DFFPOSX1 _14577_ (
    .CLK(CLK_bF$buf62),
    .D(\datapath.programcounter._1_ [17]),
    .Q(\datapath.programcounter.pc [17])
);

DFFPOSX1 _14578_ (
    .CLK(CLK_bF$buf61),
    .D(\datapath.programcounter._1_ [18]),
    .Q(\datapath.programcounter.pc [18])
);

DFFPOSX1 _14579_ (
    .CLK(CLK_bF$buf60),
    .D(\datapath.programcounter._1_ [19]),
    .Q(\datapath.programcounter.pc [19])
);

DFFPOSX1 _14580_ (
    .CLK(CLK_bF$buf59),
    .D(\datapath.programcounter._1_ [20]),
    .Q(\datapath.programcounter.pc [20])
);

DFFPOSX1 _14581_ (
    .CLK(CLK_bF$buf58),
    .D(\datapath.programcounter._1_ [21]),
    .Q(\datapath.programcounter.pc [21])
);

DFFPOSX1 _14582_ (
    .CLK(CLK_bF$buf57),
    .D(\datapath.programcounter._1_ [22]),
    .Q(\datapath.programcounter.pc [22])
);

DFFPOSX1 _14583_ (
    .CLK(CLK_bF$buf56),
    .D(\datapath.programcounter._1_ [23]),
    .Q(\datapath.programcounter.pc [23])
);

DFFPOSX1 _14584_ (
    .CLK(CLK_bF$buf55),
    .D(\datapath.programcounter._1_ [24]),
    .Q(\datapath.programcounter.pc [24])
);

DFFPOSX1 _14585_ (
    .CLK(CLK_bF$buf54),
    .D(\datapath.programcounter._1_ [25]),
    .Q(\datapath.programcounter.pc [25])
);

DFFPOSX1 _14586_ (
    .CLK(CLK_bF$buf53),
    .D(\datapath.programcounter._1_ [26]),
    .Q(\datapath.programcounter.pc [26])
);

DFFPOSX1 _14587_ (
    .CLK(CLK_bF$buf52),
    .D(\datapath.programcounter._1_ [27]),
    .Q(\datapath.programcounter.pc [27])
);

DFFPOSX1 _14588_ (
    .CLK(CLK_bF$buf51),
    .D(\datapath.programcounter._1_ [28]),
    .Q(\datapath.programcounter.pc [28])
);

DFFPOSX1 _14589_ (
    .CLK(CLK_bF$buf50),
    .D(\datapath.programcounter._1_ [29]),
    .Q(\datapath.programcounter.pc [29])
);

DFFPOSX1 _14590_ (
    .CLK(CLK_bF$buf49),
    .D(\datapath.programcounter._1_ [30]),
    .Q(\datapath.programcounter.pc [30])
);

DFFPOSX1 _14591_ (
    .CLK(CLK_bF$buf48),
    .D(\datapath.programcounter._1_ [31]),
    .Q(\datapath.programcounter.pc [31])
);

INVX8 _14592_ (
    .A(\datapath.rd [0]),
    .Y(_4786_)
);

INVX1 _14593_ (
    .A(\datapath.wbinstr [7]),
    .Y(_4787_)
);

NOR2X1 _14594_ (
    .A(\datapath.wbinstr [8]),
    .B(_4787_),
    .Y(_4788_)
);

NOR2X1 _14595_ (
    .A(\datapath.wbinstr [8]),
    .B(\datapath.wbinstr [7]),
    .Y(_4789_)
);

INVX2 _14596_ (
    .A(_4789_),
    .Y(_4790_)
);

INVX1 _14597_ (
    .A(\datapath.wbinstr [9]),
    .Y(_4791_)
);

INVX1 _14598_ (
    .A(\datapath.wbinstr [10]),
    .Y(_4792_)
);

INVX1 _14599_ (
    .A(\datapath.wbinstr [11]),
    .Y(_4793_)
);

NAND3X1 _14600_ (
    .A(_4791_),
    .B(_4792_),
    .C(_4793_),
    .Y(_4794_)
);

OAI21X1 _14601_ (
    .A(_4790_),
    .B(_4794__bF$buf7),
    .C(\controlunit.regfile_wen ),
    .Y(_4795_)
);

NOR2X1 _14602_ (
    .A(\datapath.wbinstr [10]),
    .B(_4793_),
    .Y(_4796_)
);

NAND2X1 _14603_ (
    .A(\datapath.wbinstr [9]),
    .B(_4796_),
    .Y(_4797_)
);

NOR2X1 _14604_ (
    .A(_4797_),
    .B(_4795_),
    .Y(_4798_)
);

NAND2X1 _14605_ (
    .A(_4788_),
    .B(_4798_),
    .Y(_4799_)
);

NAND2X1 _14606_ (
    .A(\datapath.registers.838[21] [0]),
    .B(_4799__bF$buf7),
    .Y(_4800_)
);

OAI21X1 _14607_ (
    .A(_4786__bF$buf4),
    .B(_4799__bF$buf6),
    .C(_4800_),
    .Y(_4178_)
);

INVX8 _14608_ (
    .A(\datapath.rd [1]),
    .Y(_4801_)
);

NAND2X1 _14609_ (
    .A(\datapath.registers.838[21] [1]),
    .B(_4799__bF$buf5),
    .Y(_4802_)
);

OAI21X1 _14610_ (
    .A(_4801__bF$buf4),
    .B(_4799__bF$buf4),
    .C(_4802_),
    .Y(_4189_)
);

INVX8 _14611_ (
    .A(\datapath.rd [2]),
    .Y(_4803_)
);

NAND2X1 _14612_ (
    .A(\datapath.registers.838[21] [2]),
    .B(_4799__bF$buf3),
    .Y(_4804_)
);

OAI21X1 _14613_ (
    .A(_4803__bF$buf4),
    .B(_4799__bF$buf2),
    .C(_4804_),
    .Y(_4200_)
);

INVX8 _14614_ (
    .A(\datapath.rd [3]),
    .Y(_4805_)
);

NAND2X1 _14615_ (
    .A(\datapath.registers.838[21] [3]),
    .B(_4799__bF$buf1),
    .Y(_4806_)
);

OAI21X1 _14616_ (
    .A(_4805__bF$buf4),
    .B(_4799__bF$buf0),
    .C(_4806_),
    .Y(_4203_)
);

INVX8 _14617_ (
    .A(\datapath.rd [4]),
    .Y(_4807_)
);

NAND2X1 _14618_ (
    .A(\datapath.registers.838[21] [4]),
    .B(_4799__bF$buf7),
    .Y(_4808_)
);

OAI21X1 _14619_ (
    .A(_4807__bF$buf4),
    .B(_4799__bF$buf6),
    .C(_4808_),
    .Y(_4204_)
);

INVX8 _14620_ (
    .A(\datapath.rd [5]),
    .Y(_4809_)
);

NAND2X1 _14621_ (
    .A(\datapath.registers.838[21] [5]),
    .B(_4799__bF$buf5),
    .Y(_4810_)
);

OAI21X1 _14622_ (
    .A(_4809__bF$buf4),
    .B(_4799__bF$buf4),
    .C(_4810_),
    .Y(_4205_)
);

INVX8 _14623_ (
    .A(\datapath.rd [6]),
    .Y(_4811_)
);

NAND2X1 _14624_ (
    .A(\datapath.registers.838[21] [6]),
    .B(_4799__bF$buf3),
    .Y(_4812_)
);

OAI21X1 _14625_ (
    .A(_4811__bF$buf4),
    .B(_4799__bF$buf2),
    .C(_4812_),
    .Y(_4206_)
);

INVX8 _14626_ (
    .A(\datapath.rd [7]),
    .Y(_4813_)
);

NAND2X1 _14627_ (
    .A(\datapath.registers.838[21] [7]),
    .B(_4799__bF$buf1),
    .Y(_4814_)
);

OAI21X1 _14628_ (
    .A(_4813__bF$buf4),
    .B(_4799__bF$buf0),
    .C(_4814_),
    .Y(_4207_)
);

INVX8 _14629_ (
    .A(\datapath.rd [8]),
    .Y(_4815_)
);

NAND2X1 _14630_ (
    .A(\datapath.registers.838[21] [8]),
    .B(_4799__bF$buf7),
    .Y(_4816_)
);

OAI21X1 _14631_ (
    .A(_4815__bF$buf4),
    .B(_4799__bF$buf6),
    .C(_4816_),
    .Y(_4208_)
);

INVX8 _14632_ (
    .A(\datapath.rd [9]),
    .Y(_4817_)
);

NAND2X1 _14633_ (
    .A(\datapath.registers.838[21] [9]),
    .B(_4799__bF$buf5),
    .Y(_4818_)
);

OAI21X1 _14634_ (
    .A(_4817__bF$buf4),
    .B(_4799__bF$buf4),
    .C(_4818_),
    .Y(_4209_)
);

INVX8 _14635_ (
    .A(\datapath.rd [10]),
    .Y(_4819_)
);

NAND2X1 _14636_ (
    .A(\datapath.registers.838[21] [10]),
    .B(_4799__bF$buf3),
    .Y(_4820_)
);

OAI21X1 _14637_ (
    .A(_4819__bF$buf4),
    .B(_4799__bF$buf2),
    .C(_4820_),
    .Y(_4179_)
);

INVX8 _14638_ (
    .A(\datapath.rd [11]),
    .Y(_4821_)
);

NAND2X1 _14639_ (
    .A(\datapath.registers.838[21] [11]),
    .B(_4799__bF$buf1),
    .Y(_4822_)
);

OAI21X1 _14640_ (
    .A(_4821__bF$buf4),
    .B(_4799__bF$buf0),
    .C(_4822_),
    .Y(_4180_)
);

INVX8 _14641_ (
    .A(\datapath.rd [12]),
    .Y(_4823_)
);

NAND2X1 _14642_ (
    .A(\datapath.registers.838[21] [12]),
    .B(_4799__bF$buf7),
    .Y(_4824_)
);

OAI21X1 _14643_ (
    .A(_4823__bF$buf4),
    .B(_4799__bF$buf6),
    .C(_4824_),
    .Y(_4181_)
);

INVX8 _14644_ (
    .A(\datapath.rd [13]),
    .Y(_4825_)
);

NAND2X1 _14645_ (
    .A(\datapath.registers.838[21] [13]),
    .B(_4799__bF$buf5),
    .Y(_4826_)
);

OAI21X1 _14646_ (
    .A(_4825__bF$buf4),
    .B(_4799__bF$buf4),
    .C(_4826_),
    .Y(_4182_)
);

INVX8 _14647_ (
    .A(\datapath.rd [14]),
    .Y(_4827_)
);

NAND2X1 _14648_ (
    .A(\datapath.registers.838[21] [14]),
    .B(_4799__bF$buf3),
    .Y(_4828_)
);

OAI21X1 _14649_ (
    .A(_4827__bF$buf4),
    .B(_4799__bF$buf2),
    .C(_4828_),
    .Y(_4183_)
);

INVX8 _14650_ (
    .A(\datapath.rd [15]),
    .Y(_4829_)
);

NAND2X1 _14651_ (
    .A(\datapath.registers.838[21] [15]),
    .B(_4799__bF$buf1),
    .Y(_4830_)
);

OAI21X1 _14652_ (
    .A(_4829__bF$buf4),
    .B(_4799__bF$buf0),
    .C(_4830_),
    .Y(_4184_)
);

INVX8 _14653_ (
    .A(\datapath.rd [16]),
    .Y(_4831_)
);

NAND2X1 _14654_ (
    .A(\datapath.registers.838[21] [16]),
    .B(_4799__bF$buf7),
    .Y(_4832_)
);

OAI21X1 _14655_ (
    .A(_4831__bF$buf4),
    .B(_4799__bF$buf6),
    .C(_4832_),
    .Y(_4185_)
);

INVX8 _14656_ (
    .A(\datapath.rd [17]),
    .Y(_4833_)
);

NAND2X1 _14657_ (
    .A(\datapath.registers.838[21] [17]),
    .B(_4799__bF$buf5),
    .Y(_4834_)
);

OAI21X1 _14658_ (
    .A(_4833__bF$buf4),
    .B(_4799__bF$buf4),
    .C(_4834_),
    .Y(_4186_)
);

INVX8 _14659_ (
    .A(\datapath.rd [18]),
    .Y(_4835_)
);

NAND2X1 _14660_ (
    .A(\datapath.registers.838[21] [18]),
    .B(_4799__bF$buf3),
    .Y(_4836_)
);

OAI21X1 _14661_ (
    .A(_4835__bF$buf4),
    .B(_4799__bF$buf2),
    .C(_4836_),
    .Y(_4187_)
);

INVX8 _14662_ (
    .A(\datapath.rd [19]),
    .Y(_4837_)
);

NAND2X1 _14663_ (
    .A(\datapath.registers.838[21] [19]),
    .B(_4799__bF$buf1),
    .Y(_4838_)
);

OAI21X1 _14664_ (
    .A(_4837__bF$buf4),
    .B(_4799__bF$buf0),
    .C(_4838_),
    .Y(_4188_)
);

INVX8 _14665_ (
    .A(\datapath.rd [20]),
    .Y(_4839_)
);

NAND2X1 _14666_ (
    .A(\datapath.registers.838[21] [20]),
    .B(_4799__bF$buf7),
    .Y(_4840_)
);

OAI21X1 _14667_ (
    .A(_4839__bF$buf4),
    .B(_4799__bF$buf6),
    .C(_4840_),
    .Y(_4190_)
);

INVX8 _14668_ (
    .A(\datapath.rd [21]),
    .Y(_4841_)
);

NAND2X1 _14669_ (
    .A(\datapath.registers.838[21] [21]),
    .B(_4799__bF$buf5),
    .Y(_4842_)
);

OAI21X1 _14670_ (
    .A(_4841__bF$buf4),
    .B(_4799__bF$buf4),
    .C(_4842_),
    .Y(_4191_)
);

INVX8 _14671_ (
    .A(\datapath.rd [22]),
    .Y(_4843_)
);

NAND2X1 _14672_ (
    .A(\datapath.registers.838[21] [22]),
    .B(_4799__bF$buf3),
    .Y(_4844_)
);

OAI21X1 _14673_ (
    .A(_4843__bF$buf4),
    .B(_4799__bF$buf2),
    .C(_4844_),
    .Y(_4192_)
);

INVX8 _14674_ (
    .A(\datapath.rd [23]),
    .Y(_4845_)
);

NAND2X1 _14675_ (
    .A(\datapath.registers.838[21] [23]),
    .B(_4799__bF$buf1),
    .Y(_4846_)
);

OAI21X1 _14676_ (
    .A(_4845__bF$buf4),
    .B(_4799__bF$buf0),
    .C(_4846_),
    .Y(_4193_)
);

INVX8 _14677_ (
    .A(\datapath.rd [24]),
    .Y(_4847_)
);

NAND2X1 _14678_ (
    .A(\datapath.registers.838[21] [24]),
    .B(_4799__bF$buf7),
    .Y(_4848_)
);

OAI21X1 _14679_ (
    .A(_4847__bF$buf4),
    .B(_4799__bF$buf6),
    .C(_4848_),
    .Y(_4194_)
);

INVX8 _14680_ (
    .A(\datapath.rd [25]),
    .Y(_4849_)
);

NAND2X1 _14681_ (
    .A(\datapath.registers.838[21] [25]),
    .B(_4799__bF$buf5),
    .Y(_4850_)
);

OAI21X1 _14682_ (
    .A(_4849__bF$buf4),
    .B(_4799__bF$buf4),
    .C(_4850_),
    .Y(_4195_)
);

INVX8 _14683_ (
    .A(\datapath.rd [26]),
    .Y(_4851_)
);

NAND2X1 _14684_ (
    .A(\datapath.registers.838[21] [26]),
    .B(_4799__bF$buf3),
    .Y(_4852_)
);

OAI21X1 _14685_ (
    .A(_4851__bF$buf4),
    .B(_4799__bF$buf2),
    .C(_4852_),
    .Y(_4196_)
);

INVX8 _14686_ (
    .A(\datapath.rd [27]),
    .Y(_4853_)
);

NAND2X1 _14687_ (
    .A(\datapath.registers.838[21] [27]),
    .B(_4799__bF$buf1),
    .Y(_4854_)
);

OAI21X1 _14688_ (
    .A(_4853__bF$buf4),
    .B(_4799__bF$buf0),
    .C(_4854_),
    .Y(_4197_)
);

INVX8 _14689_ (
    .A(\datapath.rd [28]),
    .Y(_4855_)
);

NAND2X1 _14690_ (
    .A(\datapath.registers.838[21] [28]),
    .B(_4799__bF$buf7),
    .Y(_4856_)
);

OAI21X1 _14691_ (
    .A(_4855__bF$buf4),
    .B(_4799__bF$buf6),
    .C(_4856_),
    .Y(_4198_)
);

INVX8 _14692_ (
    .A(\datapath.rd [29]),
    .Y(_4857_)
);

NAND2X1 _14693_ (
    .A(\datapath.registers.838[21] [29]),
    .B(_4799__bF$buf5),
    .Y(_4858_)
);

OAI21X1 _14694_ (
    .A(_4857__bF$buf4),
    .B(_4799__bF$buf4),
    .C(_4858_),
    .Y(_4199_)
);

INVX8 _14695_ (
    .A(\datapath.rd [30]),
    .Y(_4859_)
);

NAND2X1 _14696_ (
    .A(\datapath.registers.838[21] [30]),
    .B(_4799__bF$buf3),
    .Y(_4860_)
);

OAI21X1 _14697_ (
    .A(_4859__bF$buf4),
    .B(_4799__bF$buf2),
    .C(_4860_),
    .Y(_4201_)
);

INVX8 _14698_ (
    .A(\datapath.rd [31]),
    .Y(_4861_)
);

NAND2X1 _14699_ (
    .A(\datapath.registers.838[21] [31]),
    .B(_4799__bF$buf1),
    .Y(_4862_)
);

OAI21X1 _14700_ (
    .A(_4861__bF$buf4),
    .B(_4799__bF$buf0),
    .C(_4862_),
    .Y(_4202_)
);

NAND2X1 _14701_ (
    .A(_4789_),
    .B(_4798_),
    .Y(_4863_)
);

NAND2X1 _14702_ (
    .A(\datapath.registers.838[20] [0]),
    .B(_4863__bF$buf7),
    .Y(_4864_)
);

OAI21X1 _14703_ (
    .A(_4786__bF$buf3),
    .B(_4863__bF$buf6),
    .C(_4864_),
    .Y(_4146_)
);

NAND2X1 _14704_ (
    .A(\datapath.registers.838[20] [1]),
    .B(_4863__bF$buf5),
    .Y(_4865_)
);

OAI21X1 _14705_ (
    .A(_4801__bF$buf3),
    .B(_4863__bF$buf4),
    .C(_4865_),
    .Y(_4157_)
);

NAND2X1 _14706_ (
    .A(\datapath.registers.838[20] [2]),
    .B(_4863__bF$buf3),
    .Y(_4866_)
);

OAI21X1 _14707_ (
    .A(_4803__bF$buf3),
    .B(_4863__bF$buf2),
    .C(_4866_),
    .Y(_4168_)
);

NAND2X1 _14708_ (
    .A(\datapath.registers.838[20] [3]),
    .B(_4863__bF$buf1),
    .Y(_4867_)
);

OAI21X1 _14709_ (
    .A(_4805__bF$buf3),
    .B(_4863__bF$buf0),
    .C(_4867_),
    .Y(_4171_)
);

NAND2X1 _14710_ (
    .A(\datapath.registers.838[20] [4]),
    .B(_4863__bF$buf7),
    .Y(_4868_)
);

OAI21X1 _14711_ (
    .A(_4807__bF$buf3),
    .B(_4863__bF$buf6),
    .C(_4868_),
    .Y(_4172_)
);

NAND2X1 _14712_ (
    .A(\datapath.registers.838[20] [5]),
    .B(_4863__bF$buf5),
    .Y(_4869_)
);

OAI21X1 _14713_ (
    .A(_4809__bF$buf3),
    .B(_4863__bF$buf4),
    .C(_4869_),
    .Y(_4173_)
);

NAND2X1 _14714_ (
    .A(\datapath.registers.838[20] [6]),
    .B(_4863__bF$buf3),
    .Y(_4870_)
);

OAI21X1 _14715_ (
    .A(_4811__bF$buf3),
    .B(_4863__bF$buf2),
    .C(_4870_),
    .Y(_4174_)
);

NAND2X1 _14716_ (
    .A(\datapath.registers.838[20] [7]),
    .B(_4863__bF$buf1),
    .Y(_4871_)
);

OAI21X1 _14717_ (
    .A(_4813__bF$buf3),
    .B(_4863__bF$buf0),
    .C(_4871_),
    .Y(_4175_)
);

NAND2X1 _14718_ (
    .A(\datapath.registers.838[20] [8]),
    .B(_4863__bF$buf7),
    .Y(_4872_)
);

OAI21X1 _14719_ (
    .A(_4815__bF$buf3),
    .B(_4863__bF$buf6),
    .C(_4872_),
    .Y(_4176_)
);

NAND2X1 _14720_ (
    .A(\datapath.registers.838[20] [9]),
    .B(_4863__bF$buf5),
    .Y(_4873_)
);

OAI21X1 _14721_ (
    .A(_4817__bF$buf3),
    .B(_4863__bF$buf4),
    .C(_4873_),
    .Y(_4177_)
);

NAND2X1 _14722_ (
    .A(\datapath.registers.838[20] [10]),
    .B(_4863__bF$buf3),
    .Y(_4874_)
);

OAI21X1 _14723_ (
    .A(_4819__bF$buf3),
    .B(_4863__bF$buf2),
    .C(_4874_),
    .Y(_4147_)
);

NAND2X1 _14724_ (
    .A(\datapath.registers.838[20] [11]),
    .B(_4863__bF$buf1),
    .Y(_4875_)
);

OAI21X1 _14725_ (
    .A(_4821__bF$buf3),
    .B(_4863__bF$buf0),
    .C(_4875_),
    .Y(_4148_)
);

NAND2X1 _14726_ (
    .A(\datapath.registers.838[20] [12]),
    .B(_4863__bF$buf7),
    .Y(_4876_)
);

OAI21X1 _14727_ (
    .A(_4823__bF$buf3),
    .B(_4863__bF$buf6),
    .C(_4876_),
    .Y(_4149_)
);

NAND2X1 _14728_ (
    .A(\datapath.registers.838[20] [13]),
    .B(_4863__bF$buf5),
    .Y(_4877_)
);

OAI21X1 _14729_ (
    .A(_4825__bF$buf3),
    .B(_4863__bF$buf4),
    .C(_4877_),
    .Y(_4150_)
);

NAND2X1 _14730_ (
    .A(\datapath.registers.838[20] [14]),
    .B(_4863__bF$buf3),
    .Y(_4878_)
);

OAI21X1 _14731_ (
    .A(_4827__bF$buf3),
    .B(_4863__bF$buf2),
    .C(_4878_),
    .Y(_4151_)
);

NAND2X1 _14732_ (
    .A(\datapath.registers.838[20] [15]),
    .B(_4863__bF$buf1),
    .Y(_4879_)
);

OAI21X1 _14733_ (
    .A(_4829__bF$buf3),
    .B(_4863__bF$buf0),
    .C(_4879_),
    .Y(_4152_)
);

NAND2X1 _14734_ (
    .A(\datapath.registers.838[20] [16]),
    .B(_4863__bF$buf7),
    .Y(_4880_)
);

OAI21X1 _14735_ (
    .A(_4831__bF$buf3),
    .B(_4863__bF$buf6),
    .C(_4880_),
    .Y(_4153_)
);

NAND2X1 _14736_ (
    .A(\datapath.registers.838[20] [17]),
    .B(_4863__bF$buf5),
    .Y(_4881_)
);

OAI21X1 _14737_ (
    .A(_4833__bF$buf3),
    .B(_4863__bF$buf4),
    .C(_4881_),
    .Y(_4154_)
);

NAND2X1 _14738_ (
    .A(\datapath.registers.838[20] [18]),
    .B(_4863__bF$buf3),
    .Y(_4882_)
);

OAI21X1 _14739_ (
    .A(_4835__bF$buf3),
    .B(_4863__bF$buf2),
    .C(_4882_),
    .Y(_4155_)
);

NAND2X1 _14740_ (
    .A(\datapath.registers.838[20] [19]),
    .B(_4863__bF$buf1),
    .Y(_4883_)
);

OAI21X1 _14741_ (
    .A(_4837__bF$buf3),
    .B(_4863__bF$buf0),
    .C(_4883_),
    .Y(_4156_)
);

NAND2X1 _14742_ (
    .A(\datapath.registers.838[20] [20]),
    .B(_4863__bF$buf7),
    .Y(_4884_)
);

OAI21X1 _14743_ (
    .A(_4839__bF$buf3),
    .B(_4863__bF$buf6),
    .C(_4884_),
    .Y(_4158_)
);

NAND2X1 _14744_ (
    .A(\datapath.registers.838[20] [21]),
    .B(_4863__bF$buf5),
    .Y(_4885_)
);

OAI21X1 _14745_ (
    .A(_4841__bF$buf3),
    .B(_4863__bF$buf4),
    .C(_4885_),
    .Y(_4159_)
);

NAND2X1 _14746_ (
    .A(\datapath.registers.838[20] [22]),
    .B(_4863__bF$buf3),
    .Y(_4886_)
);

OAI21X1 _14747_ (
    .A(_4843__bF$buf3),
    .B(_4863__bF$buf2),
    .C(_4886_),
    .Y(_4160_)
);

NAND2X1 _14748_ (
    .A(\datapath.registers.838[20] [23]),
    .B(_4863__bF$buf1),
    .Y(_4887_)
);

OAI21X1 _14749_ (
    .A(_4845__bF$buf3),
    .B(_4863__bF$buf0),
    .C(_4887_),
    .Y(_4161_)
);

NAND2X1 _14750_ (
    .A(\datapath.registers.838[20] [24]),
    .B(_4863__bF$buf7),
    .Y(_4888_)
);

OAI21X1 _14751_ (
    .A(_4847__bF$buf3),
    .B(_4863__bF$buf6),
    .C(_4888_),
    .Y(_4162_)
);

NAND2X1 _14752_ (
    .A(\datapath.registers.838[20] [25]),
    .B(_4863__bF$buf5),
    .Y(_4889_)
);

OAI21X1 _14753_ (
    .A(_4849__bF$buf3),
    .B(_4863__bF$buf4),
    .C(_4889_),
    .Y(_4163_)
);

NAND2X1 _14754_ (
    .A(\datapath.registers.838[20] [26]),
    .B(_4863__bF$buf3),
    .Y(_4890_)
);

OAI21X1 _14755_ (
    .A(_4851__bF$buf3),
    .B(_4863__bF$buf2),
    .C(_4890_),
    .Y(_4164_)
);

NAND2X1 _14756_ (
    .A(\datapath.registers.838[20] [27]),
    .B(_4863__bF$buf1),
    .Y(_4891_)
);

OAI21X1 _14757_ (
    .A(_4853__bF$buf3),
    .B(_4863__bF$buf0),
    .C(_4891_),
    .Y(_4165_)
);

NAND2X1 _14758_ (
    .A(\datapath.registers.838[20] [28]),
    .B(_4863__bF$buf7),
    .Y(_4892_)
);

OAI21X1 _14759_ (
    .A(_4855__bF$buf3),
    .B(_4863__bF$buf6),
    .C(_4892_),
    .Y(_4166_)
);

NAND2X1 _14760_ (
    .A(\datapath.registers.838[20] [29]),
    .B(_4863__bF$buf5),
    .Y(_4893_)
);

OAI21X1 _14761_ (
    .A(_4857__bF$buf3),
    .B(_4863__bF$buf4),
    .C(_4893_),
    .Y(_4167_)
);

NAND2X1 _14762_ (
    .A(\datapath.registers.838[20] [30]),
    .B(_4863__bF$buf3),
    .Y(_4894_)
);

OAI21X1 _14763_ (
    .A(_4859__bF$buf3),
    .B(_4863__bF$buf2),
    .C(_4894_),
    .Y(_4169_)
);

NAND2X1 _14764_ (
    .A(\datapath.registers.838[20] [31]),
    .B(_4863__bF$buf1),
    .Y(_4895_)
);

OAI21X1 _14765_ (
    .A(_4861__bF$buf3),
    .B(_4863__bF$buf0),
    .C(_4895_),
    .Y(_4170_)
);

NAND2X1 _14766_ (
    .A(_4791_),
    .B(_4796_),
    .Y(_4896_)
);

INVX1 _14767_ (
    .A(\datapath.wbinstr [8]),
    .Y(_4897_)
);

NOR2X1 _14768_ (
    .A(_4897_),
    .B(_4787_),
    .Y(_4898_)
);

NAND2X1 _14769_ (
    .A(\controlunit.regfile_wen ),
    .B(_4898_),
    .Y(_4899_)
);

OR2X2 _14770_ (
    .A(_4899__bF$buf13),
    .B(_4896__bF$buf5),
    .Y(_4900_)
);

OAI21X1 _14771_ (
    .A(_4896__bF$buf4),
    .B(_4899__bF$buf12),
    .C(\datapath.registers.838[19] [0]),
    .Y(_4901_)
);

OAI21X1 _14772_ (
    .A(_4786__bF$buf2),
    .B(_4900__bF$buf4),
    .C(_4901_),
    .Y(_4082_)
);

OAI21X1 _14773_ (
    .A(_4896__bF$buf3),
    .B(_4899__bF$buf11),
    .C(\datapath.registers.838[19] [1]),
    .Y(_4902_)
);

OAI21X1 _14774_ (
    .A(_4801__bF$buf2),
    .B(_4900__bF$buf3),
    .C(_4902_),
    .Y(_4093_)
);

OAI21X1 _14775_ (
    .A(_4896__bF$buf2),
    .B(_4899__bF$buf10),
    .C(\datapath.registers.838[19] [2]),
    .Y(_4903_)
);

OAI21X1 _14776_ (
    .A(_4803__bF$buf2),
    .B(_4900__bF$buf2),
    .C(_4903_),
    .Y(_4104_)
);

OAI21X1 _14777_ (
    .A(_4896__bF$buf1),
    .B(_4899__bF$buf9),
    .C(\datapath.registers.838[19] [3]),
    .Y(_4904_)
);

OAI21X1 _14778_ (
    .A(_4805__bF$buf2),
    .B(_4900__bF$buf1),
    .C(_4904_),
    .Y(_4107_)
);

OAI21X1 _14779_ (
    .A(_4896__bF$buf0),
    .B(_4899__bF$buf8),
    .C(\datapath.registers.838[19] [4]),
    .Y(_4905_)
);

OAI21X1 _14780_ (
    .A(_4807__bF$buf2),
    .B(_4900__bF$buf0),
    .C(_4905_),
    .Y(_4108_)
);

OAI21X1 _14781_ (
    .A(_4896__bF$buf5),
    .B(_4899__bF$buf7),
    .C(\datapath.registers.838[19] [5]),
    .Y(_4906_)
);

OAI21X1 _14782_ (
    .A(_4809__bF$buf2),
    .B(_4900__bF$buf4),
    .C(_4906_),
    .Y(_4109_)
);

OAI21X1 _14783_ (
    .A(_4896__bF$buf4),
    .B(_4899__bF$buf6),
    .C(\datapath.registers.838[19] [6]),
    .Y(_4907_)
);

OAI21X1 _14784_ (
    .A(_4811__bF$buf2),
    .B(_4900__bF$buf3),
    .C(_4907_),
    .Y(_4110_)
);

OAI21X1 _14785_ (
    .A(_4896__bF$buf3),
    .B(_4899__bF$buf5),
    .C(\datapath.registers.838[19] [7]),
    .Y(_4908_)
);

OAI21X1 _14786_ (
    .A(_4813__bF$buf2),
    .B(_4900__bF$buf2),
    .C(_4908_),
    .Y(_4111_)
);

OAI21X1 _14787_ (
    .A(_4896__bF$buf2),
    .B(_4899__bF$buf4),
    .C(\datapath.registers.838[19] [8]),
    .Y(_4909_)
);

OAI21X1 _14788_ (
    .A(_4815__bF$buf2),
    .B(_4900__bF$buf1),
    .C(_4909_),
    .Y(_4112_)
);

OAI21X1 _14789_ (
    .A(_4896__bF$buf1),
    .B(_4899__bF$buf3),
    .C(\datapath.registers.838[19] [9]),
    .Y(_4910_)
);

OAI21X1 _14790_ (
    .A(_4817__bF$buf2),
    .B(_4900__bF$buf0),
    .C(_4910_),
    .Y(_4113_)
);

OAI21X1 _14791_ (
    .A(_4896__bF$buf0),
    .B(_4899__bF$buf2),
    .C(\datapath.registers.838[19] [10]),
    .Y(_4911_)
);

OAI21X1 _14792_ (
    .A(_4819__bF$buf2),
    .B(_4900__bF$buf4),
    .C(_4911_),
    .Y(_4083_)
);

OAI21X1 _14793_ (
    .A(_4896__bF$buf5),
    .B(_4899__bF$buf1),
    .C(\datapath.registers.838[19] [11]),
    .Y(_4912_)
);

OAI21X1 _14794_ (
    .A(_4821__bF$buf2),
    .B(_4900__bF$buf3),
    .C(_4912_),
    .Y(_4084_)
);

OAI21X1 _14795_ (
    .A(_4896__bF$buf4),
    .B(_4899__bF$buf0),
    .C(\datapath.registers.838[19] [12]),
    .Y(_4913_)
);

OAI21X1 _14796_ (
    .A(_4823__bF$buf2),
    .B(_4900__bF$buf2),
    .C(_4913_),
    .Y(_4085_)
);

OAI21X1 _14797_ (
    .A(_4896__bF$buf3),
    .B(_4899__bF$buf13),
    .C(\datapath.registers.838[19] [13]),
    .Y(_4914_)
);

OAI21X1 _14798_ (
    .A(_4825__bF$buf2),
    .B(_4900__bF$buf1),
    .C(_4914_),
    .Y(_4086_)
);

OAI21X1 _14799_ (
    .A(_4896__bF$buf2),
    .B(_4899__bF$buf12),
    .C(\datapath.registers.838[19] [14]),
    .Y(_4915_)
);

OAI21X1 _14800_ (
    .A(_4827__bF$buf2),
    .B(_4900__bF$buf0),
    .C(_4915_),
    .Y(_4087_)
);

OAI21X1 _14801_ (
    .A(_4896__bF$buf1),
    .B(_4899__bF$buf11),
    .C(\datapath.registers.838[19] [15]),
    .Y(_4916_)
);

OAI21X1 _14802_ (
    .A(_4829__bF$buf2),
    .B(_4900__bF$buf4),
    .C(_4916_),
    .Y(_4088_)
);

OAI21X1 _14803_ (
    .A(_4896__bF$buf0),
    .B(_4899__bF$buf10),
    .C(\datapath.registers.838[19] [16]),
    .Y(_4917_)
);

OAI21X1 _14804_ (
    .A(_4831__bF$buf2),
    .B(_4900__bF$buf3),
    .C(_4917_),
    .Y(_4089_)
);

OAI21X1 _14805_ (
    .A(_4896__bF$buf5),
    .B(_4899__bF$buf9),
    .C(\datapath.registers.838[19] [17]),
    .Y(_4918_)
);

OAI21X1 _14806_ (
    .A(_4833__bF$buf2),
    .B(_4900__bF$buf2),
    .C(_4918_),
    .Y(_4090_)
);

OAI21X1 _14807_ (
    .A(_4896__bF$buf4),
    .B(_4899__bF$buf8),
    .C(\datapath.registers.838[19] [18]),
    .Y(_4919_)
);

OAI21X1 _14808_ (
    .A(_4835__bF$buf2),
    .B(_4900__bF$buf1),
    .C(_4919_),
    .Y(_4091_)
);

OAI21X1 _14809_ (
    .A(_4896__bF$buf3),
    .B(_4899__bF$buf7),
    .C(\datapath.registers.838[19] [19]),
    .Y(_4920_)
);

OAI21X1 _14810_ (
    .A(_4837__bF$buf2),
    .B(_4900__bF$buf0),
    .C(_4920_),
    .Y(_4092_)
);

OAI21X1 _14811_ (
    .A(_4896__bF$buf2),
    .B(_4899__bF$buf6),
    .C(\datapath.registers.838[19] [20]),
    .Y(_4921_)
);

OAI21X1 _14812_ (
    .A(_4839__bF$buf2),
    .B(_4900__bF$buf4),
    .C(_4921_),
    .Y(_4094_)
);

OAI21X1 _14813_ (
    .A(_4896__bF$buf1),
    .B(_4899__bF$buf5),
    .C(\datapath.registers.838[19] [21]),
    .Y(_4922_)
);

OAI21X1 _14814_ (
    .A(_4841__bF$buf2),
    .B(_4900__bF$buf3),
    .C(_4922_),
    .Y(_4095_)
);

OAI21X1 _14815_ (
    .A(_4896__bF$buf0),
    .B(_4899__bF$buf4),
    .C(\datapath.registers.838[19] [22]),
    .Y(_4923_)
);

OAI21X1 _14816_ (
    .A(_4843__bF$buf2),
    .B(_4900__bF$buf2),
    .C(_4923_),
    .Y(_4096_)
);

OAI21X1 _14817_ (
    .A(_4896__bF$buf5),
    .B(_4899__bF$buf3),
    .C(\datapath.registers.838[19] [23]),
    .Y(_4924_)
);

OAI21X1 _14818_ (
    .A(_4845__bF$buf2),
    .B(_4900__bF$buf1),
    .C(_4924_),
    .Y(_4097_)
);

OAI21X1 _14819_ (
    .A(_4896__bF$buf4),
    .B(_4899__bF$buf2),
    .C(\datapath.registers.838[19] [24]),
    .Y(_4925_)
);

OAI21X1 _14820_ (
    .A(_4847__bF$buf2),
    .B(_4900__bF$buf0),
    .C(_4925_),
    .Y(_4098_)
);

OAI21X1 _14821_ (
    .A(_4896__bF$buf3),
    .B(_4899__bF$buf1),
    .C(\datapath.registers.838[19] [25]),
    .Y(_4926_)
);

OAI21X1 _14822_ (
    .A(_4849__bF$buf2),
    .B(_4900__bF$buf4),
    .C(_4926_),
    .Y(_4099_)
);

OAI21X1 _14823_ (
    .A(_4896__bF$buf2),
    .B(_4899__bF$buf0),
    .C(\datapath.registers.838[19] [26]),
    .Y(_4927_)
);

OAI21X1 _14824_ (
    .A(_4851__bF$buf2),
    .B(_4900__bF$buf3),
    .C(_4927_),
    .Y(_4100_)
);

OAI21X1 _14825_ (
    .A(_4896__bF$buf1),
    .B(_4899__bF$buf13),
    .C(\datapath.registers.838[19] [27]),
    .Y(_4928_)
);

OAI21X1 _14826_ (
    .A(_4853__bF$buf2),
    .B(_4900__bF$buf2),
    .C(_4928_),
    .Y(_4101_)
);

OAI21X1 _14827_ (
    .A(_4896__bF$buf0),
    .B(_4899__bF$buf12),
    .C(\datapath.registers.838[19] [28]),
    .Y(_4929_)
);

OAI21X1 _14828_ (
    .A(_4855__bF$buf2),
    .B(_4900__bF$buf1),
    .C(_4929_),
    .Y(_4102_)
);

OAI21X1 _14829_ (
    .A(_4896__bF$buf5),
    .B(_4899__bF$buf11),
    .C(\datapath.registers.838[19] [29]),
    .Y(_4930_)
);

OAI21X1 _14830_ (
    .A(_4857__bF$buf2),
    .B(_4900__bF$buf0),
    .C(_4930_),
    .Y(_4103_)
);

OAI21X1 _14831_ (
    .A(_4896__bF$buf4),
    .B(_4899__bF$buf10),
    .C(\datapath.registers.838[19] [30]),
    .Y(_4931_)
);

OAI21X1 _14832_ (
    .A(_4859__bF$buf2),
    .B(_4900__bF$buf4),
    .C(_4931_),
    .Y(_4105_)
);

OAI21X1 _14833_ (
    .A(_4896__bF$buf3),
    .B(_4899__bF$buf9),
    .C(\datapath.registers.838[19] [31]),
    .Y(_4932_)
);

OAI21X1 _14834_ (
    .A(_4861__bF$buf2),
    .B(_4900__bF$buf3),
    .C(_4932_),
    .Y(_4106_)
);

NOR2X1 _14835_ (
    .A(\datapath.wbinstr [7]),
    .B(_4897_),
    .Y(_4933_)
);

NAND2X1 _14836_ (
    .A(\controlunit.regfile_wen ),
    .B(_4933_),
    .Y(_4934_)
);

NOR2X1 _14837_ (
    .A(_4896__bF$buf2),
    .B(_4934__bF$buf9),
    .Y(_4935_)
);

NOR2X1 _14838_ (
    .A(\datapath.registers.838[18] [0]),
    .B(_4935__bF$buf7),
    .Y(_4936_)
);

AOI21X1 _14839_ (
    .A(_4786__bF$buf1),
    .B(_4935__bF$buf6),
    .C(_4936_),
    .Y(_4050_)
);

NOR2X1 _14840_ (
    .A(\datapath.registers.838[18] [1]),
    .B(_4935__bF$buf5),
    .Y(_4937_)
);

AOI21X1 _14841_ (
    .A(_4801__bF$buf1),
    .B(_4935__bF$buf4),
    .C(_4937_),
    .Y(_4061_)
);

NOR2X1 _14842_ (
    .A(\datapath.registers.838[18] [2]),
    .B(_4935__bF$buf3),
    .Y(_4938_)
);

AOI21X1 _14843_ (
    .A(_4803__bF$buf1),
    .B(_4935__bF$buf2),
    .C(_4938_),
    .Y(_4072_)
);

NOR2X1 _14844_ (
    .A(\datapath.registers.838[18] [3]),
    .B(_4935__bF$buf1),
    .Y(_4939_)
);

AOI21X1 _14845_ (
    .A(_4805__bF$buf1),
    .B(_4935__bF$buf0),
    .C(_4939_),
    .Y(_4075_)
);

NOR2X1 _14846_ (
    .A(\datapath.registers.838[18] [4]),
    .B(_4935__bF$buf7),
    .Y(_4940_)
);

AOI21X1 _14847_ (
    .A(_4807__bF$buf1),
    .B(_4935__bF$buf6),
    .C(_4940_),
    .Y(_4076_)
);

NOR2X1 _14848_ (
    .A(\datapath.registers.838[18] [5]),
    .B(_4935__bF$buf5),
    .Y(_4941_)
);

AOI21X1 _14849_ (
    .A(_4809__bF$buf1),
    .B(_4935__bF$buf4),
    .C(_4941_),
    .Y(_4077_)
);

NOR2X1 _14850_ (
    .A(\datapath.registers.838[18] [6]),
    .B(_4935__bF$buf3),
    .Y(_4942_)
);

AOI21X1 _14851_ (
    .A(_4811__bF$buf1),
    .B(_4935__bF$buf2),
    .C(_4942_),
    .Y(_4078_)
);

NOR2X1 _14852_ (
    .A(\datapath.registers.838[18] [7]),
    .B(_4935__bF$buf1),
    .Y(_4943_)
);

AOI21X1 _14853_ (
    .A(_4813__bF$buf1),
    .B(_4935__bF$buf0),
    .C(_4943_),
    .Y(_4079_)
);

NOR2X1 _14854_ (
    .A(\datapath.registers.838[18] [8]),
    .B(_4935__bF$buf7),
    .Y(_4944_)
);

AOI21X1 _14855_ (
    .A(_4815__bF$buf1),
    .B(_4935__bF$buf6),
    .C(_4944_),
    .Y(_4080_)
);

NOR2X1 _14856_ (
    .A(\datapath.registers.838[18] [9]),
    .B(_4935__bF$buf5),
    .Y(_4945_)
);

AOI21X1 _14857_ (
    .A(_4817__bF$buf1),
    .B(_4935__bF$buf4),
    .C(_4945_),
    .Y(_4081_)
);

NOR2X1 _14858_ (
    .A(\datapath.registers.838[18] [10]),
    .B(_4935__bF$buf3),
    .Y(_4946_)
);

AOI21X1 _14859_ (
    .A(_4819__bF$buf1),
    .B(_4935__bF$buf2),
    .C(_4946_),
    .Y(_4051_)
);

NOR2X1 _14860_ (
    .A(\datapath.registers.838[18] [11]),
    .B(_4935__bF$buf1),
    .Y(_4947_)
);

AOI21X1 _14861_ (
    .A(_4821__bF$buf1),
    .B(_4935__bF$buf0),
    .C(_4947_),
    .Y(_4052_)
);

NOR2X1 _14862_ (
    .A(\datapath.registers.838[18] [12]),
    .B(_4935__bF$buf7),
    .Y(_4948_)
);

AOI21X1 _14863_ (
    .A(_4823__bF$buf1),
    .B(_4935__bF$buf6),
    .C(_4948_),
    .Y(_4053_)
);

NOR2X1 _14864_ (
    .A(\datapath.registers.838[18] [13]),
    .B(_4935__bF$buf5),
    .Y(_4949_)
);

AOI21X1 _14865_ (
    .A(_4825__bF$buf1),
    .B(_4935__bF$buf4),
    .C(_4949_),
    .Y(_4054_)
);

NOR2X1 _14866_ (
    .A(\datapath.registers.838[18] [14]),
    .B(_4935__bF$buf3),
    .Y(_4950_)
);

AOI21X1 _14867_ (
    .A(_4827__bF$buf1),
    .B(_4935__bF$buf2),
    .C(_4950_),
    .Y(_4055_)
);

NOR2X1 _14868_ (
    .A(\datapath.registers.838[18] [15]),
    .B(_4935__bF$buf1),
    .Y(_4951_)
);

AOI21X1 _14869_ (
    .A(_4829__bF$buf1),
    .B(_4935__bF$buf0),
    .C(_4951_),
    .Y(_4056_)
);

NOR2X1 _14870_ (
    .A(\datapath.registers.838[18] [16]),
    .B(_4935__bF$buf7),
    .Y(_4952_)
);

AOI21X1 _14871_ (
    .A(_4831__bF$buf1),
    .B(_4935__bF$buf6),
    .C(_4952_),
    .Y(_4057_)
);

NOR2X1 _14872_ (
    .A(\datapath.registers.838[18] [17]),
    .B(_4935__bF$buf5),
    .Y(_4953_)
);

AOI21X1 _14873_ (
    .A(_4833__bF$buf1),
    .B(_4935__bF$buf4),
    .C(_4953_),
    .Y(_4058_)
);

NOR2X1 _14874_ (
    .A(\datapath.registers.838[18] [18]),
    .B(_4935__bF$buf3),
    .Y(_4954_)
);

AOI21X1 _14875_ (
    .A(_4835__bF$buf1),
    .B(_4935__bF$buf2),
    .C(_4954_),
    .Y(_4059_)
);

NOR2X1 _14876_ (
    .A(\datapath.registers.838[18] [19]),
    .B(_4935__bF$buf1),
    .Y(_4955_)
);

AOI21X1 _14877_ (
    .A(_4837__bF$buf1),
    .B(_4935__bF$buf0),
    .C(_4955_),
    .Y(_4060_)
);

NOR2X1 _14878_ (
    .A(\datapath.registers.838[18] [20]),
    .B(_4935__bF$buf7),
    .Y(_4956_)
);

AOI21X1 _14879_ (
    .A(_4839__bF$buf1),
    .B(_4935__bF$buf6),
    .C(_4956_),
    .Y(_4062_)
);

NOR2X1 _14880_ (
    .A(\datapath.registers.838[18] [21]),
    .B(_4935__bF$buf5),
    .Y(_4957_)
);

AOI21X1 _14881_ (
    .A(_4841__bF$buf1),
    .B(_4935__bF$buf4),
    .C(_4957_),
    .Y(_4063_)
);

NOR2X1 _14882_ (
    .A(\datapath.registers.838[18] [22]),
    .B(_4935__bF$buf3),
    .Y(_4958_)
);

AOI21X1 _14883_ (
    .A(_4843__bF$buf1),
    .B(_4935__bF$buf2),
    .C(_4958_),
    .Y(_4064_)
);

NOR2X1 _14884_ (
    .A(\datapath.registers.838[18] [23]),
    .B(_4935__bF$buf1),
    .Y(_4959_)
);

AOI21X1 _14885_ (
    .A(_4845__bF$buf1),
    .B(_4935__bF$buf0),
    .C(_4959_),
    .Y(_4065_)
);

NOR2X1 _14886_ (
    .A(\datapath.registers.838[18] [24]),
    .B(_4935__bF$buf7),
    .Y(_4960_)
);

AOI21X1 _14887_ (
    .A(_4847__bF$buf1),
    .B(_4935__bF$buf6),
    .C(_4960_),
    .Y(_4066_)
);

NOR2X1 _14888_ (
    .A(\datapath.registers.838[18] [25]),
    .B(_4935__bF$buf5),
    .Y(_4961_)
);

AOI21X1 _14889_ (
    .A(_4849__bF$buf1),
    .B(_4935__bF$buf4),
    .C(_4961_),
    .Y(_4067_)
);

NOR2X1 _14890_ (
    .A(\datapath.registers.838[18] [26]),
    .B(_4935__bF$buf3),
    .Y(_4962_)
);

AOI21X1 _14891_ (
    .A(_4851__bF$buf1),
    .B(_4935__bF$buf2),
    .C(_4962_),
    .Y(_4068_)
);

NOR2X1 _14892_ (
    .A(\datapath.registers.838[18] [27]),
    .B(_4935__bF$buf1),
    .Y(_4963_)
);

AOI21X1 _14893_ (
    .A(_4853__bF$buf1),
    .B(_4935__bF$buf0),
    .C(_4963_),
    .Y(_4069_)
);

NOR2X1 _14894_ (
    .A(\datapath.registers.838[18] [28]),
    .B(_4935__bF$buf7),
    .Y(_4964_)
);

AOI21X1 _14895_ (
    .A(_4855__bF$buf1),
    .B(_4935__bF$buf6),
    .C(_4964_),
    .Y(_4070_)
);

NOR2X1 _14896_ (
    .A(\datapath.registers.838[18] [29]),
    .B(_4935__bF$buf5),
    .Y(_4965_)
);

AOI21X1 _14897_ (
    .A(_4857__bF$buf1),
    .B(_4935__bF$buf4),
    .C(_4965_),
    .Y(_4071_)
);

NOR2X1 _14898_ (
    .A(\datapath.registers.838[18] [30]),
    .B(_4935__bF$buf3),
    .Y(_4966_)
);

AOI21X1 _14899_ (
    .A(_4859__bF$buf1),
    .B(_4935__bF$buf2),
    .C(_4966_),
    .Y(_4073_)
);

NOR2X1 _14900_ (
    .A(\datapath.registers.838[18] [31]),
    .B(_4935__bF$buf1),
    .Y(_4967_)
);

AOI21X1 _14901_ (
    .A(_4861__bF$buf1),
    .B(_4935__bF$buf0),
    .C(_4967_),
    .Y(_4074_)
);

NAND2X1 _14902_ (
    .A(\controlunit.regfile_wen ),
    .B(_4788_),
    .Y(_4968_)
);

NOR2X1 _14903_ (
    .A(_4896__bF$buf1),
    .B(_4968__bF$buf9),
    .Y(_4969_)
);

NOR2X1 _14904_ (
    .A(\datapath.registers.838[17] [0]),
    .B(_4969__bF$buf7),
    .Y(_4970_)
);

AOI21X1 _14905_ (
    .A(_4786__bF$buf0),
    .B(_4969__bF$buf6),
    .C(_4970_),
    .Y(_4018_)
);

NOR2X1 _14906_ (
    .A(\datapath.registers.838[17] [1]),
    .B(_4969__bF$buf5),
    .Y(_4971_)
);

AOI21X1 _14907_ (
    .A(_4801__bF$buf0),
    .B(_4969__bF$buf4),
    .C(_4971_),
    .Y(_4029_)
);

NOR2X1 _14908_ (
    .A(\datapath.registers.838[17] [2]),
    .B(_4969__bF$buf3),
    .Y(_4972_)
);

AOI21X1 _14909_ (
    .A(_4803__bF$buf0),
    .B(_4969__bF$buf2),
    .C(_4972_),
    .Y(_4040_)
);

INVX1 _14910_ (
    .A(\datapath.registers.838[17] [3]),
    .Y(_4973_)
);

NAND2X1 _14911_ (
    .A(\datapath.rd [3]),
    .B(_4969__bF$buf1),
    .Y(_4974_)
);

OAI21X1 _14912_ (
    .A(_4973_),
    .B(_4969__bF$buf0),
    .C(_4974_),
    .Y(_4043_)
);

INVX1 _14913_ (
    .A(\datapath.registers.838[17] [4]),
    .Y(_4975_)
);

NAND2X1 _14914_ (
    .A(\datapath.rd [4]),
    .B(_4969__bF$buf7),
    .Y(_4976_)
);

OAI21X1 _14915_ (
    .A(_4975_),
    .B(_4969__bF$buf6),
    .C(_4976_),
    .Y(_4044_)
);

INVX1 _14916_ (
    .A(\datapath.registers.838[17] [5]),
    .Y(_4977_)
);

NAND2X1 _14917_ (
    .A(\datapath.rd [5]),
    .B(_4969__bF$buf5),
    .Y(_4978_)
);

OAI21X1 _14918_ (
    .A(_4977_),
    .B(_4969__bF$buf4),
    .C(_4978_),
    .Y(_4045_)
);

INVX1 _14919_ (
    .A(\datapath.registers.838[17] [6]),
    .Y(_4979_)
);

NAND2X1 _14920_ (
    .A(\datapath.rd [6]),
    .B(_4969__bF$buf3),
    .Y(_4980_)
);

OAI21X1 _14921_ (
    .A(_4979_),
    .B(_4969__bF$buf2),
    .C(_4980_),
    .Y(_4046_)
);

NOR2X1 _14922_ (
    .A(\datapath.registers.838[17] [7]),
    .B(_4969__bF$buf1),
    .Y(_4981_)
);

AOI21X1 _14923_ (
    .A(_4813__bF$buf0),
    .B(_4969__bF$buf0),
    .C(_4981_),
    .Y(_4047_)
);

NOR2X1 _14924_ (
    .A(\datapath.registers.838[17] [8]),
    .B(_4969__bF$buf7),
    .Y(_4982_)
);

AOI21X1 _14925_ (
    .A(_4815__bF$buf0),
    .B(_4969__bF$buf6),
    .C(_4982_),
    .Y(_4048_)
);

INVX1 _14926_ (
    .A(\datapath.registers.838[17] [9]),
    .Y(_4983_)
);

NAND2X1 _14927_ (
    .A(\datapath.rd [9]),
    .B(_4969__bF$buf5),
    .Y(_4984_)
);

OAI21X1 _14928_ (
    .A(_4983_),
    .B(_4969__bF$buf4),
    .C(_4984_),
    .Y(_4049_)
);

INVX1 _14929_ (
    .A(\datapath.registers.838[17] [10]),
    .Y(_4985_)
);

NAND2X1 _14930_ (
    .A(\datapath.rd [10]),
    .B(_4969__bF$buf3),
    .Y(_4986_)
);

OAI21X1 _14931_ (
    .A(_4985_),
    .B(_4969__bF$buf2),
    .C(_4986_),
    .Y(_4019_)
);

NOR2X1 _14932_ (
    .A(\datapath.registers.838[17] [11]),
    .B(_4969__bF$buf1),
    .Y(_4987_)
);

AOI21X1 _14933_ (
    .A(_4821__bF$buf0),
    .B(_4969__bF$buf0),
    .C(_4987_),
    .Y(_4020_)
);

NOR2X1 _14934_ (
    .A(\datapath.registers.838[17] [12]),
    .B(_4969__bF$buf7),
    .Y(_4988_)
);

AOI21X1 _14935_ (
    .A(_4823__bF$buf0),
    .B(_4969__bF$buf6),
    .C(_4988_),
    .Y(_4021_)
);

NOR2X1 _14936_ (
    .A(\datapath.registers.838[17] [13]),
    .B(_4969__bF$buf5),
    .Y(_4989_)
);

AOI21X1 _14937_ (
    .A(_4825__bF$buf0),
    .B(_4969__bF$buf4),
    .C(_4989_),
    .Y(_4022_)
);

NOR2X1 _14938_ (
    .A(\datapath.registers.838[17] [14]),
    .B(_4969__bF$buf3),
    .Y(_4990_)
);

AOI21X1 _14939_ (
    .A(_4827__bF$buf0),
    .B(_4969__bF$buf2),
    .C(_4990_),
    .Y(_4023_)
);

NOR2X1 _14940_ (
    .A(\datapath.registers.838[17] [15]),
    .B(_4969__bF$buf1),
    .Y(_4991_)
);

AOI21X1 _14941_ (
    .A(_4829__bF$buf0),
    .B(_4969__bF$buf0),
    .C(_4991_),
    .Y(_4024_)
);

NOR2X1 _14942_ (
    .A(\datapath.registers.838[17] [16]),
    .B(_4969__bF$buf7),
    .Y(_4992_)
);

AOI21X1 _14943_ (
    .A(_4831__bF$buf0),
    .B(_4969__bF$buf6),
    .C(_4992_),
    .Y(_4025_)
);

NOR2X1 _14944_ (
    .A(\datapath.registers.838[17] [17]),
    .B(_4969__bF$buf5),
    .Y(_4993_)
);

AOI21X1 _14945_ (
    .A(_4833__bF$buf0),
    .B(_4969__bF$buf4),
    .C(_4993_),
    .Y(_4026_)
);

NOR2X1 _14946_ (
    .A(\datapath.registers.838[17] [18]),
    .B(_4969__bF$buf3),
    .Y(_4994_)
);

AOI21X1 _14947_ (
    .A(_4835__bF$buf0),
    .B(_4969__bF$buf2),
    .C(_4994_),
    .Y(_4027_)
);

INVX1 _14948_ (
    .A(\datapath.registers.838[17] [19]),
    .Y(_4995_)
);

NAND2X1 _14949_ (
    .A(\datapath.rd [19]),
    .B(_4969__bF$buf1),
    .Y(_4996_)
);

OAI21X1 _14950_ (
    .A(_4995_),
    .B(_4969__bF$buf0),
    .C(_4996_),
    .Y(_4028_)
);

NOR2X1 _14951_ (
    .A(\datapath.registers.838[17] [20]),
    .B(_4969__bF$buf7),
    .Y(_4997_)
);

AOI21X1 _14952_ (
    .A(_4839__bF$buf0),
    .B(_4969__bF$buf6),
    .C(_4997_),
    .Y(_4030_)
);

INVX1 _14953_ (
    .A(\datapath.registers.838[17] [21]),
    .Y(_4998_)
);

NAND2X1 _14954_ (
    .A(\datapath.rd [21]),
    .B(_4969__bF$buf5),
    .Y(_4999_)
);

OAI21X1 _14955_ (
    .A(_4998_),
    .B(_4969__bF$buf4),
    .C(_4999_),
    .Y(_4031_)
);

INVX1 _14956_ (
    .A(\datapath.registers.838[17] [22]),
    .Y(_5000_)
);

NAND2X1 _14957_ (
    .A(\datapath.rd [22]),
    .B(_4969__bF$buf3),
    .Y(_5001_)
);

OAI21X1 _14958_ (
    .A(_5000_),
    .B(_4969__bF$buf2),
    .C(_5001_),
    .Y(_4032_)
);

INVX1 _14959_ (
    .A(\datapath.registers.838[17] [23]),
    .Y(_5002_)
);

NAND2X1 _14960_ (
    .A(\datapath.rd [23]),
    .B(_4969__bF$buf1),
    .Y(_5003_)
);

OAI21X1 _14961_ (
    .A(_5002_),
    .B(_4969__bF$buf0),
    .C(_5003_),
    .Y(_4033_)
);

INVX1 _14962_ (
    .A(\datapath.registers.838[17] [24]),
    .Y(_5004_)
);

NAND2X1 _14963_ (
    .A(\datapath.rd [24]),
    .B(_4969__bF$buf7),
    .Y(_5005_)
);

OAI21X1 _14964_ (
    .A(_5004_),
    .B(_4969__bF$buf6),
    .C(_5005_),
    .Y(_4034_)
);

INVX1 _14965_ (
    .A(\datapath.registers.838[17] [25]),
    .Y(_5006_)
);

NAND2X1 _14966_ (
    .A(\datapath.rd [25]),
    .B(_4969__bF$buf5),
    .Y(_5007_)
);

OAI21X1 _14967_ (
    .A(_5006_),
    .B(_4969__bF$buf4),
    .C(_5007_),
    .Y(_4035_)
);

NOR2X1 _14968_ (
    .A(\datapath.registers.838[17] [26]),
    .B(_4969__bF$buf3),
    .Y(_5008_)
);

AOI21X1 _14969_ (
    .A(_4851__bF$buf0),
    .B(_4969__bF$buf2),
    .C(_5008_),
    .Y(_4036_)
);

INVX1 _14970_ (
    .A(\datapath.registers.838[17] [27]),
    .Y(_5009_)
);

NAND2X1 _14971_ (
    .A(\datapath.rd [27]),
    .B(_4969__bF$buf1),
    .Y(_5010_)
);

OAI21X1 _14972_ (
    .A(_5009_),
    .B(_4969__bF$buf0),
    .C(_5010_),
    .Y(_4037_)
);

NOR2X1 _14973_ (
    .A(\datapath.registers.838[17] [28]),
    .B(_4969__bF$buf7),
    .Y(_5011_)
);

AOI21X1 _14974_ (
    .A(_4855__bF$buf0),
    .B(_4969__bF$buf6),
    .C(_5011_),
    .Y(_4038_)
);

NOR2X1 _14975_ (
    .A(\datapath.registers.838[17] [29]),
    .B(_4969__bF$buf5),
    .Y(_5012_)
);

AOI21X1 _14976_ (
    .A(_4857__bF$buf0),
    .B(_4969__bF$buf4),
    .C(_5012_),
    .Y(_4039_)
);

NOR2X1 _14977_ (
    .A(\datapath.registers.838[17] [30]),
    .B(_4969__bF$buf3),
    .Y(_5013_)
);

AOI21X1 _14978_ (
    .A(_4859__bF$buf0),
    .B(_4969__bF$buf2),
    .C(_5013_),
    .Y(_4041_)
);

NOR2X1 _14979_ (
    .A(\datapath.registers.838[17] [31]),
    .B(_4969__bF$buf1),
    .Y(_5014_)
);

AOI21X1 _14980_ (
    .A(_4861__bF$buf0),
    .B(_4969__bF$buf0),
    .C(_5014_),
    .Y(_4042_)
);

INVX2 _14981_ (
    .A(_4795_),
    .Y(_5015_)
);

NOR2X1 _14982_ (
    .A(_4790_),
    .B(_4896__bF$buf0),
    .Y(_5016_)
);

NAND2X1 _14983_ (
    .A(_5016_),
    .B(_5015_),
    .Y(_5017_)
);

NAND2X1 _14984_ (
    .A(\datapath.registers.838[16] [0]),
    .B(_5017__bF$buf7),
    .Y(_5018_)
);

OAI21X1 _14985_ (
    .A(_4786__bF$buf4),
    .B(_5017__bF$buf6),
    .C(_5018_),
    .Y(_3986_)
);

NAND2X1 _14986_ (
    .A(\datapath.registers.838[16] [1]),
    .B(_5017__bF$buf5),
    .Y(_5019_)
);

OAI21X1 _14987_ (
    .A(_4801__bF$buf4),
    .B(_5017__bF$buf4),
    .C(_5019_),
    .Y(_3997_)
);

NAND2X1 _14988_ (
    .A(\datapath.registers.838[16] [2]),
    .B(_5017__bF$buf3),
    .Y(_5020_)
);

OAI21X1 _14989_ (
    .A(_4803__bF$buf4),
    .B(_5017__bF$buf2),
    .C(_5020_),
    .Y(_4008_)
);

NAND2X1 _14990_ (
    .A(\datapath.registers.838[16] [3]),
    .B(_5017__bF$buf1),
    .Y(_5021_)
);

OAI21X1 _14991_ (
    .A(_4805__bF$buf0),
    .B(_5017__bF$buf0),
    .C(_5021_),
    .Y(_4011_)
);

NAND2X1 _14992_ (
    .A(\datapath.registers.838[16] [4]),
    .B(_5017__bF$buf7),
    .Y(_5022_)
);

OAI21X1 _14993_ (
    .A(_4807__bF$buf0),
    .B(_5017__bF$buf6),
    .C(_5022_),
    .Y(_4012_)
);

NAND2X1 _14994_ (
    .A(\datapath.registers.838[16] [5]),
    .B(_5017__bF$buf5),
    .Y(_5023_)
);

OAI21X1 _14995_ (
    .A(_4809__bF$buf0),
    .B(_5017__bF$buf4),
    .C(_5023_),
    .Y(_4013_)
);

NAND2X1 _14996_ (
    .A(\datapath.registers.838[16] [6]),
    .B(_5017__bF$buf3),
    .Y(_5024_)
);

OAI21X1 _14997_ (
    .A(_4811__bF$buf0),
    .B(_5017__bF$buf2),
    .C(_5024_),
    .Y(_4014_)
);

NAND2X1 _14998_ (
    .A(\datapath.registers.838[16] [7]),
    .B(_5017__bF$buf1),
    .Y(_5025_)
);

OAI21X1 _14999_ (
    .A(_4813__bF$buf4),
    .B(_5017__bF$buf0),
    .C(_5025_),
    .Y(_4015_)
);

NAND2X1 _15000_ (
    .A(\datapath.registers.838[16] [8]),
    .B(_5017__bF$buf7),
    .Y(_5026_)
);

OAI21X1 _15001_ (
    .A(_4815__bF$buf4),
    .B(_5017__bF$buf6),
    .C(_5026_),
    .Y(_4016_)
);

NAND2X1 _15002_ (
    .A(\datapath.registers.838[16] [9]),
    .B(_5017__bF$buf5),
    .Y(_5027_)
);

OAI21X1 _15003_ (
    .A(_4817__bF$buf0),
    .B(_5017__bF$buf4),
    .C(_5027_),
    .Y(_4017_)
);

NAND2X1 _15004_ (
    .A(\datapath.registers.838[16] [10]),
    .B(_5017__bF$buf3),
    .Y(_5028_)
);

OAI21X1 _15005_ (
    .A(_4819__bF$buf0),
    .B(_5017__bF$buf2),
    .C(_5028_),
    .Y(_3987_)
);

NAND2X1 _15006_ (
    .A(\datapath.registers.838[16] [11]),
    .B(_5017__bF$buf1),
    .Y(_5029_)
);

OAI21X1 _15007_ (
    .A(_4821__bF$buf4),
    .B(_5017__bF$buf0),
    .C(_5029_),
    .Y(_3988_)
);

NAND2X1 _15008_ (
    .A(\datapath.registers.838[16] [12]),
    .B(_5017__bF$buf7),
    .Y(_5030_)
);

OAI21X1 _15009_ (
    .A(_4823__bF$buf4),
    .B(_5017__bF$buf6),
    .C(_5030_),
    .Y(_3989_)
);

NAND2X1 _15010_ (
    .A(\datapath.registers.838[16] [13]),
    .B(_5017__bF$buf5),
    .Y(_5031_)
);

OAI21X1 _15011_ (
    .A(_4825__bF$buf4),
    .B(_5017__bF$buf4),
    .C(_5031_),
    .Y(_3990_)
);

NAND2X1 _15012_ (
    .A(\datapath.registers.838[16] [14]),
    .B(_5017__bF$buf3),
    .Y(_5032_)
);

OAI21X1 _15013_ (
    .A(_4827__bF$buf4),
    .B(_5017__bF$buf2),
    .C(_5032_),
    .Y(_3991_)
);

NAND2X1 _15014_ (
    .A(\datapath.registers.838[16] [15]),
    .B(_5017__bF$buf1),
    .Y(_5033_)
);

OAI21X1 _15015_ (
    .A(_4829__bF$buf4),
    .B(_5017__bF$buf0),
    .C(_5033_),
    .Y(_3992_)
);

NAND2X1 _15016_ (
    .A(\datapath.registers.838[16] [16]),
    .B(_5017__bF$buf7),
    .Y(_5034_)
);

OAI21X1 _15017_ (
    .A(_4831__bF$buf4),
    .B(_5017__bF$buf6),
    .C(_5034_),
    .Y(_3993_)
);

NAND2X1 _15018_ (
    .A(\datapath.registers.838[16] [17]),
    .B(_5017__bF$buf5),
    .Y(_5035_)
);

OAI21X1 _15019_ (
    .A(_4833__bF$buf4),
    .B(_5017__bF$buf4),
    .C(_5035_),
    .Y(_3994_)
);

NAND2X1 _15020_ (
    .A(\datapath.registers.838[16] [18]),
    .B(_5017__bF$buf3),
    .Y(_5036_)
);

OAI21X1 _15021_ (
    .A(_4835__bF$buf4),
    .B(_5017__bF$buf2),
    .C(_5036_),
    .Y(_3995_)
);

NAND2X1 _15022_ (
    .A(\datapath.registers.838[16] [19]),
    .B(_5017__bF$buf1),
    .Y(_5037_)
);

OAI21X1 _15023_ (
    .A(_4837__bF$buf0),
    .B(_5017__bF$buf0),
    .C(_5037_),
    .Y(_3996_)
);

NAND2X1 _15024_ (
    .A(\datapath.registers.838[16] [20]),
    .B(_5017__bF$buf7),
    .Y(_5038_)
);

OAI21X1 _15025_ (
    .A(_4839__bF$buf4),
    .B(_5017__bF$buf6),
    .C(_5038_),
    .Y(_3998_)
);

NAND2X1 _15026_ (
    .A(\datapath.registers.838[16] [21]),
    .B(_5017__bF$buf5),
    .Y(_5039_)
);

OAI21X1 _15027_ (
    .A(_4841__bF$buf0),
    .B(_5017__bF$buf4),
    .C(_5039_),
    .Y(_3999_)
);

NAND2X1 _15028_ (
    .A(\datapath.registers.838[16] [22]),
    .B(_5017__bF$buf3),
    .Y(_5040_)
);

OAI21X1 _15029_ (
    .A(_4843__bF$buf0),
    .B(_5017__bF$buf2),
    .C(_5040_),
    .Y(_4000_)
);

NAND2X1 _15030_ (
    .A(\datapath.registers.838[16] [23]),
    .B(_5017__bF$buf1),
    .Y(_5041_)
);

OAI21X1 _15031_ (
    .A(_4845__bF$buf0),
    .B(_5017__bF$buf0),
    .C(_5041_),
    .Y(_4001_)
);

NAND2X1 _15032_ (
    .A(\datapath.registers.838[16] [24]),
    .B(_5017__bF$buf7),
    .Y(_5042_)
);

OAI21X1 _15033_ (
    .A(_4847__bF$buf0),
    .B(_5017__bF$buf6),
    .C(_5042_),
    .Y(_4002_)
);

NAND2X1 _15034_ (
    .A(\datapath.registers.838[16] [25]),
    .B(_5017__bF$buf5),
    .Y(_5043_)
);

OAI21X1 _15035_ (
    .A(_4849__bF$buf0),
    .B(_5017__bF$buf4),
    .C(_5043_),
    .Y(_4003_)
);

NAND2X1 _15036_ (
    .A(\datapath.registers.838[16] [26]),
    .B(_5017__bF$buf3),
    .Y(_5044_)
);

OAI21X1 _15037_ (
    .A(_4851__bF$buf4),
    .B(_5017__bF$buf2),
    .C(_5044_),
    .Y(_4004_)
);

NAND2X1 _15038_ (
    .A(\datapath.registers.838[16] [27]),
    .B(_5017__bF$buf1),
    .Y(_5045_)
);

OAI21X1 _15039_ (
    .A(_4853__bF$buf0),
    .B(_5017__bF$buf0),
    .C(_5045_),
    .Y(_4005_)
);

NAND2X1 _15040_ (
    .A(\datapath.registers.838[16] [28]),
    .B(_5017__bF$buf7),
    .Y(_5046_)
);

OAI21X1 _15041_ (
    .A(_4855__bF$buf4),
    .B(_5017__bF$buf6),
    .C(_5046_),
    .Y(_4006_)
);

NAND2X1 _15042_ (
    .A(\datapath.registers.838[16] [29]),
    .B(_5017__bF$buf5),
    .Y(_5047_)
);

OAI21X1 _15043_ (
    .A(_4857__bF$buf4),
    .B(_5017__bF$buf4),
    .C(_5047_),
    .Y(_4007_)
);

NAND2X1 _15044_ (
    .A(\datapath.registers.838[16] [30]),
    .B(_5017__bF$buf3),
    .Y(_5048_)
);

OAI21X1 _15045_ (
    .A(_4859__bF$buf4),
    .B(_5017__bF$buf2),
    .C(_5048_),
    .Y(_4009_)
);

NAND2X1 _15046_ (
    .A(\datapath.registers.838[16] [31]),
    .B(_5017__bF$buf1),
    .Y(_5049_)
);

OAI21X1 _15047_ (
    .A(_4861__bF$buf4),
    .B(_5017__bF$buf0),
    .C(_5049_),
    .Y(_4010_)
);

NAND2X1 _15048_ (
    .A(\datapath.wbinstr [10]),
    .B(_4793_),
    .Y(_5050_)
);

OR2X2 _15049_ (
    .A(_5050_),
    .B(_4791_),
    .Y(_5051_)
);

OR2X2 _15050_ (
    .A(_5051__bF$buf5),
    .B(_4899__bF$buf8),
    .Y(_5052_)
);

OAI21X1 _15051_ (
    .A(_4899__bF$buf7),
    .B(_5051__bF$buf4),
    .C(\datapath.registers.838[15] [0]),
    .Y(_5053_)
);

OAI21X1 _15052_ (
    .A(_4786__bF$buf3),
    .B(_5052__bF$buf4),
    .C(_5053_),
    .Y(_3954_)
);

OAI21X1 _15053_ (
    .A(_4899__bF$buf6),
    .B(_5051__bF$buf3),
    .C(\datapath.registers.838[15] [1]),
    .Y(_5054_)
);

OAI21X1 _15054_ (
    .A(_4801__bF$buf3),
    .B(_5052__bF$buf3),
    .C(_5054_),
    .Y(_3965_)
);

OAI21X1 _15055_ (
    .A(_4899__bF$buf5),
    .B(_5051__bF$buf2),
    .C(\datapath.registers.838[15] [2]),
    .Y(_5055_)
);

OAI21X1 _15056_ (
    .A(_4803__bF$buf3),
    .B(_5052__bF$buf2),
    .C(_5055_),
    .Y(_3976_)
);

OAI21X1 _15057_ (
    .A(_4899__bF$buf4),
    .B(_5051__bF$buf1),
    .C(\datapath.registers.838[15] [3]),
    .Y(_5056_)
);

OAI21X1 _15058_ (
    .A(_4805__bF$buf4),
    .B(_5052__bF$buf1),
    .C(_5056_),
    .Y(_3979_)
);

OAI21X1 _15059_ (
    .A(_4899__bF$buf3),
    .B(_5051__bF$buf0),
    .C(\datapath.registers.838[15] [4]),
    .Y(_5057_)
);

OAI21X1 _15060_ (
    .A(_4807__bF$buf4),
    .B(_5052__bF$buf0),
    .C(_5057_),
    .Y(_3980_)
);

OAI21X1 _15061_ (
    .A(_4899__bF$buf2),
    .B(_5051__bF$buf5),
    .C(\datapath.registers.838[15] [5]),
    .Y(_5058_)
);

OAI21X1 _15062_ (
    .A(_4809__bF$buf4),
    .B(_5052__bF$buf4),
    .C(_5058_),
    .Y(_3981_)
);

OAI21X1 _15063_ (
    .A(_4899__bF$buf1),
    .B(_5051__bF$buf4),
    .C(\datapath.registers.838[15] [6]),
    .Y(_5059_)
);

OAI21X1 _15064_ (
    .A(_4811__bF$buf4),
    .B(_5052__bF$buf3),
    .C(_5059_),
    .Y(_3982_)
);

OAI21X1 _15065_ (
    .A(_4899__bF$buf0),
    .B(_5051__bF$buf3),
    .C(\datapath.registers.838[15] [7]),
    .Y(_5060_)
);

OAI21X1 _15066_ (
    .A(_4813__bF$buf3),
    .B(_5052__bF$buf2),
    .C(_5060_),
    .Y(_3983_)
);

OAI21X1 _15067_ (
    .A(_4899__bF$buf13),
    .B(_5051__bF$buf2),
    .C(\datapath.registers.838[15] [8]),
    .Y(_5061_)
);

OAI21X1 _15068_ (
    .A(_4815__bF$buf3),
    .B(_5052__bF$buf1),
    .C(_5061_),
    .Y(_3984_)
);

OAI21X1 _15069_ (
    .A(_4899__bF$buf12),
    .B(_5051__bF$buf1),
    .C(\datapath.registers.838[15] [9]),
    .Y(_5062_)
);

OAI21X1 _15070_ (
    .A(_4817__bF$buf4),
    .B(_5052__bF$buf0),
    .C(_5062_),
    .Y(_3985_)
);

OAI21X1 _15071_ (
    .A(_4899__bF$buf11),
    .B(_5051__bF$buf0),
    .C(\datapath.registers.838[15] [10]),
    .Y(_5063_)
);

OAI21X1 _15072_ (
    .A(_4819__bF$buf4),
    .B(_5052__bF$buf4),
    .C(_5063_),
    .Y(_3955_)
);

OAI21X1 _15073_ (
    .A(_4899__bF$buf10),
    .B(_5051__bF$buf5),
    .C(\datapath.registers.838[15] [11]),
    .Y(_5064_)
);

OAI21X1 _15074_ (
    .A(_4821__bF$buf3),
    .B(_5052__bF$buf3),
    .C(_5064_),
    .Y(_3956_)
);

OAI21X1 _15075_ (
    .A(_4899__bF$buf9),
    .B(_5051__bF$buf4),
    .C(\datapath.registers.838[15] [12]),
    .Y(_5065_)
);

OAI21X1 _15076_ (
    .A(_4823__bF$buf3),
    .B(_5052__bF$buf2),
    .C(_5065_),
    .Y(_3957_)
);

OAI21X1 _15077_ (
    .A(_4899__bF$buf8),
    .B(_5051__bF$buf3),
    .C(\datapath.registers.838[15] [13]),
    .Y(_5066_)
);

OAI21X1 _15078_ (
    .A(_4825__bF$buf3),
    .B(_5052__bF$buf1),
    .C(_5066_),
    .Y(_3958_)
);

OAI21X1 _15079_ (
    .A(_4899__bF$buf7),
    .B(_5051__bF$buf2),
    .C(\datapath.registers.838[15] [14]),
    .Y(_5067_)
);

OAI21X1 _15080_ (
    .A(_4827__bF$buf3),
    .B(_5052__bF$buf0),
    .C(_5067_),
    .Y(_3959_)
);

OAI21X1 _15081_ (
    .A(_4899__bF$buf6),
    .B(_5051__bF$buf1),
    .C(\datapath.registers.838[15] [15]),
    .Y(_5068_)
);

OAI21X1 _15082_ (
    .A(_4829__bF$buf3),
    .B(_5052__bF$buf4),
    .C(_5068_),
    .Y(_3960_)
);

OAI21X1 _15083_ (
    .A(_4899__bF$buf5),
    .B(_5051__bF$buf0),
    .C(\datapath.registers.838[15] [16]),
    .Y(_5069_)
);

OAI21X1 _15084_ (
    .A(_4831__bF$buf3),
    .B(_5052__bF$buf3),
    .C(_5069_),
    .Y(_3961_)
);

OAI21X1 _15085_ (
    .A(_4899__bF$buf4),
    .B(_5051__bF$buf5),
    .C(\datapath.registers.838[15] [17]),
    .Y(_5070_)
);

OAI21X1 _15086_ (
    .A(_4833__bF$buf3),
    .B(_5052__bF$buf2),
    .C(_5070_),
    .Y(_3962_)
);

OAI21X1 _15087_ (
    .A(_4899__bF$buf3),
    .B(_5051__bF$buf4),
    .C(\datapath.registers.838[15] [18]),
    .Y(_5071_)
);

OAI21X1 _15088_ (
    .A(_4835__bF$buf3),
    .B(_5052__bF$buf1),
    .C(_5071_),
    .Y(_3963_)
);

OAI21X1 _15089_ (
    .A(_4899__bF$buf2),
    .B(_5051__bF$buf3),
    .C(\datapath.registers.838[15] [19]),
    .Y(_5072_)
);

OAI21X1 _15090_ (
    .A(_4837__bF$buf4),
    .B(_5052__bF$buf0),
    .C(_5072_),
    .Y(_3964_)
);

OAI21X1 _15091_ (
    .A(_4899__bF$buf1),
    .B(_5051__bF$buf2),
    .C(\datapath.registers.838[15] [20]),
    .Y(_5073_)
);

OAI21X1 _15092_ (
    .A(_4839__bF$buf3),
    .B(_5052__bF$buf4),
    .C(_5073_),
    .Y(_3966_)
);

OAI21X1 _15093_ (
    .A(_4899__bF$buf0),
    .B(_5051__bF$buf1),
    .C(\datapath.registers.838[15] [21]),
    .Y(_5074_)
);

OAI21X1 _15094_ (
    .A(_4841__bF$buf4),
    .B(_5052__bF$buf3),
    .C(_5074_),
    .Y(_3967_)
);

OAI21X1 _15095_ (
    .A(_4899__bF$buf13),
    .B(_5051__bF$buf0),
    .C(\datapath.registers.838[15] [22]),
    .Y(_5075_)
);

OAI21X1 _15096_ (
    .A(_4843__bF$buf4),
    .B(_5052__bF$buf2),
    .C(_5075_),
    .Y(_3968_)
);

OAI21X1 _15097_ (
    .A(_4899__bF$buf12),
    .B(_5051__bF$buf5),
    .C(\datapath.registers.838[15] [23]),
    .Y(_5076_)
);

OAI21X1 _15098_ (
    .A(_4845__bF$buf4),
    .B(_5052__bF$buf1),
    .C(_5076_),
    .Y(_3969_)
);

OAI21X1 _15099_ (
    .A(_4899__bF$buf11),
    .B(_5051__bF$buf4),
    .C(\datapath.registers.838[15] [24]),
    .Y(_5077_)
);

OAI21X1 _15100_ (
    .A(_4847__bF$buf4),
    .B(_5052__bF$buf0),
    .C(_5077_),
    .Y(_3970_)
);

OAI21X1 _15101_ (
    .A(_4899__bF$buf10),
    .B(_5051__bF$buf3),
    .C(\datapath.registers.838[15] [25]),
    .Y(_5078_)
);

OAI21X1 _15102_ (
    .A(_4849__bF$buf4),
    .B(_5052__bF$buf4),
    .C(_5078_),
    .Y(_3971_)
);

OAI21X1 _15103_ (
    .A(_4899__bF$buf9),
    .B(_5051__bF$buf2),
    .C(\datapath.registers.838[15] [26]),
    .Y(_5079_)
);

OAI21X1 _15104_ (
    .A(_4851__bF$buf3),
    .B(_5052__bF$buf3),
    .C(_5079_),
    .Y(_3972_)
);

OAI21X1 _15105_ (
    .A(_4899__bF$buf8),
    .B(_5051__bF$buf1),
    .C(\datapath.registers.838[15] [27]),
    .Y(_5080_)
);

OAI21X1 _15106_ (
    .A(_4853__bF$buf4),
    .B(_5052__bF$buf2),
    .C(_5080_),
    .Y(_3973_)
);

OAI21X1 _15107_ (
    .A(_4899__bF$buf7),
    .B(_5051__bF$buf0),
    .C(\datapath.registers.838[15] [28]),
    .Y(_5081_)
);

OAI21X1 _15108_ (
    .A(_4855__bF$buf3),
    .B(_5052__bF$buf1),
    .C(_5081_),
    .Y(_3974_)
);

OAI21X1 _15109_ (
    .A(_4899__bF$buf6),
    .B(_5051__bF$buf5),
    .C(\datapath.registers.838[15] [29]),
    .Y(_5082_)
);

OAI21X1 _15110_ (
    .A(_4857__bF$buf3),
    .B(_5052__bF$buf0),
    .C(_5082_),
    .Y(_3975_)
);

OAI21X1 _15111_ (
    .A(_4899__bF$buf5),
    .B(_5051__bF$buf4),
    .C(\datapath.registers.838[15] [30]),
    .Y(_5083_)
);

OAI21X1 _15112_ (
    .A(_4859__bF$buf3),
    .B(_5052__bF$buf4),
    .C(_5083_),
    .Y(_3977_)
);

OAI21X1 _15113_ (
    .A(_4899__bF$buf4),
    .B(_5051__bF$buf3),
    .C(\datapath.registers.838[15] [31]),
    .Y(_5084_)
);

OAI21X1 _15114_ (
    .A(_4861__bF$buf3),
    .B(_5052__bF$buf3),
    .C(_5084_),
    .Y(_3978_)
);

NOR2X1 _15115_ (
    .A(_4934__bF$buf8),
    .B(_5051__bF$buf2),
    .Y(_5085_)
);

NOR2X1 _15116_ (
    .A(\datapath.registers.838[14] [0]),
    .B(_5085__bF$buf7),
    .Y(_5086_)
);

AOI21X1 _15117_ (
    .A(_4786__bF$buf2),
    .B(_5085__bF$buf6),
    .C(_5086_),
    .Y(_3922_)
);

NOR2X1 _15118_ (
    .A(\datapath.registers.838[14] [1]),
    .B(_5085__bF$buf5),
    .Y(_5087_)
);

AOI21X1 _15119_ (
    .A(_4801__bF$buf2),
    .B(_5085__bF$buf4),
    .C(_5087_),
    .Y(_3933_)
);

NOR2X1 _15120_ (
    .A(\datapath.registers.838[14] [2]),
    .B(_5085__bF$buf3),
    .Y(_5088_)
);

AOI21X1 _15121_ (
    .A(_4803__bF$buf2),
    .B(_5085__bF$buf2),
    .C(_5088_),
    .Y(_3944_)
);

NOR2X1 _15122_ (
    .A(\datapath.registers.838[14] [3]),
    .B(_5085__bF$buf1),
    .Y(_5089_)
);

AOI21X1 _15123_ (
    .A(_4805__bF$buf3),
    .B(_5085__bF$buf0),
    .C(_5089_),
    .Y(_3947_)
);

NOR2X1 _15124_ (
    .A(\datapath.registers.838[14] [4]),
    .B(_5085__bF$buf7),
    .Y(_5090_)
);

AOI21X1 _15125_ (
    .A(_4807__bF$buf3),
    .B(_5085__bF$buf6),
    .C(_5090_),
    .Y(_3948_)
);

NOR2X1 _15126_ (
    .A(\datapath.registers.838[14] [5]),
    .B(_5085__bF$buf5),
    .Y(_5091_)
);

AOI21X1 _15127_ (
    .A(_4809__bF$buf3),
    .B(_5085__bF$buf4),
    .C(_5091_),
    .Y(_3949_)
);

NOR2X1 _15128_ (
    .A(\datapath.registers.838[14] [6]),
    .B(_5085__bF$buf3),
    .Y(_5092_)
);

AOI21X1 _15129_ (
    .A(_4811__bF$buf3),
    .B(_5085__bF$buf2),
    .C(_5092_),
    .Y(_3950_)
);

NOR2X1 _15130_ (
    .A(\datapath.registers.838[14] [7]),
    .B(_5085__bF$buf1),
    .Y(_5093_)
);

AOI21X1 _15131_ (
    .A(_4813__bF$buf2),
    .B(_5085__bF$buf0),
    .C(_5093_),
    .Y(_3951_)
);

NOR2X1 _15132_ (
    .A(\datapath.registers.838[14] [8]),
    .B(_5085__bF$buf7),
    .Y(_5094_)
);

AOI21X1 _15133_ (
    .A(_4815__bF$buf2),
    .B(_5085__bF$buf6),
    .C(_5094_),
    .Y(_3952_)
);

NOR2X1 _15134_ (
    .A(\datapath.registers.838[14] [9]),
    .B(_5085__bF$buf5),
    .Y(_5095_)
);

AOI21X1 _15135_ (
    .A(_4817__bF$buf3),
    .B(_5085__bF$buf4),
    .C(_5095_),
    .Y(_3953_)
);

NOR2X1 _15136_ (
    .A(\datapath.registers.838[14] [10]),
    .B(_5085__bF$buf3),
    .Y(_5096_)
);

AOI21X1 _15137_ (
    .A(_4819__bF$buf3),
    .B(_5085__bF$buf2),
    .C(_5096_),
    .Y(_3923_)
);

NOR2X1 _15138_ (
    .A(\datapath.registers.838[14] [11]),
    .B(_5085__bF$buf1),
    .Y(_5097_)
);

AOI21X1 _15139_ (
    .A(_4821__bF$buf2),
    .B(_5085__bF$buf0),
    .C(_5097_),
    .Y(_3924_)
);

NOR2X1 _15140_ (
    .A(\datapath.registers.838[14] [12]),
    .B(_5085__bF$buf7),
    .Y(_5098_)
);

AOI21X1 _15141_ (
    .A(_4823__bF$buf2),
    .B(_5085__bF$buf6),
    .C(_5098_),
    .Y(_3925_)
);

NOR2X1 _15142_ (
    .A(\datapath.registers.838[14] [13]),
    .B(_5085__bF$buf5),
    .Y(_5099_)
);

AOI21X1 _15143_ (
    .A(_4825__bF$buf2),
    .B(_5085__bF$buf4),
    .C(_5099_),
    .Y(_3926_)
);

NOR2X1 _15144_ (
    .A(\datapath.registers.838[14] [14]),
    .B(_5085__bF$buf3),
    .Y(_5100_)
);

AOI21X1 _15145_ (
    .A(_4827__bF$buf2),
    .B(_5085__bF$buf2),
    .C(_5100_),
    .Y(_3927_)
);

NOR2X1 _15146_ (
    .A(\datapath.registers.838[14] [15]),
    .B(_5085__bF$buf1),
    .Y(_5101_)
);

AOI21X1 _15147_ (
    .A(_4829__bF$buf2),
    .B(_5085__bF$buf0),
    .C(_5101_),
    .Y(_3928_)
);

NOR2X1 _15148_ (
    .A(\datapath.registers.838[14] [16]),
    .B(_5085__bF$buf7),
    .Y(_5102_)
);

AOI21X1 _15149_ (
    .A(_4831__bF$buf2),
    .B(_5085__bF$buf6),
    .C(_5102_),
    .Y(_3929_)
);

NOR2X1 _15150_ (
    .A(\datapath.registers.838[14] [17]),
    .B(_5085__bF$buf5),
    .Y(_5103_)
);

AOI21X1 _15151_ (
    .A(_4833__bF$buf2),
    .B(_5085__bF$buf4),
    .C(_5103_),
    .Y(_3930_)
);

NOR2X1 _15152_ (
    .A(\datapath.registers.838[14] [18]),
    .B(_5085__bF$buf3),
    .Y(_5104_)
);

AOI21X1 _15153_ (
    .A(_4835__bF$buf2),
    .B(_5085__bF$buf2),
    .C(_5104_),
    .Y(_3931_)
);

NOR2X1 _15154_ (
    .A(\datapath.registers.838[14] [19]),
    .B(_5085__bF$buf1),
    .Y(_5105_)
);

AOI21X1 _15155_ (
    .A(_4837__bF$buf3),
    .B(_5085__bF$buf0),
    .C(_5105_),
    .Y(_3932_)
);

NOR2X1 _15156_ (
    .A(\datapath.registers.838[14] [20]),
    .B(_5085__bF$buf7),
    .Y(_5106_)
);

AOI21X1 _15157_ (
    .A(_4839__bF$buf2),
    .B(_5085__bF$buf6),
    .C(_5106_),
    .Y(_3934_)
);

NOR2X1 _15158_ (
    .A(\datapath.registers.838[14] [21]),
    .B(_5085__bF$buf5),
    .Y(_5107_)
);

AOI21X1 _15159_ (
    .A(_4841__bF$buf3),
    .B(_5085__bF$buf4),
    .C(_5107_),
    .Y(_3935_)
);

NOR2X1 _15160_ (
    .A(\datapath.registers.838[14] [22]),
    .B(_5085__bF$buf3),
    .Y(_5108_)
);

AOI21X1 _15161_ (
    .A(_4843__bF$buf3),
    .B(_5085__bF$buf2),
    .C(_5108_),
    .Y(_3936_)
);

NOR2X1 _15162_ (
    .A(\datapath.registers.838[14] [23]),
    .B(_5085__bF$buf1),
    .Y(_5109_)
);

AOI21X1 _15163_ (
    .A(_4845__bF$buf3),
    .B(_5085__bF$buf0),
    .C(_5109_),
    .Y(_3937_)
);

NOR2X1 _15164_ (
    .A(\datapath.registers.838[14] [24]),
    .B(_5085__bF$buf7),
    .Y(_5110_)
);

AOI21X1 _15165_ (
    .A(_4847__bF$buf3),
    .B(_5085__bF$buf6),
    .C(_5110_),
    .Y(_3938_)
);

NOR2X1 _15166_ (
    .A(\datapath.registers.838[14] [25]),
    .B(_5085__bF$buf5),
    .Y(_5111_)
);

AOI21X1 _15167_ (
    .A(_4849__bF$buf3),
    .B(_5085__bF$buf4),
    .C(_5111_),
    .Y(_3939_)
);

NOR2X1 _15168_ (
    .A(\datapath.registers.838[14] [26]),
    .B(_5085__bF$buf3),
    .Y(_5112_)
);

AOI21X1 _15169_ (
    .A(_4851__bF$buf2),
    .B(_5085__bF$buf2),
    .C(_5112_),
    .Y(_3940_)
);

NOR2X1 _15170_ (
    .A(\datapath.registers.838[14] [27]),
    .B(_5085__bF$buf1),
    .Y(_5113_)
);

AOI21X1 _15171_ (
    .A(_4853__bF$buf3),
    .B(_5085__bF$buf0),
    .C(_5113_),
    .Y(_3941_)
);

NOR2X1 _15172_ (
    .A(\datapath.registers.838[14] [28]),
    .B(_5085__bF$buf7),
    .Y(_5114_)
);

AOI21X1 _15173_ (
    .A(_4855__bF$buf2),
    .B(_5085__bF$buf6),
    .C(_5114_),
    .Y(_3942_)
);

NOR2X1 _15174_ (
    .A(\datapath.registers.838[14] [29]),
    .B(_5085__bF$buf5),
    .Y(_5115_)
);

AOI21X1 _15175_ (
    .A(_4857__bF$buf2),
    .B(_5085__bF$buf4),
    .C(_5115_),
    .Y(_3943_)
);

NOR2X1 _15176_ (
    .A(\datapath.registers.838[14] [30]),
    .B(_5085__bF$buf3),
    .Y(_5116_)
);

AOI21X1 _15177_ (
    .A(_4859__bF$buf2),
    .B(_5085__bF$buf2),
    .C(_5116_),
    .Y(_3945_)
);

NOR2X1 _15178_ (
    .A(\datapath.registers.838[14] [31]),
    .B(_5085__bF$buf1),
    .Y(_5117_)
);

AOI21X1 _15179_ (
    .A(_4861__bF$buf2),
    .B(_5085__bF$buf0),
    .C(_5117_),
    .Y(_3946_)
);

NOR2X1 _15180_ (
    .A(_4968__bF$buf8),
    .B(_5051__bF$buf1),
    .Y(_5118_)
);

NOR2X1 _15181_ (
    .A(\datapath.registers.838[13] [0]),
    .B(_5118__bF$buf7),
    .Y(_5119_)
);

AOI21X1 _15182_ (
    .A(_4786__bF$buf1),
    .B(_5118__bF$buf6),
    .C(_5119_),
    .Y(_3890_)
);

NOR2X1 _15183_ (
    .A(\datapath.registers.838[13] [1]),
    .B(_5118__bF$buf5),
    .Y(_5120_)
);

AOI21X1 _15184_ (
    .A(_4801__bF$buf1),
    .B(_5118__bF$buf4),
    .C(_5120_),
    .Y(_3901_)
);

NOR2X1 _15185_ (
    .A(\datapath.registers.838[13] [2]),
    .B(_5118__bF$buf3),
    .Y(_5121_)
);

AOI21X1 _15186_ (
    .A(_4803__bF$buf1),
    .B(_5118__bF$buf2),
    .C(_5121_),
    .Y(_3912_)
);

NOR2X1 _15187_ (
    .A(\datapath.registers.838[13] [3]),
    .B(_5118__bF$buf1),
    .Y(_5122_)
);

AOI21X1 _15188_ (
    .A(_4805__bF$buf2),
    .B(_5118__bF$buf0),
    .C(_5122_),
    .Y(_3915_)
);

NOR2X1 _15189_ (
    .A(\datapath.registers.838[13] [4]),
    .B(_5118__bF$buf7),
    .Y(_5123_)
);

AOI21X1 _15190_ (
    .A(_4807__bF$buf2),
    .B(_5118__bF$buf6),
    .C(_5123_),
    .Y(_3916_)
);

NOR2X1 _15191_ (
    .A(\datapath.registers.838[13] [5]),
    .B(_5118__bF$buf5),
    .Y(_5124_)
);

AOI21X1 _15192_ (
    .A(_4809__bF$buf2),
    .B(_5118__bF$buf4),
    .C(_5124_),
    .Y(_3917_)
);

NOR2X1 _15193_ (
    .A(\datapath.registers.838[13] [6]),
    .B(_5118__bF$buf3),
    .Y(_5125_)
);

AOI21X1 _15194_ (
    .A(_4811__bF$buf2),
    .B(_5118__bF$buf2),
    .C(_5125_),
    .Y(_3918_)
);

NOR2X1 _15195_ (
    .A(\datapath.registers.838[13] [7]),
    .B(_5118__bF$buf1),
    .Y(_5126_)
);

AOI21X1 _15196_ (
    .A(_4813__bF$buf1),
    .B(_5118__bF$buf0),
    .C(_5126_),
    .Y(_3919_)
);

NOR2X1 _15197_ (
    .A(\datapath.registers.838[13] [8]),
    .B(_5118__bF$buf7),
    .Y(_5127_)
);

AOI21X1 _15198_ (
    .A(_4815__bF$buf1),
    .B(_5118__bF$buf6),
    .C(_5127_),
    .Y(_3920_)
);

NOR2X1 _15199_ (
    .A(\datapath.registers.838[13] [9]),
    .B(_5118__bF$buf5),
    .Y(_5128_)
);

AOI21X1 _15200_ (
    .A(_4817__bF$buf2),
    .B(_5118__bF$buf4),
    .C(_5128_),
    .Y(_3921_)
);

NOR2X1 _15201_ (
    .A(\datapath.registers.838[13] [10]),
    .B(_5118__bF$buf3),
    .Y(_5129_)
);

AOI21X1 _15202_ (
    .A(_4819__bF$buf2),
    .B(_5118__bF$buf2),
    .C(_5129_),
    .Y(_3891_)
);

NOR2X1 _15203_ (
    .A(\datapath.registers.838[13] [11]),
    .B(_5118__bF$buf1),
    .Y(_5130_)
);

AOI21X1 _15204_ (
    .A(_4821__bF$buf1),
    .B(_5118__bF$buf0),
    .C(_5130_),
    .Y(_3892_)
);

NOR2X1 _15205_ (
    .A(\datapath.registers.838[13] [12]),
    .B(_5118__bF$buf7),
    .Y(_5131_)
);

AOI21X1 _15206_ (
    .A(_4823__bF$buf1),
    .B(_5118__bF$buf6),
    .C(_5131_),
    .Y(_3893_)
);

NOR2X1 _15207_ (
    .A(\datapath.registers.838[13] [13]),
    .B(_5118__bF$buf5),
    .Y(_5132_)
);

AOI21X1 _15208_ (
    .A(_4825__bF$buf1),
    .B(_5118__bF$buf4),
    .C(_5132_),
    .Y(_3894_)
);

NOR2X1 _15209_ (
    .A(\datapath.registers.838[13] [14]),
    .B(_5118__bF$buf3),
    .Y(_5133_)
);

AOI21X1 _15210_ (
    .A(_4827__bF$buf1),
    .B(_5118__bF$buf2),
    .C(_5133_),
    .Y(_3895_)
);

NOR2X1 _15211_ (
    .A(\datapath.registers.838[13] [15]),
    .B(_5118__bF$buf1),
    .Y(_5134_)
);

AOI21X1 _15212_ (
    .A(_4829__bF$buf1),
    .B(_5118__bF$buf0),
    .C(_5134_),
    .Y(_3896_)
);

NOR2X1 _15213_ (
    .A(\datapath.registers.838[13] [16]),
    .B(_5118__bF$buf7),
    .Y(_5135_)
);

AOI21X1 _15214_ (
    .A(_4831__bF$buf1),
    .B(_5118__bF$buf6),
    .C(_5135_),
    .Y(_3897_)
);

NOR2X1 _15215_ (
    .A(\datapath.registers.838[13] [17]),
    .B(_5118__bF$buf5),
    .Y(_5136_)
);

AOI21X1 _15216_ (
    .A(_4833__bF$buf1),
    .B(_5118__bF$buf4),
    .C(_5136_),
    .Y(_3898_)
);

NOR2X1 _15217_ (
    .A(\datapath.registers.838[13] [18]),
    .B(_5118__bF$buf3),
    .Y(_5137_)
);

AOI21X1 _15218_ (
    .A(_4835__bF$buf1),
    .B(_5118__bF$buf2),
    .C(_5137_),
    .Y(_3899_)
);

NOR2X1 _15219_ (
    .A(\datapath.registers.838[13] [19]),
    .B(_5118__bF$buf1),
    .Y(_5138_)
);

AOI21X1 _15220_ (
    .A(_4837__bF$buf2),
    .B(_5118__bF$buf0),
    .C(_5138_),
    .Y(_3900_)
);

NOR2X1 _15221_ (
    .A(\datapath.registers.838[13] [20]),
    .B(_5118__bF$buf7),
    .Y(_5139_)
);

AOI21X1 _15222_ (
    .A(_4839__bF$buf1),
    .B(_5118__bF$buf6),
    .C(_5139_),
    .Y(_3902_)
);

NOR2X1 _15223_ (
    .A(\datapath.registers.838[13] [21]),
    .B(_5118__bF$buf5),
    .Y(_5140_)
);

AOI21X1 _15224_ (
    .A(_4841__bF$buf2),
    .B(_5118__bF$buf4),
    .C(_5140_),
    .Y(_3903_)
);

NOR2X1 _15225_ (
    .A(\datapath.registers.838[13] [22]),
    .B(_5118__bF$buf3),
    .Y(_5141_)
);

AOI21X1 _15226_ (
    .A(_4843__bF$buf2),
    .B(_5118__bF$buf2),
    .C(_5141_),
    .Y(_3904_)
);

NOR2X1 _15227_ (
    .A(\datapath.registers.838[13] [23]),
    .B(_5118__bF$buf1),
    .Y(_5142_)
);

AOI21X1 _15228_ (
    .A(_4845__bF$buf2),
    .B(_5118__bF$buf0),
    .C(_5142_),
    .Y(_3905_)
);

NOR2X1 _15229_ (
    .A(\datapath.registers.838[13] [24]),
    .B(_5118__bF$buf7),
    .Y(_5143_)
);

AOI21X1 _15230_ (
    .A(_4847__bF$buf2),
    .B(_5118__bF$buf6),
    .C(_5143_),
    .Y(_3906_)
);

NOR2X1 _15231_ (
    .A(\datapath.registers.838[13] [25]),
    .B(_5118__bF$buf5),
    .Y(_5144_)
);

AOI21X1 _15232_ (
    .A(_4849__bF$buf2),
    .B(_5118__bF$buf4),
    .C(_5144_),
    .Y(_3907_)
);

NOR2X1 _15233_ (
    .A(\datapath.registers.838[13] [26]),
    .B(_5118__bF$buf3),
    .Y(_5145_)
);

AOI21X1 _15234_ (
    .A(_4851__bF$buf1),
    .B(_5118__bF$buf2),
    .C(_5145_),
    .Y(_3908_)
);

NOR2X1 _15235_ (
    .A(\datapath.registers.838[13] [27]),
    .B(_5118__bF$buf1),
    .Y(_5146_)
);

AOI21X1 _15236_ (
    .A(_4853__bF$buf2),
    .B(_5118__bF$buf0),
    .C(_5146_),
    .Y(_3909_)
);

NOR2X1 _15237_ (
    .A(\datapath.registers.838[13] [28]),
    .B(_5118__bF$buf7),
    .Y(_5147_)
);

AOI21X1 _15238_ (
    .A(_4855__bF$buf1),
    .B(_5118__bF$buf6),
    .C(_5147_),
    .Y(_3910_)
);

NOR2X1 _15239_ (
    .A(\datapath.registers.838[13] [29]),
    .B(_5118__bF$buf5),
    .Y(_5148_)
);

AOI21X1 _15240_ (
    .A(_4857__bF$buf1),
    .B(_5118__bF$buf4),
    .C(_5148_),
    .Y(_3911_)
);

NOR2X1 _15241_ (
    .A(\datapath.registers.838[13] [30]),
    .B(_5118__bF$buf3),
    .Y(_5149_)
);

AOI21X1 _15242_ (
    .A(_4859__bF$buf1),
    .B(_5118__bF$buf2),
    .C(_5149_),
    .Y(_3913_)
);

NOR2X1 _15243_ (
    .A(\datapath.registers.838[13] [31]),
    .B(_5118__bF$buf1),
    .Y(_5150_)
);

AOI21X1 _15244_ (
    .A(_4861__bF$buf1),
    .B(_5118__bF$buf0),
    .C(_5150_),
    .Y(_3914_)
);

NOR2X1 _15245_ (
    .A(_4790_),
    .B(_5051__bF$buf0),
    .Y(_5151_)
);

NAND2X1 _15246_ (
    .A(_5015_),
    .B(_5151_),
    .Y(_5152_)
);

NAND2X1 _15247_ (
    .A(\datapath.registers.838[12] [0]),
    .B(_5152__bF$buf7),
    .Y(_5153_)
);

OAI21X1 _15248_ (
    .A(_4786__bF$buf0),
    .B(_5152__bF$buf6),
    .C(_5153_),
    .Y(_3858_)
);

NAND2X1 _15249_ (
    .A(\datapath.registers.838[12] [1]),
    .B(_5152__bF$buf5),
    .Y(_5154_)
);

OAI21X1 _15250_ (
    .A(_4801__bF$buf0),
    .B(_5152__bF$buf4),
    .C(_5154_),
    .Y(_3869_)
);

NAND2X1 _15251_ (
    .A(\datapath.registers.838[12] [2]),
    .B(_5152__bF$buf3),
    .Y(_5155_)
);

OAI21X1 _15252_ (
    .A(_4803__bF$buf0),
    .B(_5152__bF$buf2),
    .C(_5155_),
    .Y(_3880_)
);

NAND2X1 _15253_ (
    .A(\datapath.registers.838[12] [3]),
    .B(_5152__bF$buf1),
    .Y(_5156_)
);

OAI21X1 _15254_ (
    .A(_4805__bF$buf1),
    .B(_5152__bF$buf0),
    .C(_5156_),
    .Y(_3883_)
);

NAND2X1 _15255_ (
    .A(\datapath.registers.838[12] [4]),
    .B(_5152__bF$buf7),
    .Y(_5157_)
);

OAI21X1 _15256_ (
    .A(_4807__bF$buf1),
    .B(_5152__bF$buf6),
    .C(_5157_),
    .Y(_3884_)
);

NAND2X1 _15257_ (
    .A(\datapath.registers.838[12] [5]),
    .B(_5152__bF$buf5),
    .Y(_5158_)
);

OAI21X1 _15258_ (
    .A(_4809__bF$buf1),
    .B(_5152__bF$buf4),
    .C(_5158_),
    .Y(_3885_)
);

NAND2X1 _15259_ (
    .A(\datapath.registers.838[12] [6]),
    .B(_5152__bF$buf3),
    .Y(_5159_)
);

OAI21X1 _15260_ (
    .A(_4811__bF$buf1),
    .B(_5152__bF$buf2),
    .C(_5159_),
    .Y(_3886_)
);

NAND2X1 _15261_ (
    .A(\datapath.registers.838[12] [7]),
    .B(_5152__bF$buf1),
    .Y(_5160_)
);

OAI21X1 _15262_ (
    .A(_4813__bF$buf0),
    .B(_5152__bF$buf0),
    .C(_5160_),
    .Y(_3887_)
);

NAND2X1 _15263_ (
    .A(\datapath.registers.838[12] [8]),
    .B(_5152__bF$buf7),
    .Y(_5161_)
);

OAI21X1 _15264_ (
    .A(_4815__bF$buf0),
    .B(_5152__bF$buf6),
    .C(_5161_),
    .Y(_3888_)
);

NAND2X1 _15265_ (
    .A(\datapath.registers.838[12] [9]),
    .B(_5152__bF$buf5),
    .Y(_5162_)
);

OAI21X1 _15266_ (
    .A(_4817__bF$buf1),
    .B(_5152__bF$buf4),
    .C(_5162_),
    .Y(_3889_)
);

NAND2X1 _15267_ (
    .A(\datapath.registers.838[12] [10]),
    .B(_5152__bF$buf3),
    .Y(_5163_)
);

OAI21X1 _15268_ (
    .A(_4819__bF$buf1),
    .B(_5152__bF$buf2),
    .C(_5163_),
    .Y(_3859_)
);

NAND2X1 _15269_ (
    .A(\datapath.registers.838[12] [11]),
    .B(_5152__bF$buf1),
    .Y(_5164_)
);

OAI21X1 _15270_ (
    .A(_4821__bF$buf0),
    .B(_5152__bF$buf0),
    .C(_5164_),
    .Y(_3860_)
);

NAND2X1 _15271_ (
    .A(\datapath.registers.838[12] [12]),
    .B(_5152__bF$buf7),
    .Y(_5165_)
);

OAI21X1 _15272_ (
    .A(_4823__bF$buf0),
    .B(_5152__bF$buf6),
    .C(_5165_),
    .Y(_3861_)
);

NAND2X1 _15273_ (
    .A(\datapath.registers.838[12] [13]),
    .B(_5152__bF$buf5),
    .Y(_5166_)
);

OAI21X1 _15274_ (
    .A(_4825__bF$buf0),
    .B(_5152__bF$buf4),
    .C(_5166_),
    .Y(_3862_)
);

NAND2X1 _15275_ (
    .A(\datapath.registers.838[12] [14]),
    .B(_5152__bF$buf3),
    .Y(_5167_)
);

OAI21X1 _15276_ (
    .A(_4827__bF$buf0),
    .B(_5152__bF$buf2),
    .C(_5167_),
    .Y(_3863_)
);

NAND2X1 _15277_ (
    .A(\datapath.registers.838[12] [15]),
    .B(_5152__bF$buf1),
    .Y(_5168_)
);

OAI21X1 _15278_ (
    .A(_4829__bF$buf0),
    .B(_5152__bF$buf0),
    .C(_5168_),
    .Y(_3864_)
);

NAND2X1 _15279_ (
    .A(\datapath.registers.838[12] [16]),
    .B(_5152__bF$buf7),
    .Y(_5169_)
);

OAI21X1 _15280_ (
    .A(_4831__bF$buf0),
    .B(_5152__bF$buf6),
    .C(_5169_),
    .Y(_3865_)
);

NAND2X1 _15281_ (
    .A(\datapath.registers.838[12] [17]),
    .B(_5152__bF$buf5),
    .Y(_5170_)
);

OAI21X1 _15282_ (
    .A(_4833__bF$buf0),
    .B(_5152__bF$buf4),
    .C(_5170_),
    .Y(_3866_)
);

NAND2X1 _15283_ (
    .A(\datapath.registers.838[12] [18]),
    .B(_5152__bF$buf3),
    .Y(_5171_)
);

OAI21X1 _15284_ (
    .A(_4835__bF$buf0),
    .B(_5152__bF$buf2),
    .C(_5171_),
    .Y(_3867_)
);

NAND2X1 _15285_ (
    .A(\datapath.registers.838[12] [19]),
    .B(_5152__bF$buf1),
    .Y(_5172_)
);

OAI21X1 _15286_ (
    .A(_4837__bF$buf1),
    .B(_5152__bF$buf0),
    .C(_5172_),
    .Y(_3868_)
);

NAND2X1 _15287_ (
    .A(\datapath.registers.838[12] [20]),
    .B(_5152__bF$buf7),
    .Y(_5173_)
);

OAI21X1 _15288_ (
    .A(_4839__bF$buf0),
    .B(_5152__bF$buf6),
    .C(_5173_),
    .Y(_3870_)
);

NAND2X1 _15289_ (
    .A(\datapath.registers.838[12] [21]),
    .B(_5152__bF$buf5),
    .Y(_5174_)
);

OAI21X1 _15290_ (
    .A(_4841__bF$buf1),
    .B(_5152__bF$buf4),
    .C(_5174_),
    .Y(_3871_)
);

NAND2X1 _15291_ (
    .A(\datapath.registers.838[12] [22]),
    .B(_5152__bF$buf3),
    .Y(_5175_)
);

OAI21X1 _15292_ (
    .A(_4843__bF$buf1),
    .B(_5152__bF$buf2),
    .C(_5175_),
    .Y(_3872_)
);

NAND2X1 _15293_ (
    .A(\datapath.registers.838[12] [23]),
    .B(_5152__bF$buf1),
    .Y(_5176_)
);

OAI21X1 _15294_ (
    .A(_4845__bF$buf1),
    .B(_5152__bF$buf0),
    .C(_5176_),
    .Y(_3873_)
);

NAND2X1 _15295_ (
    .A(\datapath.registers.838[12] [24]),
    .B(_5152__bF$buf7),
    .Y(_5177_)
);

OAI21X1 _15296_ (
    .A(_4847__bF$buf1),
    .B(_5152__bF$buf6),
    .C(_5177_),
    .Y(_3874_)
);

NAND2X1 _15297_ (
    .A(\datapath.registers.838[12] [25]),
    .B(_5152__bF$buf5),
    .Y(_5178_)
);

OAI21X1 _15298_ (
    .A(_4849__bF$buf1),
    .B(_5152__bF$buf4),
    .C(_5178_),
    .Y(_3875_)
);

NAND2X1 _15299_ (
    .A(\datapath.registers.838[12] [26]),
    .B(_5152__bF$buf3),
    .Y(_5179_)
);

OAI21X1 _15300_ (
    .A(_4851__bF$buf0),
    .B(_5152__bF$buf2),
    .C(_5179_),
    .Y(_3876_)
);

NAND2X1 _15301_ (
    .A(\datapath.registers.838[12] [27]),
    .B(_5152__bF$buf1),
    .Y(_5180_)
);

OAI21X1 _15302_ (
    .A(_4853__bF$buf1),
    .B(_5152__bF$buf0),
    .C(_5180_),
    .Y(_3877_)
);

NAND2X1 _15303_ (
    .A(\datapath.registers.838[12] [28]),
    .B(_5152__bF$buf7),
    .Y(_5181_)
);

OAI21X1 _15304_ (
    .A(_4855__bF$buf0),
    .B(_5152__bF$buf6),
    .C(_5181_),
    .Y(_3878_)
);

NAND2X1 _15305_ (
    .A(\datapath.registers.838[12] [29]),
    .B(_5152__bF$buf5),
    .Y(_5182_)
);

OAI21X1 _15306_ (
    .A(_4857__bF$buf0),
    .B(_5152__bF$buf4),
    .C(_5182_),
    .Y(_3879_)
);

NAND2X1 _15307_ (
    .A(\datapath.registers.838[12] [30]),
    .B(_5152__bF$buf3),
    .Y(_5183_)
);

OAI21X1 _15308_ (
    .A(_4859__bF$buf0),
    .B(_5152__bF$buf2),
    .C(_5183_),
    .Y(_3881_)
);

NAND2X1 _15309_ (
    .A(\datapath.registers.838[12] [31]),
    .B(_5152__bF$buf1),
    .Y(_5184_)
);

OAI21X1 _15310_ (
    .A(_4861__bF$buf0),
    .B(_5152__bF$buf0),
    .C(_5184_),
    .Y(_3882_)
);

OR2X2 _15311_ (
    .A(_5050_),
    .B(\datapath.wbinstr [9]),
    .Y(_5185_)
);

OR2X2 _15312_ (
    .A(_5185__bF$buf5),
    .B(_4899__bF$buf3),
    .Y(_5186_)
);

OAI21X1 _15313_ (
    .A(_4899__bF$buf2),
    .B(_5185__bF$buf4),
    .C(\datapath.registers.838[11] [0]),
    .Y(_5187_)
);

OAI21X1 _15314_ (
    .A(_4786__bF$buf4),
    .B(_5186__bF$buf4),
    .C(_5187_),
    .Y(_3826_)
);

OAI21X1 _15315_ (
    .A(_4899__bF$buf1),
    .B(_5185__bF$buf3),
    .C(\datapath.registers.838[11] [1]),
    .Y(_5188_)
);

OAI21X1 _15316_ (
    .A(_4801__bF$buf4),
    .B(_5186__bF$buf3),
    .C(_5188_),
    .Y(_3837_)
);

OAI21X1 _15317_ (
    .A(_4899__bF$buf0),
    .B(_5185__bF$buf2),
    .C(\datapath.registers.838[11] [2]),
    .Y(_5189_)
);

OAI21X1 _15318_ (
    .A(_4803__bF$buf4),
    .B(_5186__bF$buf2),
    .C(_5189_),
    .Y(_3848_)
);

OAI21X1 _15319_ (
    .A(_4899__bF$buf13),
    .B(_5185__bF$buf1),
    .C(\datapath.registers.838[11] [3]),
    .Y(_5190_)
);

OAI21X1 _15320_ (
    .A(_4805__bF$buf0),
    .B(_5186__bF$buf1),
    .C(_5190_),
    .Y(_3851_)
);

OAI21X1 _15321_ (
    .A(_4899__bF$buf12),
    .B(_5185__bF$buf0),
    .C(\datapath.registers.838[11] [4]),
    .Y(_5191_)
);

OAI21X1 _15322_ (
    .A(_4807__bF$buf0),
    .B(_5186__bF$buf0),
    .C(_5191_),
    .Y(_3852_)
);

OAI21X1 _15323_ (
    .A(_4899__bF$buf11),
    .B(_5185__bF$buf5),
    .C(\datapath.registers.838[11] [5]),
    .Y(_5192_)
);

OAI21X1 _15324_ (
    .A(_4809__bF$buf0),
    .B(_5186__bF$buf4),
    .C(_5192_),
    .Y(_3853_)
);

OAI21X1 _15325_ (
    .A(_4899__bF$buf10),
    .B(_5185__bF$buf4),
    .C(\datapath.registers.838[11] [6]),
    .Y(_5193_)
);

OAI21X1 _15326_ (
    .A(_4811__bF$buf0),
    .B(_5186__bF$buf3),
    .C(_5193_),
    .Y(_3854_)
);

OAI21X1 _15327_ (
    .A(_4899__bF$buf9),
    .B(_5185__bF$buf3),
    .C(\datapath.registers.838[11] [7]),
    .Y(_5194_)
);

OAI21X1 _15328_ (
    .A(_4813__bF$buf4),
    .B(_5186__bF$buf2),
    .C(_5194_),
    .Y(_3855_)
);

OAI21X1 _15329_ (
    .A(_4899__bF$buf8),
    .B(_5185__bF$buf2),
    .C(\datapath.registers.838[11] [8]),
    .Y(_5195_)
);

OAI21X1 _15330_ (
    .A(_4815__bF$buf4),
    .B(_5186__bF$buf1),
    .C(_5195_),
    .Y(_3856_)
);

OAI21X1 _15331_ (
    .A(_4899__bF$buf7),
    .B(_5185__bF$buf1),
    .C(\datapath.registers.838[11] [9]),
    .Y(_5196_)
);

OAI21X1 _15332_ (
    .A(_4817__bF$buf0),
    .B(_5186__bF$buf0),
    .C(_5196_),
    .Y(_3857_)
);

OAI21X1 _15333_ (
    .A(_4899__bF$buf6),
    .B(_5185__bF$buf0),
    .C(\datapath.registers.838[11] [10]),
    .Y(_5197_)
);

OAI21X1 _15334_ (
    .A(_4819__bF$buf0),
    .B(_5186__bF$buf4),
    .C(_5197_),
    .Y(_3827_)
);

OAI21X1 _15335_ (
    .A(_4899__bF$buf5),
    .B(_5185__bF$buf5),
    .C(\datapath.registers.838[11] [11]),
    .Y(_5198_)
);

OAI21X1 _15336_ (
    .A(_4821__bF$buf4),
    .B(_5186__bF$buf3),
    .C(_5198_),
    .Y(_3828_)
);

OAI21X1 _15337_ (
    .A(_4899__bF$buf4),
    .B(_5185__bF$buf4),
    .C(\datapath.registers.838[11] [12]),
    .Y(_5199_)
);

OAI21X1 _15338_ (
    .A(_4823__bF$buf4),
    .B(_5186__bF$buf2),
    .C(_5199_),
    .Y(_3829_)
);

OAI21X1 _15339_ (
    .A(_4899__bF$buf3),
    .B(_5185__bF$buf3),
    .C(\datapath.registers.838[11] [13]),
    .Y(_5200_)
);

OAI21X1 _15340_ (
    .A(_4825__bF$buf4),
    .B(_5186__bF$buf1),
    .C(_5200_),
    .Y(_3830_)
);

OAI21X1 _15341_ (
    .A(_4899__bF$buf2),
    .B(_5185__bF$buf2),
    .C(\datapath.registers.838[11] [14]),
    .Y(_5201_)
);

OAI21X1 _15342_ (
    .A(_4827__bF$buf4),
    .B(_5186__bF$buf0),
    .C(_5201_),
    .Y(_3831_)
);

OAI21X1 _15343_ (
    .A(_4899__bF$buf1),
    .B(_5185__bF$buf1),
    .C(\datapath.registers.838[11] [15]),
    .Y(_5202_)
);

OAI21X1 _15344_ (
    .A(_4829__bF$buf4),
    .B(_5186__bF$buf4),
    .C(_5202_),
    .Y(_3832_)
);

OAI21X1 _15345_ (
    .A(_4899__bF$buf0),
    .B(_5185__bF$buf0),
    .C(\datapath.registers.838[11] [16]),
    .Y(_5203_)
);

OAI21X1 _15346_ (
    .A(_4831__bF$buf4),
    .B(_5186__bF$buf3),
    .C(_5203_),
    .Y(_3833_)
);

OAI21X1 _15347_ (
    .A(_4899__bF$buf13),
    .B(_5185__bF$buf5),
    .C(\datapath.registers.838[11] [17]),
    .Y(_5204_)
);

OAI21X1 _15348_ (
    .A(_4833__bF$buf4),
    .B(_5186__bF$buf2),
    .C(_5204_),
    .Y(_3834_)
);

OAI21X1 _15349_ (
    .A(_4899__bF$buf12),
    .B(_5185__bF$buf4),
    .C(\datapath.registers.838[11] [18]),
    .Y(_5205_)
);

OAI21X1 _15350_ (
    .A(_4835__bF$buf4),
    .B(_5186__bF$buf1),
    .C(_5205_),
    .Y(_3835_)
);

OAI21X1 _15351_ (
    .A(_4899__bF$buf11),
    .B(_5185__bF$buf3),
    .C(\datapath.registers.838[11] [19]),
    .Y(_5206_)
);

OAI21X1 _15352_ (
    .A(_4837__bF$buf0),
    .B(_5186__bF$buf0),
    .C(_5206_),
    .Y(_3836_)
);

OAI21X1 _15353_ (
    .A(_4899__bF$buf10),
    .B(_5185__bF$buf2),
    .C(\datapath.registers.838[11] [20]),
    .Y(_5207_)
);

OAI21X1 _15354_ (
    .A(_4839__bF$buf4),
    .B(_5186__bF$buf4),
    .C(_5207_),
    .Y(_3838_)
);

OAI21X1 _15355_ (
    .A(_4899__bF$buf9),
    .B(_5185__bF$buf1),
    .C(\datapath.registers.838[11] [21]),
    .Y(_5208_)
);

OAI21X1 _15356_ (
    .A(_4841__bF$buf0),
    .B(_5186__bF$buf3),
    .C(_5208_),
    .Y(_3839_)
);

OAI21X1 _15357_ (
    .A(_4899__bF$buf8),
    .B(_5185__bF$buf0),
    .C(\datapath.registers.838[11] [22]),
    .Y(_5209_)
);

OAI21X1 _15358_ (
    .A(_4843__bF$buf0),
    .B(_5186__bF$buf2),
    .C(_5209_),
    .Y(_3840_)
);

OAI21X1 _15359_ (
    .A(_4899__bF$buf7),
    .B(_5185__bF$buf5),
    .C(\datapath.registers.838[11] [23]),
    .Y(_5210_)
);

OAI21X1 _15360_ (
    .A(_4845__bF$buf0),
    .B(_5186__bF$buf1),
    .C(_5210_),
    .Y(_3841_)
);

OAI21X1 _15361_ (
    .A(_4899__bF$buf6),
    .B(_5185__bF$buf4),
    .C(\datapath.registers.838[11] [24]),
    .Y(_5211_)
);

OAI21X1 _15362_ (
    .A(_4847__bF$buf0),
    .B(_5186__bF$buf0),
    .C(_5211_),
    .Y(_3842_)
);

OAI21X1 _15363_ (
    .A(_4899__bF$buf5),
    .B(_5185__bF$buf3),
    .C(\datapath.registers.838[11] [25]),
    .Y(_5212_)
);

OAI21X1 _15364_ (
    .A(_4849__bF$buf0),
    .B(_5186__bF$buf4),
    .C(_5212_),
    .Y(_3843_)
);

OAI21X1 _15365_ (
    .A(_4899__bF$buf4),
    .B(_5185__bF$buf2),
    .C(\datapath.registers.838[11] [26]),
    .Y(_5213_)
);

OAI21X1 _15366_ (
    .A(_4851__bF$buf4),
    .B(_5186__bF$buf3),
    .C(_5213_),
    .Y(_3844_)
);

OAI21X1 _15367_ (
    .A(_4899__bF$buf3),
    .B(_5185__bF$buf1),
    .C(\datapath.registers.838[11] [27]),
    .Y(_5214_)
);

OAI21X1 _15368_ (
    .A(_4853__bF$buf0),
    .B(_5186__bF$buf2),
    .C(_5214_),
    .Y(_3845_)
);

OAI21X1 _15369_ (
    .A(_4899__bF$buf2),
    .B(_5185__bF$buf0),
    .C(\datapath.registers.838[11] [28]),
    .Y(_5215_)
);

OAI21X1 _15370_ (
    .A(_4855__bF$buf4),
    .B(_5186__bF$buf1),
    .C(_5215_),
    .Y(_3846_)
);

OAI21X1 _15371_ (
    .A(_4899__bF$buf1),
    .B(_5185__bF$buf5),
    .C(\datapath.registers.838[11] [29]),
    .Y(_5216_)
);

OAI21X1 _15372_ (
    .A(_4857__bF$buf4),
    .B(_5186__bF$buf0),
    .C(_5216_),
    .Y(_3847_)
);

OAI21X1 _15373_ (
    .A(_4899__bF$buf0),
    .B(_5185__bF$buf4),
    .C(\datapath.registers.838[11] [30]),
    .Y(_5217_)
);

OAI21X1 _15374_ (
    .A(_4859__bF$buf4),
    .B(_5186__bF$buf4),
    .C(_5217_),
    .Y(_3849_)
);

OAI21X1 _15375_ (
    .A(_4899__bF$buf13),
    .B(_5185__bF$buf3),
    .C(\datapath.registers.838[11] [31]),
    .Y(_5218_)
);

OAI21X1 _15376_ (
    .A(_4861__bF$buf4),
    .B(_5186__bF$buf3),
    .C(_5218_),
    .Y(_3850_)
);

INVX1 _15377_ (
    .A(\datapath.registers.838[10] [0]),
    .Y(_5219_)
);

NOR2X1 _15378_ (
    .A(_4934__bF$buf7),
    .B(_5185__bF$buf2),
    .Y(_5220_)
);

NAND2X1 _15379_ (
    .A(\datapath.rd [0]),
    .B(_5220__bF$buf7),
    .Y(_5221_)
);

OAI21X1 _15380_ (
    .A(_5219_),
    .B(_5220__bF$buf6),
    .C(_5221_),
    .Y(_3794_)
);

NOR2X1 _15381_ (
    .A(\datapath.registers.838[10] [1]),
    .B(_5220__bF$buf5),
    .Y(_5222_)
);

AOI21X1 _15382_ (
    .A(_4801__bF$buf3),
    .B(_5220__bF$buf4),
    .C(_5222_),
    .Y(_3805_)
);

INVX1 _15383_ (
    .A(\datapath.registers.838[10] [2]),
    .Y(_5223_)
);

NAND2X1 _15384_ (
    .A(\datapath.rd [2]),
    .B(_5220__bF$buf3),
    .Y(_5224_)
);

OAI21X1 _15385_ (
    .A(_5223_),
    .B(_5220__bF$buf2),
    .C(_5224_),
    .Y(_3816_)
);

INVX1 _15386_ (
    .A(\datapath.registers.838[10] [3]),
    .Y(_5225_)
);

NAND2X1 _15387_ (
    .A(\datapath.rd [3]),
    .B(_5220__bF$buf1),
    .Y(_5226_)
);

OAI21X1 _15388_ (
    .A(_5225_),
    .B(_5220__bF$buf0),
    .C(_5226_),
    .Y(_3819_)
);

NOR2X1 _15389_ (
    .A(\datapath.registers.838[10] [4]),
    .B(_5220__bF$buf7),
    .Y(_5227_)
);

AOI21X1 _15390_ (
    .A(_4807__bF$buf4),
    .B(_5220__bF$buf6),
    .C(_5227_),
    .Y(_3820_)
);

NOR2X1 _15391_ (
    .A(\datapath.registers.838[10] [5]),
    .B(_5220__bF$buf5),
    .Y(_5228_)
);

AOI21X1 _15392_ (
    .A(_4809__bF$buf4),
    .B(_5220__bF$buf4),
    .C(_5228_),
    .Y(_3821_)
);

INVX1 _15393_ (
    .A(\datapath.registers.838[10] [6]),
    .Y(_5229_)
);

NAND2X1 _15394_ (
    .A(\datapath.rd [6]),
    .B(_5220__bF$buf3),
    .Y(_5230_)
);

OAI21X1 _15395_ (
    .A(_5229_),
    .B(_5220__bF$buf2),
    .C(_5230_),
    .Y(_3822_)
);

NOR2X1 _15396_ (
    .A(\datapath.registers.838[10] [7]),
    .B(_5220__bF$buf1),
    .Y(_5231_)
);

AOI21X1 _15397_ (
    .A(_4813__bF$buf3),
    .B(_5220__bF$buf0),
    .C(_5231_),
    .Y(_3823_)
);

NOR2X1 _15398_ (
    .A(\datapath.registers.838[10] [8]),
    .B(_5220__bF$buf7),
    .Y(_5232_)
);

AOI21X1 _15399_ (
    .A(_4815__bF$buf3),
    .B(_5220__bF$buf6),
    .C(_5232_),
    .Y(_3824_)
);

INVX1 _15400_ (
    .A(\datapath.registers.838[10] [9]),
    .Y(_5233_)
);

NAND2X1 _15401_ (
    .A(\datapath.rd [9]),
    .B(_5220__bF$buf5),
    .Y(_5234_)
);

OAI21X1 _15402_ (
    .A(_5233_),
    .B(_5220__bF$buf4),
    .C(_5234_),
    .Y(_3825_)
);

NOR2X1 _15403_ (
    .A(\datapath.registers.838[10] [10]),
    .B(_5220__bF$buf3),
    .Y(_5235_)
);

AOI21X1 _15404_ (
    .A(_4819__bF$buf4),
    .B(_5220__bF$buf2),
    .C(_5235_),
    .Y(_3795_)
);

NOR2X1 _15405_ (
    .A(\datapath.registers.838[10] [11]),
    .B(_5220__bF$buf1),
    .Y(_5236_)
);

AOI21X1 _15406_ (
    .A(_4821__bF$buf3),
    .B(_5220__bF$buf0),
    .C(_5236_),
    .Y(_3796_)
);

INVX1 _15407_ (
    .A(\datapath.registers.838[10] [12]),
    .Y(_5237_)
);

NAND2X1 _15408_ (
    .A(\datapath.rd [12]),
    .B(_5220__bF$buf7),
    .Y(_5238_)
);

OAI21X1 _15409_ (
    .A(_5237_),
    .B(_5220__bF$buf6),
    .C(_5238_),
    .Y(_3797_)
);

NOR2X1 _15410_ (
    .A(\datapath.registers.838[10] [13]),
    .B(_5220__bF$buf5),
    .Y(_5239_)
);

AOI21X1 _15411_ (
    .A(_4825__bF$buf3),
    .B(_5220__bF$buf4),
    .C(_5239_),
    .Y(_3798_)
);

NOR2X1 _15412_ (
    .A(\datapath.registers.838[10] [14]),
    .B(_5220__bF$buf3),
    .Y(_5240_)
);

AOI21X1 _15413_ (
    .A(_4827__bF$buf3),
    .B(_5220__bF$buf2),
    .C(_5240_),
    .Y(_3799_)
);

NOR2X1 _15414_ (
    .A(\datapath.registers.838[10] [15]),
    .B(_5220__bF$buf1),
    .Y(_5241_)
);

AOI21X1 _15415_ (
    .A(_4829__bF$buf3),
    .B(_5220__bF$buf0),
    .C(_5241_),
    .Y(_3800_)
);

NOR2X1 _15416_ (
    .A(\datapath.registers.838[10] [16]),
    .B(_5220__bF$buf7),
    .Y(_5242_)
);

AOI21X1 _15417_ (
    .A(_4831__bF$buf3),
    .B(_5220__bF$buf6),
    .C(_5242_),
    .Y(_3801_)
);

INVX1 _15418_ (
    .A(\datapath.registers.838[10] [17]),
    .Y(_5243_)
);

NAND2X1 _15419_ (
    .A(\datapath.rd [17]),
    .B(_5220__bF$buf5),
    .Y(_5244_)
);

OAI21X1 _15420_ (
    .A(_5243_),
    .B(_5220__bF$buf4),
    .C(_5244_),
    .Y(_3802_)
);

INVX1 _15421_ (
    .A(\datapath.registers.838[10] [18]),
    .Y(_5245_)
);

NAND2X1 _15422_ (
    .A(\datapath.rd [18]),
    .B(_5220__bF$buf3),
    .Y(_5246_)
);

OAI21X1 _15423_ (
    .A(_5245_),
    .B(_5220__bF$buf2),
    .C(_5246_),
    .Y(_3803_)
);

INVX1 _15424_ (
    .A(\datapath.registers.838[10] [19]),
    .Y(_5247_)
);

NAND2X1 _15425_ (
    .A(\datapath.rd [19]),
    .B(_5220__bF$buf1),
    .Y(_5248_)
);

OAI21X1 _15426_ (
    .A(_5247_),
    .B(_5220__bF$buf0),
    .C(_5248_),
    .Y(_3804_)
);

NOR2X1 _15427_ (
    .A(\datapath.registers.838[10] [20]),
    .B(_5220__bF$buf7),
    .Y(_5249_)
);

AOI21X1 _15428_ (
    .A(_4839__bF$buf3),
    .B(_5220__bF$buf6),
    .C(_5249_),
    .Y(_3806_)
);

NOR2X1 _15429_ (
    .A(\datapath.registers.838[10] [21]),
    .B(_5220__bF$buf5),
    .Y(_5250_)
);

AOI21X1 _15430_ (
    .A(_4841__bF$buf4),
    .B(_5220__bF$buf4),
    .C(_5250_),
    .Y(_3807_)
);

NOR2X1 _15431_ (
    .A(\datapath.registers.838[10] [22]),
    .B(_5220__bF$buf3),
    .Y(_5251_)
);

AOI21X1 _15432_ (
    .A(_4843__bF$buf4),
    .B(_5220__bF$buf2),
    .C(_5251_),
    .Y(_3808_)
);

NOR2X1 _15433_ (
    .A(\datapath.registers.838[10] [23]),
    .B(_5220__bF$buf1),
    .Y(_5252_)
);

AOI21X1 _15434_ (
    .A(_4845__bF$buf4),
    .B(_5220__bF$buf0),
    .C(_5252_),
    .Y(_3809_)
);

INVX1 _15435_ (
    .A(\datapath.registers.838[10] [24]),
    .Y(_5253_)
);

NAND2X1 _15436_ (
    .A(\datapath.rd [24]),
    .B(_5220__bF$buf7),
    .Y(_5254_)
);

OAI21X1 _15437_ (
    .A(_5253_),
    .B(_5220__bF$buf6),
    .C(_5254_),
    .Y(_3810_)
);

NOR2X1 _15438_ (
    .A(\datapath.registers.838[10] [25]),
    .B(_5220__bF$buf5),
    .Y(_5255_)
);

AOI21X1 _15439_ (
    .A(_4849__bF$buf4),
    .B(_5220__bF$buf4),
    .C(_5255_),
    .Y(_3811_)
);

NOR2X1 _15440_ (
    .A(\datapath.registers.838[10] [26]),
    .B(_5220__bF$buf3),
    .Y(_5256_)
);

AOI21X1 _15441_ (
    .A(_4851__bF$buf3),
    .B(_5220__bF$buf2),
    .C(_5256_),
    .Y(_3812_)
);

NOR2X1 _15442_ (
    .A(\datapath.registers.838[10] [27]),
    .B(_5220__bF$buf1),
    .Y(_5257_)
);

AOI21X1 _15443_ (
    .A(_4853__bF$buf4),
    .B(_5220__bF$buf0),
    .C(_5257_),
    .Y(_3813_)
);

NOR2X1 _15444_ (
    .A(\datapath.registers.838[10] [28]),
    .B(_5220__bF$buf7),
    .Y(_5258_)
);

AOI21X1 _15445_ (
    .A(_4855__bF$buf3),
    .B(_5220__bF$buf6),
    .C(_5258_),
    .Y(_3814_)
);

NOR2X1 _15446_ (
    .A(\datapath.registers.838[10] [29]),
    .B(_5220__bF$buf5),
    .Y(_5259_)
);

AOI21X1 _15447_ (
    .A(_4857__bF$buf3),
    .B(_5220__bF$buf4),
    .C(_5259_),
    .Y(_3815_)
);

INVX1 _15448_ (
    .A(\datapath.registers.838[10] [30]),
    .Y(_5260_)
);

NAND2X1 _15449_ (
    .A(\datapath.rd [30]),
    .B(_5220__bF$buf3),
    .Y(_5261_)
);

OAI21X1 _15450_ (
    .A(_5260_),
    .B(_5220__bF$buf2),
    .C(_5261_),
    .Y(_3817_)
);

NOR2X1 _15451_ (
    .A(\datapath.registers.838[10] [31]),
    .B(_5220__bF$buf1),
    .Y(_5262_)
);

AOI21X1 _15452_ (
    .A(_4861__bF$buf3),
    .B(_5220__bF$buf0),
    .C(_5262_),
    .Y(_3818_)
);

INVX1 _15453_ (
    .A(\datapath.registers.838[9] [0]),
    .Y(_5263_)
);

NOR2X1 _15454_ (
    .A(_4968__bF$buf7),
    .B(_5185__bF$buf1),
    .Y(_5264_)
);

NAND2X1 _15455_ (
    .A(\datapath.rd [0]),
    .B(_5264__bF$buf7),
    .Y(_5265_)
);

OAI21X1 _15456_ (
    .A(_5263_),
    .B(_5264__bF$buf6),
    .C(_5265_),
    .Y(_4754_)
);

NOR2X1 _15457_ (
    .A(\datapath.registers.838[9] [1]),
    .B(_5264__bF$buf5),
    .Y(_5266_)
);

AOI21X1 _15458_ (
    .A(_4801__bF$buf2),
    .B(_5264__bF$buf4),
    .C(_5266_),
    .Y(_4765_)
);

INVX1 _15459_ (
    .A(\datapath.registers.838[9] [2]),
    .Y(_5267_)
);

NAND2X1 _15460_ (
    .A(\datapath.rd [2]),
    .B(_5264__bF$buf3),
    .Y(_5268_)
);

OAI21X1 _15461_ (
    .A(_5267_),
    .B(_5264__bF$buf2),
    .C(_5268_),
    .Y(_4776_)
);

INVX1 _15462_ (
    .A(\datapath.registers.838[9] [3]),
    .Y(_5269_)
);

NAND2X1 _15463_ (
    .A(\datapath.rd [3]),
    .B(_5264__bF$buf1),
    .Y(_5270_)
);

OAI21X1 _15464_ (
    .A(_5269_),
    .B(_5264__bF$buf0),
    .C(_5270_),
    .Y(_4779_)
);

NOR2X1 _15465_ (
    .A(\datapath.registers.838[9] [4]),
    .B(_5264__bF$buf7),
    .Y(_5271_)
);

AOI21X1 _15466_ (
    .A(_4807__bF$buf3),
    .B(_5264__bF$buf6),
    .C(_5271_),
    .Y(_4780_)
);

NOR2X1 _15467_ (
    .A(\datapath.registers.838[9] [5]),
    .B(_5264__bF$buf5),
    .Y(_5272_)
);

AOI21X1 _15468_ (
    .A(_4809__bF$buf3),
    .B(_5264__bF$buf4),
    .C(_5272_),
    .Y(_4781_)
);

INVX1 _15469_ (
    .A(\datapath.registers.838[9] [6]),
    .Y(_5273_)
);

NAND2X1 _15470_ (
    .A(\datapath.rd [6]),
    .B(_5264__bF$buf3),
    .Y(_5274_)
);

OAI21X1 _15471_ (
    .A(_5273_),
    .B(_5264__bF$buf2),
    .C(_5274_),
    .Y(_4782_)
);

NOR2X1 _15472_ (
    .A(\datapath.registers.838[9] [7]),
    .B(_5264__bF$buf1),
    .Y(_5275_)
);

AOI21X1 _15473_ (
    .A(_4813__bF$buf2),
    .B(_5264__bF$buf0),
    .C(_5275_),
    .Y(_4783_)
);

NOR2X1 _15474_ (
    .A(\datapath.registers.838[9] [8]),
    .B(_5264__bF$buf7),
    .Y(_5276_)
);

AOI21X1 _15475_ (
    .A(_4815__bF$buf2),
    .B(_5264__bF$buf6),
    .C(_5276_),
    .Y(_4784_)
);

INVX1 _15476_ (
    .A(\datapath.registers.838[9] [9]),
    .Y(_5277_)
);

NAND2X1 _15477_ (
    .A(\datapath.rd [9]),
    .B(_5264__bF$buf5),
    .Y(_5278_)
);

OAI21X1 _15478_ (
    .A(_5277_),
    .B(_5264__bF$buf4),
    .C(_5278_),
    .Y(_4785_)
);

NOR2X1 _15479_ (
    .A(\datapath.registers.838[9] [10]),
    .B(_5264__bF$buf3),
    .Y(_5279_)
);

AOI21X1 _15480_ (
    .A(_4819__bF$buf3),
    .B(_5264__bF$buf2),
    .C(_5279_),
    .Y(_4755_)
);

NOR2X1 _15481_ (
    .A(\datapath.registers.838[9] [11]),
    .B(_5264__bF$buf1),
    .Y(_5280_)
);

AOI21X1 _15482_ (
    .A(_4821__bF$buf2),
    .B(_5264__bF$buf0),
    .C(_5280_),
    .Y(_4756_)
);

INVX1 _15483_ (
    .A(\datapath.registers.838[9] [12]),
    .Y(_5281_)
);

NAND2X1 _15484_ (
    .A(\datapath.rd [12]),
    .B(_5264__bF$buf7),
    .Y(_5282_)
);

OAI21X1 _15485_ (
    .A(_5281_),
    .B(_5264__bF$buf6),
    .C(_5282_),
    .Y(_4757_)
);

NOR2X1 _15486_ (
    .A(\datapath.registers.838[9] [13]),
    .B(_5264__bF$buf5),
    .Y(_5283_)
);

AOI21X1 _15487_ (
    .A(_4825__bF$buf2),
    .B(_5264__bF$buf4),
    .C(_5283_),
    .Y(_4758_)
);

NOR2X1 _15488_ (
    .A(\datapath.registers.838[9] [14]),
    .B(_5264__bF$buf3),
    .Y(_5284_)
);

AOI21X1 _15489_ (
    .A(_4827__bF$buf2),
    .B(_5264__bF$buf2),
    .C(_5284_),
    .Y(_4759_)
);

NOR2X1 _15490_ (
    .A(\datapath.registers.838[9] [15]),
    .B(_5264__bF$buf1),
    .Y(_5285_)
);

AOI21X1 _15491_ (
    .A(_4829__bF$buf2),
    .B(_5264__bF$buf0),
    .C(_5285_),
    .Y(_4760_)
);

NOR2X1 _15492_ (
    .A(\datapath.registers.838[9] [16]),
    .B(_5264__bF$buf7),
    .Y(_5286_)
);

AOI21X1 _15493_ (
    .A(_4831__bF$buf2),
    .B(_5264__bF$buf6),
    .C(_5286_),
    .Y(_4761_)
);

INVX1 _15494_ (
    .A(\datapath.registers.838[9] [17]),
    .Y(_5287_)
);

NAND2X1 _15495_ (
    .A(\datapath.rd [17]),
    .B(_5264__bF$buf5),
    .Y(_5288_)
);

OAI21X1 _15496_ (
    .A(_5287_),
    .B(_5264__bF$buf4),
    .C(_5288_),
    .Y(_4762_)
);

INVX1 _15497_ (
    .A(\datapath.registers.838[9] [18]),
    .Y(_5289_)
);

NAND2X1 _15498_ (
    .A(\datapath.rd [18]),
    .B(_5264__bF$buf3),
    .Y(_5290_)
);

OAI21X1 _15499_ (
    .A(_5289_),
    .B(_5264__bF$buf2),
    .C(_5290_),
    .Y(_4763_)
);

INVX1 _15500_ (
    .A(\datapath.registers.838[9] [19]),
    .Y(_5291_)
);

NAND2X1 _15501_ (
    .A(\datapath.rd [19]),
    .B(_5264__bF$buf1),
    .Y(_5292_)
);

OAI21X1 _15502_ (
    .A(_5291_),
    .B(_5264__bF$buf0),
    .C(_5292_),
    .Y(_4764_)
);

NOR2X1 _15503_ (
    .A(\datapath.registers.838[9] [20]),
    .B(_5264__bF$buf7),
    .Y(_5293_)
);

AOI21X1 _15504_ (
    .A(_4839__bF$buf2),
    .B(_5264__bF$buf6),
    .C(_5293_),
    .Y(_4766_)
);

NOR2X1 _15505_ (
    .A(\datapath.registers.838[9] [21]),
    .B(_5264__bF$buf5),
    .Y(_5294_)
);

AOI21X1 _15506_ (
    .A(_4841__bF$buf3),
    .B(_5264__bF$buf4),
    .C(_5294_),
    .Y(_4767_)
);

NOR2X1 _15507_ (
    .A(\datapath.registers.838[9] [22]),
    .B(_5264__bF$buf3),
    .Y(_5295_)
);

AOI21X1 _15508_ (
    .A(_4843__bF$buf3),
    .B(_5264__bF$buf2),
    .C(_5295_),
    .Y(_4768_)
);

NOR2X1 _15509_ (
    .A(\datapath.registers.838[9] [23]),
    .B(_5264__bF$buf1),
    .Y(_5296_)
);

AOI21X1 _15510_ (
    .A(_4845__bF$buf3),
    .B(_5264__bF$buf0),
    .C(_5296_),
    .Y(_4769_)
);

INVX1 _15511_ (
    .A(\datapath.registers.838[9] [24]),
    .Y(_5297_)
);

NAND2X1 _15512_ (
    .A(\datapath.rd [24]),
    .B(_5264__bF$buf7),
    .Y(_5298_)
);

OAI21X1 _15513_ (
    .A(_5297_),
    .B(_5264__bF$buf6),
    .C(_5298_),
    .Y(_4770_)
);

NOR2X1 _15514_ (
    .A(\datapath.registers.838[9] [25]),
    .B(_5264__bF$buf5),
    .Y(_5299_)
);

AOI21X1 _15515_ (
    .A(_4849__bF$buf3),
    .B(_5264__bF$buf4),
    .C(_5299_),
    .Y(_4771_)
);

NOR2X1 _15516_ (
    .A(\datapath.registers.838[9] [26]),
    .B(_5264__bF$buf3),
    .Y(_5300_)
);

AOI21X1 _15517_ (
    .A(_4851__bF$buf2),
    .B(_5264__bF$buf2),
    .C(_5300_),
    .Y(_4772_)
);

NOR2X1 _15518_ (
    .A(\datapath.registers.838[9] [27]),
    .B(_5264__bF$buf1),
    .Y(_5301_)
);

AOI21X1 _15519_ (
    .A(_4853__bF$buf3),
    .B(_5264__bF$buf0),
    .C(_5301_),
    .Y(_4773_)
);

NOR2X1 _15520_ (
    .A(\datapath.registers.838[9] [28]),
    .B(_5264__bF$buf7),
    .Y(_5302_)
);

AOI21X1 _15521_ (
    .A(_4855__bF$buf2),
    .B(_5264__bF$buf6),
    .C(_5302_),
    .Y(_4774_)
);

NOR2X1 _15522_ (
    .A(\datapath.registers.838[9] [29]),
    .B(_5264__bF$buf5),
    .Y(_5303_)
);

AOI21X1 _15523_ (
    .A(_4857__bF$buf2),
    .B(_5264__bF$buf4),
    .C(_5303_),
    .Y(_4775_)
);

INVX1 _15524_ (
    .A(\datapath.registers.838[9] [30]),
    .Y(_5304_)
);

NAND2X1 _15525_ (
    .A(\datapath.rd [30]),
    .B(_5264__bF$buf3),
    .Y(_5305_)
);

OAI21X1 _15526_ (
    .A(_5304_),
    .B(_5264__bF$buf2),
    .C(_5305_),
    .Y(_4777_)
);

NOR2X1 _15527_ (
    .A(\datapath.registers.838[9] [31]),
    .B(_5264__bF$buf1),
    .Y(_5306_)
);

AOI21X1 _15528_ (
    .A(_4861__bF$buf2),
    .B(_5264__bF$buf0),
    .C(_5306_),
    .Y(_4778_)
);

NOR2X1 _15529_ (
    .A(_4790_),
    .B(_5185__bF$buf0),
    .Y(_5307_)
);

NAND2X1 _15530_ (
    .A(_5015_),
    .B(_5307_),
    .Y(_5308_)
);

NAND2X1 _15531_ (
    .A(\datapath.registers.838[8] [0]),
    .B(_5308__bF$buf7),
    .Y(_5309_)
);

OAI21X1 _15532_ (
    .A(_4786__bF$buf3),
    .B(_5308__bF$buf6),
    .C(_5309_),
    .Y(_4722_)
);

NAND2X1 _15533_ (
    .A(\datapath.registers.838[8] [1]),
    .B(_5308__bF$buf5),
    .Y(_5310_)
);

OAI21X1 _15534_ (
    .A(_4801__bF$buf1),
    .B(_5308__bF$buf4),
    .C(_5310_),
    .Y(_4733_)
);

NAND2X1 _15535_ (
    .A(\datapath.registers.838[8] [2]),
    .B(_5308__bF$buf3),
    .Y(_5311_)
);

OAI21X1 _15536_ (
    .A(_4803__bF$buf3),
    .B(_5308__bF$buf2),
    .C(_5311_),
    .Y(_4744_)
);

NAND2X1 _15537_ (
    .A(\datapath.registers.838[8] [3]),
    .B(_5308__bF$buf1),
    .Y(_5312_)
);

OAI21X1 _15538_ (
    .A(_4805__bF$buf4),
    .B(_5308__bF$buf0),
    .C(_5312_),
    .Y(_4747_)
);

NAND2X1 _15539_ (
    .A(\datapath.registers.838[8] [4]),
    .B(_5308__bF$buf7),
    .Y(_5313_)
);

OAI21X1 _15540_ (
    .A(_4807__bF$buf2),
    .B(_5308__bF$buf6),
    .C(_5313_),
    .Y(_4748_)
);

NAND2X1 _15541_ (
    .A(\datapath.registers.838[8] [5]),
    .B(_5308__bF$buf5),
    .Y(_5314_)
);

OAI21X1 _15542_ (
    .A(_4809__bF$buf2),
    .B(_5308__bF$buf4),
    .C(_5314_),
    .Y(_4749_)
);

NAND2X1 _15543_ (
    .A(\datapath.registers.838[8] [6]),
    .B(_5308__bF$buf3),
    .Y(_5315_)
);

OAI21X1 _15544_ (
    .A(_4811__bF$buf4),
    .B(_5308__bF$buf2),
    .C(_5315_),
    .Y(_4750_)
);

NAND2X1 _15545_ (
    .A(\datapath.registers.838[8] [7]),
    .B(_5308__bF$buf1),
    .Y(_5316_)
);

OAI21X1 _15546_ (
    .A(_4813__bF$buf1),
    .B(_5308__bF$buf0),
    .C(_5316_),
    .Y(_4751_)
);

NAND2X1 _15547_ (
    .A(\datapath.registers.838[8] [8]),
    .B(_5308__bF$buf7),
    .Y(_5317_)
);

OAI21X1 _15548_ (
    .A(_4815__bF$buf1),
    .B(_5308__bF$buf6),
    .C(_5317_),
    .Y(_4752_)
);

NAND2X1 _15549_ (
    .A(\datapath.registers.838[8] [9]),
    .B(_5308__bF$buf5),
    .Y(_5318_)
);

OAI21X1 _15550_ (
    .A(_4817__bF$buf4),
    .B(_5308__bF$buf4),
    .C(_5318_),
    .Y(_4753_)
);

NAND2X1 _15551_ (
    .A(\datapath.registers.838[8] [10]),
    .B(_5308__bF$buf3),
    .Y(_5319_)
);

OAI21X1 _15552_ (
    .A(_4819__bF$buf2),
    .B(_5308__bF$buf2),
    .C(_5319_),
    .Y(_4723_)
);

NAND2X1 _15553_ (
    .A(\datapath.registers.838[8] [11]),
    .B(_5308__bF$buf1),
    .Y(_5320_)
);

OAI21X1 _15554_ (
    .A(_4821__bF$buf1),
    .B(_5308__bF$buf0),
    .C(_5320_),
    .Y(_4724_)
);

NAND2X1 _15555_ (
    .A(\datapath.registers.838[8] [12]),
    .B(_5308__bF$buf7),
    .Y(_5321_)
);

OAI21X1 _15556_ (
    .A(_4823__bF$buf3),
    .B(_5308__bF$buf6),
    .C(_5321_),
    .Y(_4725_)
);

NAND2X1 _15557_ (
    .A(\datapath.registers.838[8] [13]),
    .B(_5308__bF$buf5),
    .Y(_5322_)
);

OAI21X1 _15558_ (
    .A(_4825__bF$buf1),
    .B(_5308__bF$buf4),
    .C(_5322_),
    .Y(_4726_)
);

NAND2X1 _15559_ (
    .A(\datapath.registers.838[8] [14]),
    .B(_5308__bF$buf3),
    .Y(_5323_)
);

OAI21X1 _15560_ (
    .A(_4827__bF$buf1),
    .B(_5308__bF$buf2),
    .C(_5323_),
    .Y(_4727_)
);

NAND2X1 _15561_ (
    .A(\datapath.registers.838[8] [15]),
    .B(_5308__bF$buf1),
    .Y(_5324_)
);

OAI21X1 _15562_ (
    .A(_4829__bF$buf1),
    .B(_5308__bF$buf0),
    .C(_5324_),
    .Y(_4728_)
);

NAND2X1 _15563_ (
    .A(\datapath.registers.838[8] [16]),
    .B(_5308__bF$buf7),
    .Y(_5325_)
);

OAI21X1 _15564_ (
    .A(_4831__bF$buf1),
    .B(_5308__bF$buf6),
    .C(_5325_),
    .Y(_4729_)
);

NAND2X1 _15565_ (
    .A(\datapath.registers.838[8] [17]),
    .B(_5308__bF$buf5),
    .Y(_5326_)
);

OAI21X1 _15566_ (
    .A(_4833__bF$buf3),
    .B(_5308__bF$buf4),
    .C(_5326_),
    .Y(_4730_)
);

NAND2X1 _15567_ (
    .A(\datapath.registers.838[8] [18]),
    .B(_5308__bF$buf3),
    .Y(_5327_)
);

OAI21X1 _15568_ (
    .A(_4835__bF$buf3),
    .B(_5308__bF$buf2),
    .C(_5327_),
    .Y(_4731_)
);

NAND2X1 _15569_ (
    .A(\datapath.registers.838[8] [19]),
    .B(_5308__bF$buf1),
    .Y(_5328_)
);

OAI21X1 _15570_ (
    .A(_4837__bF$buf4),
    .B(_5308__bF$buf0),
    .C(_5328_),
    .Y(_4732_)
);

NAND2X1 _15571_ (
    .A(\datapath.registers.838[8] [20]),
    .B(_5308__bF$buf7),
    .Y(_5329_)
);

OAI21X1 _15572_ (
    .A(_4839__bF$buf1),
    .B(_5308__bF$buf6),
    .C(_5329_),
    .Y(_4734_)
);

NAND2X1 _15573_ (
    .A(\datapath.registers.838[8] [21]),
    .B(_5308__bF$buf5),
    .Y(_5330_)
);

OAI21X1 _15574_ (
    .A(_4841__bF$buf2),
    .B(_5308__bF$buf4),
    .C(_5330_),
    .Y(_4735_)
);

NAND2X1 _15575_ (
    .A(\datapath.registers.838[8] [22]),
    .B(_5308__bF$buf3),
    .Y(_5331_)
);

OAI21X1 _15576_ (
    .A(_4843__bF$buf2),
    .B(_5308__bF$buf2),
    .C(_5331_),
    .Y(_4736_)
);

NAND2X1 _15577_ (
    .A(\datapath.registers.838[8] [23]),
    .B(_5308__bF$buf1),
    .Y(_5332_)
);

OAI21X1 _15578_ (
    .A(_4845__bF$buf2),
    .B(_5308__bF$buf0),
    .C(_5332_),
    .Y(_4737_)
);

NAND2X1 _15579_ (
    .A(\datapath.registers.838[8] [24]),
    .B(_5308__bF$buf7),
    .Y(_5333_)
);

OAI21X1 _15580_ (
    .A(_4847__bF$buf4),
    .B(_5308__bF$buf6),
    .C(_5333_),
    .Y(_4738_)
);

NAND2X1 _15581_ (
    .A(\datapath.registers.838[8] [25]),
    .B(_5308__bF$buf5),
    .Y(_5334_)
);

OAI21X1 _15582_ (
    .A(_4849__bF$buf2),
    .B(_5308__bF$buf4),
    .C(_5334_),
    .Y(_4739_)
);

NAND2X1 _15583_ (
    .A(\datapath.registers.838[8] [26]),
    .B(_5308__bF$buf3),
    .Y(_5335_)
);

OAI21X1 _15584_ (
    .A(_4851__bF$buf1),
    .B(_5308__bF$buf2),
    .C(_5335_),
    .Y(_4740_)
);

NAND2X1 _15585_ (
    .A(\datapath.registers.838[8] [27]),
    .B(_5308__bF$buf1),
    .Y(_5336_)
);

OAI21X1 _15586_ (
    .A(_4853__bF$buf2),
    .B(_5308__bF$buf0),
    .C(_5336_),
    .Y(_4741_)
);

NAND2X1 _15587_ (
    .A(\datapath.registers.838[8] [28]),
    .B(_5308__bF$buf7),
    .Y(_5337_)
);

OAI21X1 _15588_ (
    .A(_4855__bF$buf1),
    .B(_5308__bF$buf6),
    .C(_5337_),
    .Y(_4742_)
);

NAND2X1 _15589_ (
    .A(\datapath.registers.838[8] [29]),
    .B(_5308__bF$buf5),
    .Y(_5338_)
);

OAI21X1 _15590_ (
    .A(_4857__bF$buf1),
    .B(_5308__bF$buf4),
    .C(_5338_),
    .Y(_4743_)
);

NAND2X1 _15591_ (
    .A(\datapath.registers.838[8] [30]),
    .B(_5308__bF$buf3),
    .Y(_5339_)
);

OAI21X1 _15592_ (
    .A(_4859__bF$buf3),
    .B(_5308__bF$buf2),
    .C(_5339_),
    .Y(_4745_)
);

NAND2X1 _15593_ (
    .A(\datapath.registers.838[8] [31]),
    .B(_5308__bF$buf1),
    .Y(_5340_)
);

OAI21X1 _15594_ (
    .A(_4861__bF$buf1),
    .B(_5308__bF$buf0),
    .C(_5340_),
    .Y(_4746_)
);

NAND3X1 _15595_ (
    .A(\datapath.wbinstr [9]),
    .B(_4792_),
    .C(_4793_),
    .Y(_5341_)
);

OR2X2 _15596_ (
    .A(_4899__bF$buf12),
    .B(_5341__bF$buf5),
    .Y(_5342_)
);

OAI21X1 _15597_ (
    .A(_5341__bF$buf4),
    .B(_4899__bF$buf11),
    .C(\datapath.registers.838[7] [0]),
    .Y(_5343_)
);

OAI21X1 _15598_ (
    .A(_4786__bF$buf2),
    .B(_5342__bF$buf4),
    .C(_5343_),
    .Y(_4690_)
);

OAI21X1 _15599_ (
    .A(_5341__bF$buf3),
    .B(_4899__bF$buf10),
    .C(\datapath.registers.838[7] [1]),
    .Y(_5344_)
);

OAI21X1 _15600_ (
    .A(_4801__bF$buf0),
    .B(_5342__bF$buf3),
    .C(_5344_),
    .Y(_4701_)
);

OAI21X1 _15601_ (
    .A(_5341__bF$buf2),
    .B(_4899__bF$buf9),
    .C(\datapath.registers.838[7] [2]),
    .Y(_5345_)
);

OAI21X1 _15602_ (
    .A(_4803__bF$buf2),
    .B(_5342__bF$buf2),
    .C(_5345_),
    .Y(_4712_)
);

OAI21X1 _15603_ (
    .A(_5341__bF$buf1),
    .B(_4899__bF$buf8),
    .C(\datapath.registers.838[7] [3]),
    .Y(_5346_)
);

OAI21X1 _15604_ (
    .A(_4805__bF$buf3),
    .B(_5342__bF$buf1),
    .C(_5346_),
    .Y(_4715_)
);

OAI21X1 _15605_ (
    .A(_5341__bF$buf0),
    .B(_4899__bF$buf7),
    .C(\datapath.registers.838[7] [4]),
    .Y(_5347_)
);

OAI21X1 _15606_ (
    .A(_4807__bF$buf1),
    .B(_5342__bF$buf0),
    .C(_5347_),
    .Y(_4716_)
);

OAI21X1 _15607_ (
    .A(_5341__bF$buf5),
    .B(_4899__bF$buf6),
    .C(\datapath.registers.838[7] [5]),
    .Y(_5348_)
);

OAI21X1 _15608_ (
    .A(_4809__bF$buf1),
    .B(_5342__bF$buf4),
    .C(_5348_),
    .Y(_4717_)
);

OAI21X1 _15609_ (
    .A(_5341__bF$buf4),
    .B(_4899__bF$buf5),
    .C(\datapath.registers.838[7] [6]),
    .Y(_5349_)
);

OAI21X1 _15610_ (
    .A(_4811__bF$buf3),
    .B(_5342__bF$buf3),
    .C(_5349_),
    .Y(_4718_)
);

OAI21X1 _15611_ (
    .A(_5341__bF$buf3),
    .B(_4899__bF$buf4),
    .C(\datapath.registers.838[7] [7]),
    .Y(_5350_)
);

OAI21X1 _15612_ (
    .A(_4813__bF$buf0),
    .B(_5342__bF$buf2),
    .C(_5350_),
    .Y(_4719_)
);

OAI21X1 _15613_ (
    .A(_5341__bF$buf2),
    .B(_4899__bF$buf3),
    .C(\datapath.registers.838[7] [8]),
    .Y(_5351_)
);

OAI21X1 _15614_ (
    .A(_4815__bF$buf0),
    .B(_5342__bF$buf1),
    .C(_5351_),
    .Y(_4720_)
);

OAI21X1 _15615_ (
    .A(_5341__bF$buf1),
    .B(_4899__bF$buf2),
    .C(\datapath.registers.838[7] [9]),
    .Y(_5352_)
);

OAI21X1 _15616_ (
    .A(_4817__bF$buf3),
    .B(_5342__bF$buf0),
    .C(_5352_),
    .Y(_4721_)
);

OAI21X1 _15617_ (
    .A(_5341__bF$buf0),
    .B(_4899__bF$buf1),
    .C(\datapath.registers.838[7] [10]),
    .Y(_5353_)
);

OAI21X1 _15618_ (
    .A(_4819__bF$buf1),
    .B(_5342__bF$buf4),
    .C(_5353_),
    .Y(_4691_)
);

OAI21X1 _15619_ (
    .A(_5341__bF$buf5),
    .B(_4899__bF$buf0),
    .C(\datapath.registers.838[7] [11]),
    .Y(_5354_)
);

OAI21X1 _15620_ (
    .A(_4821__bF$buf0),
    .B(_5342__bF$buf3),
    .C(_5354_),
    .Y(_4692_)
);

OAI21X1 _15621_ (
    .A(_5341__bF$buf4),
    .B(_4899__bF$buf13),
    .C(\datapath.registers.838[7] [12]),
    .Y(_5355_)
);

OAI21X1 _15622_ (
    .A(_4823__bF$buf2),
    .B(_5342__bF$buf2),
    .C(_5355_),
    .Y(_4693_)
);

OAI21X1 _15623_ (
    .A(_5341__bF$buf3),
    .B(_4899__bF$buf12),
    .C(\datapath.registers.838[7] [13]),
    .Y(_5356_)
);

OAI21X1 _15624_ (
    .A(_4825__bF$buf0),
    .B(_5342__bF$buf1),
    .C(_5356_),
    .Y(_4694_)
);

OAI21X1 _15625_ (
    .A(_5341__bF$buf2),
    .B(_4899__bF$buf11),
    .C(\datapath.registers.838[7] [14]),
    .Y(_5357_)
);

OAI21X1 _15626_ (
    .A(_4827__bF$buf0),
    .B(_5342__bF$buf0),
    .C(_5357_),
    .Y(_4695_)
);

OAI21X1 _15627_ (
    .A(_5341__bF$buf1),
    .B(_4899__bF$buf10),
    .C(\datapath.registers.838[7] [15]),
    .Y(_5358_)
);

OAI21X1 _15628_ (
    .A(_4829__bF$buf0),
    .B(_5342__bF$buf4),
    .C(_5358_),
    .Y(_4696_)
);

OAI21X1 _15629_ (
    .A(_5341__bF$buf0),
    .B(_4899__bF$buf9),
    .C(\datapath.registers.838[7] [16]),
    .Y(_5359_)
);

OAI21X1 _15630_ (
    .A(_4831__bF$buf0),
    .B(_5342__bF$buf3),
    .C(_5359_),
    .Y(_4697_)
);

OAI21X1 _15631_ (
    .A(_5341__bF$buf5),
    .B(_4899__bF$buf8),
    .C(\datapath.registers.838[7] [17]),
    .Y(_5360_)
);

OAI21X1 _15632_ (
    .A(_4833__bF$buf2),
    .B(_5342__bF$buf2),
    .C(_5360_),
    .Y(_4698_)
);

OAI21X1 _15633_ (
    .A(_5341__bF$buf4),
    .B(_4899__bF$buf7),
    .C(\datapath.registers.838[7] [18]),
    .Y(_5361_)
);

OAI21X1 _15634_ (
    .A(_4835__bF$buf2),
    .B(_5342__bF$buf1),
    .C(_5361_),
    .Y(_4699_)
);

OAI21X1 _15635_ (
    .A(_5341__bF$buf3),
    .B(_4899__bF$buf6),
    .C(\datapath.registers.838[7] [19]),
    .Y(_5362_)
);

OAI21X1 _15636_ (
    .A(_4837__bF$buf3),
    .B(_5342__bF$buf0),
    .C(_5362_),
    .Y(_4700_)
);

OAI21X1 _15637_ (
    .A(_5341__bF$buf2),
    .B(_4899__bF$buf5),
    .C(\datapath.registers.838[7] [20]),
    .Y(_5363_)
);

OAI21X1 _15638_ (
    .A(_4839__bF$buf0),
    .B(_5342__bF$buf4),
    .C(_5363_),
    .Y(_4702_)
);

OAI21X1 _15639_ (
    .A(_5341__bF$buf1),
    .B(_4899__bF$buf4),
    .C(\datapath.registers.838[7] [21]),
    .Y(_5364_)
);

OAI21X1 _15640_ (
    .A(_4841__bF$buf1),
    .B(_5342__bF$buf3),
    .C(_5364_),
    .Y(_4703_)
);

OAI21X1 _15641_ (
    .A(_5341__bF$buf0),
    .B(_4899__bF$buf3),
    .C(\datapath.registers.838[7] [22]),
    .Y(_5365_)
);

OAI21X1 _15642_ (
    .A(_4843__bF$buf1),
    .B(_5342__bF$buf2),
    .C(_5365_),
    .Y(_4704_)
);

OAI21X1 _15643_ (
    .A(_5341__bF$buf5),
    .B(_4899__bF$buf2),
    .C(\datapath.registers.838[7] [23]),
    .Y(_5366_)
);

OAI21X1 _15644_ (
    .A(_4845__bF$buf1),
    .B(_5342__bF$buf1),
    .C(_5366_),
    .Y(_4705_)
);

OAI21X1 _15645_ (
    .A(_5341__bF$buf4),
    .B(_4899__bF$buf1),
    .C(\datapath.registers.838[7] [24]),
    .Y(_5367_)
);

OAI21X1 _15646_ (
    .A(_4847__bF$buf3),
    .B(_5342__bF$buf0),
    .C(_5367_),
    .Y(_4706_)
);

OAI21X1 _15647_ (
    .A(_5341__bF$buf3),
    .B(_4899__bF$buf0),
    .C(\datapath.registers.838[7] [25]),
    .Y(_5368_)
);

OAI21X1 _15648_ (
    .A(_4849__bF$buf1),
    .B(_5342__bF$buf4),
    .C(_5368_),
    .Y(_4707_)
);

OAI21X1 _15649_ (
    .A(_5341__bF$buf2),
    .B(_4899__bF$buf13),
    .C(\datapath.registers.838[7] [26]),
    .Y(_5369_)
);

OAI21X1 _15650_ (
    .A(_4851__bF$buf0),
    .B(_5342__bF$buf3),
    .C(_5369_),
    .Y(_4708_)
);

OAI21X1 _15651_ (
    .A(_5341__bF$buf1),
    .B(_4899__bF$buf12),
    .C(\datapath.registers.838[7] [27]),
    .Y(_5370_)
);

OAI21X1 _15652_ (
    .A(_4853__bF$buf1),
    .B(_5342__bF$buf2),
    .C(_5370_),
    .Y(_4709_)
);

OAI21X1 _15653_ (
    .A(_5341__bF$buf0),
    .B(_4899__bF$buf11),
    .C(\datapath.registers.838[7] [28]),
    .Y(_5371_)
);

OAI21X1 _15654_ (
    .A(_4855__bF$buf0),
    .B(_5342__bF$buf1),
    .C(_5371_),
    .Y(_4710_)
);

OAI21X1 _15655_ (
    .A(_5341__bF$buf5),
    .B(_4899__bF$buf10),
    .C(\datapath.registers.838[7] [29]),
    .Y(_5372_)
);

OAI21X1 _15656_ (
    .A(_4857__bF$buf0),
    .B(_5342__bF$buf0),
    .C(_5372_),
    .Y(_4711_)
);

OAI21X1 _15657_ (
    .A(_5341__bF$buf4),
    .B(_4899__bF$buf9),
    .C(\datapath.registers.838[7] [30]),
    .Y(_5373_)
);

OAI21X1 _15658_ (
    .A(_4859__bF$buf2),
    .B(_5342__bF$buf4),
    .C(_5373_),
    .Y(_4713_)
);

OAI21X1 _15659_ (
    .A(_5341__bF$buf3),
    .B(_4899__bF$buf8),
    .C(\datapath.registers.838[7] [31]),
    .Y(_5374_)
);

OAI21X1 _15660_ (
    .A(_4861__bF$buf0),
    .B(_5342__bF$buf3),
    .C(_5374_),
    .Y(_4714_)
);

NOR2X1 _15661_ (
    .A(_5341__bF$buf2),
    .B(_4934__bF$buf6),
    .Y(_5375_)
);

NOR2X1 _15662_ (
    .A(\datapath.registers.838[6] [0]),
    .B(_5375__bF$buf7),
    .Y(_5376_)
);

AOI21X1 _15663_ (
    .A(_4786__bF$buf1),
    .B(_5375__bF$buf6),
    .C(_5376_),
    .Y(_4658_)
);

NOR2X1 _15664_ (
    .A(\datapath.registers.838[6] [1]),
    .B(_5375__bF$buf5),
    .Y(_5377_)
);

AOI21X1 _15665_ (
    .A(_4801__bF$buf4),
    .B(_5375__bF$buf4),
    .C(_5377_),
    .Y(_4669_)
);

NOR2X1 _15666_ (
    .A(\datapath.registers.838[6] [2]),
    .B(_5375__bF$buf3),
    .Y(_5378_)
);

AOI21X1 _15667_ (
    .A(_4803__bF$buf1),
    .B(_5375__bF$buf2),
    .C(_5378_),
    .Y(_4680_)
);

NOR2X1 _15668_ (
    .A(\datapath.registers.838[6] [3]),
    .B(_5375__bF$buf1),
    .Y(_5379_)
);

AOI21X1 _15669_ (
    .A(_4805__bF$buf2),
    .B(_5375__bF$buf0),
    .C(_5379_),
    .Y(_4683_)
);

NOR2X1 _15670_ (
    .A(\datapath.registers.838[6] [4]),
    .B(_5375__bF$buf7),
    .Y(_5380_)
);

AOI21X1 _15671_ (
    .A(_4807__bF$buf0),
    .B(_5375__bF$buf6),
    .C(_5380_),
    .Y(_4684_)
);

NOR2X1 _15672_ (
    .A(\datapath.registers.838[6] [5]),
    .B(_5375__bF$buf5),
    .Y(_5381_)
);

AOI21X1 _15673_ (
    .A(_4809__bF$buf0),
    .B(_5375__bF$buf4),
    .C(_5381_),
    .Y(_4685_)
);

NOR2X1 _15674_ (
    .A(\datapath.registers.838[6] [6]),
    .B(_5375__bF$buf3),
    .Y(_5382_)
);

AOI21X1 _15675_ (
    .A(_4811__bF$buf2),
    .B(_5375__bF$buf2),
    .C(_5382_),
    .Y(_4686_)
);

NOR2X1 _15676_ (
    .A(\datapath.registers.838[6] [7]),
    .B(_5375__bF$buf1),
    .Y(_5383_)
);

AOI21X1 _15677_ (
    .A(_4813__bF$buf4),
    .B(_5375__bF$buf0),
    .C(_5383_),
    .Y(_4687_)
);

NOR2X1 _15678_ (
    .A(\datapath.registers.838[6] [8]),
    .B(_5375__bF$buf7),
    .Y(_5384_)
);

AOI21X1 _15679_ (
    .A(_4815__bF$buf4),
    .B(_5375__bF$buf6),
    .C(_5384_),
    .Y(_4688_)
);

NOR2X1 _15680_ (
    .A(\datapath.registers.838[6] [9]),
    .B(_5375__bF$buf5),
    .Y(_5385_)
);

AOI21X1 _15681_ (
    .A(_4817__bF$buf2),
    .B(_5375__bF$buf4),
    .C(_5385_),
    .Y(_4689_)
);

NOR2X1 _15682_ (
    .A(\datapath.registers.838[6] [10]),
    .B(_5375__bF$buf3),
    .Y(_5386_)
);

AOI21X1 _15683_ (
    .A(_4819__bF$buf0),
    .B(_5375__bF$buf2),
    .C(_5386_),
    .Y(_4659_)
);

NOR2X1 _15684_ (
    .A(\datapath.registers.838[6] [11]),
    .B(_5375__bF$buf1),
    .Y(_5387_)
);

AOI21X1 _15685_ (
    .A(_4821__bF$buf4),
    .B(_5375__bF$buf0),
    .C(_5387_),
    .Y(_4660_)
);

NOR2X1 _15686_ (
    .A(\datapath.registers.838[6] [12]),
    .B(_5375__bF$buf7),
    .Y(_5388_)
);

AOI21X1 _15687_ (
    .A(_4823__bF$buf1),
    .B(_5375__bF$buf6),
    .C(_5388_),
    .Y(_4661_)
);

NOR2X1 _15688_ (
    .A(\datapath.registers.838[6] [13]),
    .B(_5375__bF$buf5),
    .Y(_5389_)
);

AOI21X1 _15689_ (
    .A(_4825__bF$buf4),
    .B(_5375__bF$buf4),
    .C(_5389_),
    .Y(_4662_)
);

NOR2X1 _15690_ (
    .A(\datapath.registers.838[6] [14]),
    .B(_5375__bF$buf3),
    .Y(_5390_)
);

AOI21X1 _15691_ (
    .A(_4827__bF$buf4),
    .B(_5375__bF$buf2),
    .C(_5390_),
    .Y(_4663_)
);

NOR2X1 _15692_ (
    .A(\datapath.registers.838[6] [15]),
    .B(_5375__bF$buf1),
    .Y(_5391_)
);

AOI21X1 _15693_ (
    .A(_4829__bF$buf4),
    .B(_5375__bF$buf0),
    .C(_5391_),
    .Y(_4664_)
);

NOR2X1 _15694_ (
    .A(\datapath.registers.838[6] [16]),
    .B(_5375__bF$buf7),
    .Y(_5392_)
);

AOI21X1 _15695_ (
    .A(_4831__bF$buf4),
    .B(_5375__bF$buf6),
    .C(_5392_),
    .Y(_4665_)
);

NOR2X1 _15696_ (
    .A(\datapath.registers.838[6] [17]),
    .B(_5375__bF$buf5),
    .Y(_5393_)
);

AOI21X1 _15697_ (
    .A(_4833__bF$buf1),
    .B(_5375__bF$buf4),
    .C(_5393_),
    .Y(_4666_)
);

NOR2X1 _15698_ (
    .A(\datapath.registers.838[6] [18]),
    .B(_5375__bF$buf3),
    .Y(_5394_)
);

AOI21X1 _15699_ (
    .A(_4835__bF$buf1),
    .B(_5375__bF$buf2),
    .C(_5394_),
    .Y(_4667_)
);

NOR2X1 _15700_ (
    .A(\datapath.registers.838[6] [19]),
    .B(_5375__bF$buf1),
    .Y(_5395_)
);

AOI21X1 _15701_ (
    .A(_4837__bF$buf2),
    .B(_5375__bF$buf0),
    .C(_5395_),
    .Y(_4668_)
);

NOR2X1 _15702_ (
    .A(\datapath.registers.838[6] [20]),
    .B(_5375__bF$buf7),
    .Y(_5396_)
);

AOI21X1 _15703_ (
    .A(_4839__bF$buf4),
    .B(_5375__bF$buf6),
    .C(_5396_),
    .Y(_4670_)
);

NOR2X1 _15704_ (
    .A(\datapath.registers.838[6] [21]),
    .B(_5375__bF$buf5),
    .Y(_5397_)
);

AOI21X1 _15705_ (
    .A(_4841__bF$buf0),
    .B(_5375__bF$buf4),
    .C(_5397_),
    .Y(_4671_)
);

NOR2X1 _15706_ (
    .A(\datapath.registers.838[6] [22]),
    .B(_5375__bF$buf3),
    .Y(_5398_)
);

AOI21X1 _15707_ (
    .A(_4843__bF$buf0),
    .B(_5375__bF$buf2),
    .C(_5398_),
    .Y(_4672_)
);

NOR2X1 _15708_ (
    .A(\datapath.registers.838[6] [23]),
    .B(_5375__bF$buf1),
    .Y(_5399_)
);

AOI21X1 _15709_ (
    .A(_4845__bF$buf0),
    .B(_5375__bF$buf0),
    .C(_5399_),
    .Y(_4673_)
);

NOR2X1 _15710_ (
    .A(\datapath.registers.838[6] [24]),
    .B(_5375__bF$buf7),
    .Y(_5400_)
);

AOI21X1 _15711_ (
    .A(_4847__bF$buf2),
    .B(_5375__bF$buf6),
    .C(_5400_),
    .Y(_4674_)
);

NOR2X1 _15712_ (
    .A(\datapath.registers.838[6] [25]),
    .B(_5375__bF$buf5),
    .Y(_5401_)
);

AOI21X1 _15713_ (
    .A(_4849__bF$buf0),
    .B(_5375__bF$buf4),
    .C(_5401_),
    .Y(_4675_)
);

NOR2X1 _15714_ (
    .A(\datapath.registers.838[6] [26]),
    .B(_5375__bF$buf3),
    .Y(_5402_)
);

AOI21X1 _15715_ (
    .A(_4851__bF$buf4),
    .B(_5375__bF$buf2),
    .C(_5402_),
    .Y(_4676_)
);

NOR2X1 _15716_ (
    .A(\datapath.registers.838[6] [27]),
    .B(_5375__bF$buf1),
    .Y(_5403_)
);

AOI21X1 _15717_ (
    .A(_4853__bF$buf0),
    .B(_5375__bF$buf0),
    .C(_5403_),
    .Y(_4677_)
);

NOR2X1 _15718_ (
    .A(\datapath.registers.838[6] [28]),
    .B(_5375__bF$buf7),
    .Y(_5404_)
);

AOI21X1 _15719_ (
    .A(_4855__bF$buf4),
    .B(_5375__bF$buf6),
    .C(_5404_),
    .Y(_4678_)
);

NOR2X1 _15720_ (
    .A(\datapath.registers.838[6] [29]),
    .B(_5375__bF$buf5),
    .Y(_5405_)
);

AOI21X1 _15721_ (
    .A(_4857__bF$buf4),
    .B(_5375__bF$buf4),
    .C(_5405_),
    .Y(_4679_)
);

NOR2X1 _15722_ (
    .A(\datapath.registers.838[6] [30]),
    .B(_5375__bF$buf3),
    .Y(_5406_)
);

AOI21X1 _15723_ (
    .A(_4859__bF$buf1),
    .B(_5375__bF$buf2),
    .C(_5406_),
    .Y(_4681_)
);

NOR2X1 _15724_ (
    .A(\datapath.registers.838[6] [31]),
    .B(_5375__bF$buf1),
    .Y(_5407_)
);

AOI21X1 _15725_ (
    .A(_4861__bF$buf4),
    .B(_5375__bF$buf0),
    .C(_5407_),
    .Y(_4682_)
);

NOR2X1 _15726_ (
    .A(_5341__bF$buf1),
    .B(_4968__bF$buf6),
    .Y(_5408_)
);

NOR2X1 _15727_ (
    .A(\datapath.registers.838[5] [0]),
    .B(_5408__bF$buf7),
    .Y(_5409_)
);

AOI21X1 _15728_ (
    .A(_4786__bF$buf0),
    .B(_5408__bF$buf6),
    .C(_5409_),
    .Y(_4626_)
);

NOR2X1 _15729_ (
    .A(\datapath.registers.838[5] [1]),
    .B(_5408__bF$buf5),
    .Y(_5410_)
);

AOI21X1 _15730_ (
    .A(_4801__bF$buf3),
    .B(_5408__bF$buf4),
    .C(_5410_),
    .Y(_4637_)
);

NOR2X1 _15731_ (
    .A(\datapath.registers.838[5] [2]),
    .B(_5408__bF$buf3),
    .Y(_5411_)
);

AOI21X1 _15732_ (
    .A(_4803__bF$buf0),
    .B(_5408__bF$buf2),
    .C(_5411_),
    .Y(_4648_)
);

NOR2X1 _15733_ (
    .A(\datapath.registers.838[5] [3]),
    .B(_5408__bF$buf1),
    .Y(_5412_)
);

AOI21X1 _15734_ (
    .A(_4805__bF$buf1),
    .B(_5408__bF$buf0),
    .C(_5412_),
    .Y(_4651_)
);

NOR2X1 _15735_ (
    .A(\datapath.registers.838[5] [4]),
    .B(_5408__bF$buf7),
    .Y(_5413_)
);

AOI21X1 _15736_ (
    .A(_4807__bF$buf4),
    .B(_5408__bF$buf6),
    .C(_5413_),
    .Y(_4652_)
);

NOR2X1 _15737_ (
    .A(\datapath.registers.838[5] [5]),
    .B(_5408__bF$buf5),
    .Y(_5414_)
);

AOI21X1 _15738_ (
    .A(_4809__bF$buf4),
    .B(_5408__bF$buf4),
    .C(_5414_),
    .Y(_4653_)
);

NOR2X1 _15739_ (
    .A(\datapath.registers.838[5] [6]),
    .B(_5408__bF$buf3),
    .Y(_5415_)
);

AOI21X1 _15740_ (
    .A(_4811__bF$buf1),
    .B(_5408__bF$buf2),
    .C(_5415_),
    .Y(_4654_)
);

NOR2X1 _15741_ (
    .A(\datapath.registers.838[5] [7]),
    .B(_5408__bF$buf1),
    .Y(_5416_)
);

AOI21X1 _15742_ (
    .A(_4813__bF$buf3),
    .B(_5408__bF$buf0),
    .C(_5416_),
    .Y(_4655_)
);

NOR2X1 _15743_ (
    .A(\datapath.registers.838[5] [8]),
    .B(_5408__bF$buf7),
    .Y(_5417_)
);

AOI21X1 _15744_ (
    .A(_4815__bF$buf3),
    .B(_5408__bF$buf6),
    .C(_5417_),
    .Y(_4656_)
);

NOR2X1 _15745_ (
    .A(\datapath.registers.838[5] [9]),
    .B(_5408__bF$buf5),
    .Y(_5418_)
);

AOI21X1 _15746_ (
    .A(_4817__bF$buf1),
    .B(_5408__bF$buf4),
    .C(_5418_),
    .Y(_4657_)
);

NOR2X1 _15747_ (
    .A(\datapath.registers.838[5] [10]),
    .B(_5408__bF$buf3),
    .Y(_5419_)
);

AOI21X1 _15748_ (
    .A(_4819__bF$buf4),
    .B(_5408__bF$buf2),
    .C(_5419_),
    .Y(_4627_)
);

NOR2X1 _15749_ (
    .A(\datapath.registers.838[5] [11]),
    .B(_5408__bF$buf1),
    .Y(_5420_)
);

AOI21X1 _15750_ (
    .A(_4821__bF$buf3),
    .B(_5408__bF$buf0),
    .C(_5420_),
    .Y(_4628_)
);

NOR2X1 _15751_ (
    .A(\datapath.registers.838[5] [12]),
    .B(_5408__bF$buf7),
    .Y(_5421_)
);

AOI21X1 _15752_ (
    .A(_4823__bF$buf0),
    .B(_5408__bF$buf6),
    .C(_5421_),
    .Y(_4629_)
);

NOR2X1 _15753_ (
    .A(\datapath.registers.838[5] [13]),
    .B(_5408__bF$buf5),
    .Y(_5422_)
);

AOI21X1 _15754_ (
    .A(_4825__bF$buf3),
    .B(_5408__bF$buf4),
    .C(_5422_),
    .Y(_4630_)
);

NOR2X1 _15755_ (
    .A(\datapath.registers.838[5] [14]),
    .B(_5408__bF$buf3),
    .Y(_5423_)
);

AOI21X1 _15756_ (
    .A(_4827__bF$buf3),
    .B(_5408__bF$buf2),
    .C(_5423_),
    .Y(_4631_)
);

NOR2X1 _15757_ (
    .A(\datapath.registers.838[5] [15]),
    .B(_5408__bF$buf1),
    .Y(_5424_)
);

AOI21X1 _15758_ (
    .A(_4829__bF$buf3),
    .B(_5408__bF$buf0),
    .C(_5424_),
    .Y(_4632_)
);

NOR2X1 _15759_ (
    .A(\datapath.registers.838[5] [16]),
    .B(_5408__bF$buf7),
    .Y(_5425_)
);

AOI21X1 _15760_ (
    .A(_4831__bF$buf3),
    .B(_5408__bF$buf6),
    .C(_5425_),
    .Y(_4633_)
);

NOR2X1 _15761_ (
    .A(\datapath.registers.838[5] [17]),
    .B(_5408__bF$buf5),
    .Y(_5426_)
);

AOI21X1 _15762_ (
    .A(_4833__bF$buf0),
    .B(_5408__bF$buf4),
    .C(_5426_),
    .Y(_4634_)
);

NOR2X1 _15763_ (
    .A(\datapath.registers.838[5] [18]),
    .B(_5408__bF$buf3),
    .Y(_5427_)
);

AOI21X1 _15764_ (
    .A(_4835__bF$buf0),
    .B(_5408__bF$buf2),
    .C(_5427_),
    .Y(_4635_)
);

NOR2X1 _15765_ (
    .A(\datapath.registers.838[5] [19]),
    .B(_5408__bF$buf1),
    .Y(_5428_)
);

AOI21X1 _15766_ (
    .A(_4837__bF$buf1),
    .B(_5408__bF$buf0),
    .C(_5428_),
    .Y(_4636_)
);

NOR2X1 _15767_ (
    .A(\datapath.registers.838[5] [20]),
    .B(_5408__bF$buf7),
    .Y(_5429_)
);

AOI21X1 _15768_ (
    .A(_4839__bF$buf3),
    .B(_5408__bF$buf6),
    .C(_5429_),
    .Y(_4638_)
);

NOR2X1 _15769_ (
    .A(\datapath.registers.838[5] [21]),
    .B(_5408__bF$buf5),
    .Y(_5430_)
);

AOI21X1 _15770_ (
    .A(_4841__bF$buf4),
    .B(_5408__bF$buf4),
    .C(_5430_),
    .Y(_4639_)
);

NOR2X1 _15771_ (
    .A(\datapath.registers.838[5] [22]),
    .B(_5408__bF$buf3),
    .Y(_5431_)
);

AOI21X1 _15772_ (
    .A(_4843__bF$buf4),
    .B(_5408__bF$buf2),
    .C(_5431_),
    .Y(_4640_)
);

NOR2X1 _15773_ (
    .A(\datapath.registers.838[5] [23]),
    .B(_5408__bF$buf1),
    .Y(_5432_)
);

AOI21X1 _15774_ (
    .A(_4845__bF$buf4),
    .B(_5408__bF$buf0),
    .C(_5432_),
    .Y(_4641_)
);

NOR2X1 _15775_ (
    .A(\datapath.registers.838[5] [24]),
    .B(_5408__bF$buf7),
    .Y(_5433_)
);

AOI21X1 _15776_ (
    .A(_4847__bF$buf1),
    .B(_5408__bF$buf6),
    .C(_5433_),
    .Y(_4642_)
);

NOR2X1 _15777_ (
    .A(\datapath.registers.838[5] [25]),
    .B(_5408__bF$buf5),
    .Y(_5434_)
);

AOI21X1 _15778_ (
    .A(_4849__bF$buf4),
    .B(_5408__bF$buf4),
    .C(_5434_),
    .Y(_4643_)
);

NOR2X1 _15779_ (
    .A(\datapath.registers.838[5] [26]),
    .B(_5408__bF$buf3),
    .Y(_5435_)
);

AOI21X1 _15780_ (
    .A(_4851__bF$buf3),
    .B(_5408__bF$buf2),
    .C(_5435_),
    .Y(_4644_)
);

NOR2X1 _15781_ (
    .A(\datapath.registers.838[5] [27]),
    .B(_5408__bF$buf1),
    .Y(_5436_)
);

AOI21X1 _15782_ (
    .A(_4853__bF$buf4),
    .B(_5408__bF$buf0),
    .C(_5436_),
    .Y(_4645_)
);

NOR2X1 _15783_ (
    .A(\datapath.registers.838[5] [28]),
    .B(_5408__bF$buf7),
    .Y(_5437_)
);

AOI21X1 _15784_ (
    .A(_4855__bF$buf3),
    .B(_5408__bF$buf6),
    .C(_5437_),
    .Y(_4646_)
);

NOR2X1 _15785_ (
    .A(\datapath.registers.838[5] [29]),
    .B(_5408__bF$buf5),
    .Y(_5438_)
);

AOI21X1 _15786_ (
    .A(_4857__bF$buf3),
    .B(_5408__bF$buf4),
    .C(_5438_),
    .Y(_4647_)
);

NOR2X1 _15787_ (
    .A(\datapath.registers.838[5] [30]),
    .B(_5408__bF$buf3),
    .Y(_5439_)
);

AOI21X1 _15788_ (
    .A(_4859__bF$buf0),
    .B(_5408__bF$buf2),
    .C(_5439_),
    .Y(_4649_)
);

NOR2X1 _15789_ (
    .A(\datapath.registers.838[5] [31]),
    .B(_5408__bF$buf1),
    .Y(_5440_)
);

AOI21X1 _15790_ (
    .A(_4861__bF$buf3),
    .B(_5408__bF$buf0),
    .C(_5440_),
    .Y(_4650_)
);

NOR2X1 _15791_ (
    .A(_5341__bF$buf0),
    .B(_4790_),
    .Y(_5441_)
);

NAND2X1 _15792_ (
    .A(_5441_),
    .B(_5015_),
    .Y(_5442_)
);

NAND2X1 _15793_ (
    .A(\datapath.registers.838[4] [0]),
    .B(_5442__bF$buf7),
    .Y(_5443_)
);

OAI21X1 _15794_ (
    .A(_4786__bF$buf4),
    .B(_5442__bF$buf6),
    .C(_5443_),
    .Y(_4594_)
);

NAND2X1 _15795_ (
    .A(\datapath.registers.838[4] [1]),
    .B(_5442__bF$buf5),
    .Y(_5444_)
);

OAI21X1 _15796_ (
    .A(_4801__bF$buf2),
    .B(_5442__bF$buf4),
    .C(_5444_),
    .Y(_4605_)
);

NAND2X1 _15797_ (
    .A(\datapath.registers.838[4] [2]),
    .B(_5442__bF$buf3),
    .Y(_5445_)
);

OAI21X1 _15798_ (
    .A(_4803__bF$buf4),
    .B(_5442__bF$buf2),
    .C(_5445_),
    .Y(_4616_)
);

NAND2X1 _15799_ (
    .A(\datapath.registers.838[4] [3]),
    .B(_5442__bF$buf1),
    .Y(_5446_)
);

OAI21X1 _15800_ (
    .A(_4805__bF$buf0),
    .B(_5442__bF$buf0),
    .C(_5446_),
    .Y(_4619_)
);

NAND2X1 _15801_ (
    .A(\datapath.registers.838[4] [4]),
    .B(_5442__bF$buf7),
    .Y(_5447_)
);

OAI21X1 _15802_ (
    .A(_4807__bF$buf3),
    .B(_5442__bF$buf6),
    .C(_5447_),
    .Y(_4620_)
);

NAND2X1 _15803_ (
    .A(\datapath.registers.838[4] [5]),
    .B(_5442__bF$buf5),
    .Y(_5448_)
);

OAI21X1 _15804_ (
    .A(_4809__bF$buf3),
    .B(_5442__bF$buf4),
    .C(_5448_),
    .Y(_4621_)
);

NAND2X1 _15805_ (
    .A(\datapath.registers.838[4] [6]),
    .B(_5442__bF$buf3),
    .Y(_5449_)
);

OAI21X1 _15806_ (
    .A(_4811__bF$buf0),
    .B(_5442__bF$buf2),
    .C(_5449_),
    .Y(_4622_)
);

NAND2X1 _15807_ (
    .A(\datapath.registers.838[4] [7]),
    .B(_5442__bF$buf1),
    .Y(_5450_)
);

OAI21X1 _15808_ (
    .A(_4813__bF$buf2),
    .B(_5442__bF$buf0),
    .C(_5450_),
    .Y(_4623_)
);

NAND2X1 _15809_ (
    .A(\datapath.registers.838[4] [8]),
    .B(_5442__bF$buf7),
    .Y(_5451_)
);

OAI21X1 _15810_ (
    .A(_4815__bF$buf2),
    .B(_5442__bF$buf6),
    .C(_5451_),
    .Y(_4624_)
);

NAND2X1 _15811_ (
    .A(\datapath.registers.838[4] [9]),
    .B(_5442__bF$buf5),
    .Y(_5452_)
);

OAI21X1 _15812_ (
    .A(_4817__bF$buf0),
    .B(_5442__bF$buf4),
    .C(_5452_),
    .Y(_4625_)
);

NAND2X1 _15813_ (
    .A(\datapath.registers.838[4] [10]),
    .B(_5442__bF$buf3),
    .Y(_5453_)
);

OAI21X1 _15814_ (
    .A(_4819__bF$buf3),
    .B(_5442__bF$buf2),
    .C(_5453_),
    .Y(_4595_)
);

NAND2X1 _15815_ (
    .A(\datapath.registers.838[4] [11]),
    .B(_5442__bF$buf1),
    .Y(_5454_)
);

OAI21X1 _15816_ (
    .A(_4821__bF$buf2),
    .B(_5442__bF$buf0),
    .C(_5454_),
    .Y(_4596_)
);

NAND2X1 _15817_ (
    .A(\datapath.registers.838[4] [12]),
    .B(_5442__bF$buf7),
    .Y(_5455_)
);

OAI21X1 _15818_ (
    .A(_4823__bF$buf4),
    .B(_5442__bF$buf6),
    .C(_5455_),
    .Y(_4597_)
);

NAND2X1 _15819_ (
    .A(\datapath.registers.838[4] [13]),
    .B(_5442__bF$buf5),
    .Y(_5456_)
);

OAI21X1 _15820_ (
    .A(_4825__bF$buf2),
    .B(_5442__bF$buf4),
    .C(_5456_),
    .Y(_4598_)
);

NAND2X1 _15821_ (
    .A(\datapath.registers.838[4] [14]),
    .B(_5442__bF$buf3),
    .Y(_5457_)
);

OAI21X1 _15822_ (
    .A(_4827__bF$buf2),
    .B(_5442__bF$buf2),
    .C(_5457_),
    .Y(_4599_)
);

NAND2X1 _15823_ (
    .A(\datapath.registers.838[4] [15]),
    .B(_5442__bF$buf1),
    .Y(_5458_)
);

OAI21X1 _15824_ (
    .A(_4829__bF$buf2),
    .B(_5442__bF$buf0),
    .C(_5458_),
    .Y(_4600_)
);

NAND2X1 _15825_ (
    .A(\datapath.registers.838[4] [16]),
    .B(_5442__bF$buf7),
    .Y(_5459_)
);

OAI21X1 _15826_ (
    .A(_4831__bF$buf2),
    .B(_5442__bF$buf6),
    .C(_5459_),
    .Y(_4601_)
);

NAND2X1 _15827_ (
    .A(\datapath.registers.838[4] [17]),
    .B(_5442__bF$buf5),
    .Y(_5460_)
);

OAI21X1 _15828_ (
    .A(_4833__bF$buf4),
    .B(_5442__bF$buf4),
    .C(_5460_),
    .Y(_4602_)
);

NAND2X1 _15829_ (
    .A(\datapath.registers.838[4] [18]),
    .B(_5442__bF$buf3),
    .Y(_5461_)
);

OAI21X1 _15830_ (
    .A(_4835__bF$buf4),
    .B(_5442__bF$buf2),
    .C(_5461_),
    .Y(_4603_)
);

NAND2X1 _15831_ (
    .A(\datapath.registers.838[4] [19]),
    .B(_5442__bF$buf1),
    .Y(_5462_)
);

OAI21X1 _15832_ (
    .A(_4837__bF$buf0),
    .B(_5442__bF$buf0),
    .C(_5462_),
    .Y(_4604_)
);

NAND2X1 _15833_ (
    .A(\datapath.registers.838[4] [20]),
    .B(_5442__bF$buf7),
    .Y(_5463_)
);

OAI21X1 _15834_ (
    .A(_4839__bF$buf2),
    .B(_5442__bF$buf6),
    .C(_5463_),
    .Y(_4606_)
);

NAND2X1 _15835_ (
    .A(\datapath.registers.838[4] [21]),
    .B(_5442__bF$buf5),
    .Y(_5464_)
);

OAI21X1 _15836_ (
    .A(_4841__bF$buf3),
    .B(_5442__bF$buf4),
    .C(_5464_),
    .Y(_4607_)
);

NAND2X1 _15837_ (
    .A(\datapath.registers.838[4] [22]),
    .B(_5442__bF$buf3),
    .Y(_5465_)
);

OAI21X1 _15838_ (
    .A(_4843__bF$buf3),
    .B(_5442__bF$buf2),
    .C(_5465_),
    .Y(_4608_)
);

NAND2X1 _15839_ (
    .A(\datapath.registers.838[4] [23]),
    .B(_5442__bF$buf1),
    .Y(_5466_)
);

OAI21X1 _15840_ (
    .A(_4845__bF$buf3),
    .B(_5442__bF$buf0),
    .C(_5466_),
    .Y(_4609_)
);

NAND2X1 _15841_ (
    .A(\datapath.registers.838[4] [24]),
    .B(_5442__bF$buf7),
    .Y(_5467_)
);

OAI21X1 _15842_ (
    .A(_4847__bF$buf0),
    .B(_5442__bF$buf6),
    .C(_5467_),
    .Y(_4610_)
);

NAND2X1 _15843_ (
    .A(\datapath.registers.838[4] [25]),
    .B(_5442__bF$buf5),
    .Y(_5468_)
);

OAI21X1 _15844_ (
    .A(_4849__bF$buf3),
    .B(_5442__bF$buf4),
    .C(_5468_),
    .Y(_4611_)
);

NAND2X1 _15845_ (
    .A(\datapath.registers.838[4] [26]),
    .B(_5442__bF$buf3),
    .Y(_5469_)
);

OAI21X1 _15846_ (
    .A(_4851__bF$buf2),
    .B(_5442__bF$buf2),
    .C(_5469_),
    .Y(_4612_)
);

NAND2X1 _15847_ (
    .A(\datapath.registers.838[4] [27]),
    .B(_5442__bF$buf1),
    .Y(_5470_)
);

OAI21X1 _15848_ (
    .A(_4853__bF$buf3),
    .B(_5442__bF$buf0),
    .C(_5470_),
    .Y(_4613_)
);

NAND2X1 _15849_ (
    .A(\datapath.registers.838[4] [28]),
    .B(_5442__bF$buf7),
    .Y(_5471_)
);

OAI21X1 _15850_ (
    .A(_4855__bF$buf2),
    .B(_5442__bF$buf6),
    .C(_5471_),
    .Y(_4614_)
);

NAND2X1 _15851_ (
    .A(\datapath.registers.838[4] [29]),
    .B(_5442__bF$buf5),
    .Y(_5472_)
);

OAI21X1 _15852_ (
    .A(_4857__bF$buf2),
    .B(_5442__bF$buf4),
    .C(_5472_),
    .Y(_4615_)
);

NAND2X1 _15853_ (
    .A(\datapath.registers.838[4] [30]),
    .B(_5442__bF$buf3),
    .Y(_5473_)
);

OAI21X1 _15854_ (
    .A(_4859__bF$buf4),
    .B(_5442__bF$buf2),
    .C(_5473_),
    .Y(_4617_)
);

NAND2X1 _15855_ (
    .A(\datapath.registers.838[4] [31]),
    .B(_5442__bF$buf1),
    .Y(_5474_)
);

OAI21X1 _15856_ (
    .A(_4861__bF$buf2),
    .B(_5442__bF$buf0),
    .C(_5474_),
    .Y(_4618_)
);

NAND2X1 _15857_ (
    .A(\datapath.wbinstr [10]),
    .B(\datapath.wbinstr [11]),
    .Y(_5475_)
);

NOR2X1 _15858_ (
    .A(\datapath.wbinstr [9]),
    .B(_5475_),
    .Y(_5476_)
);

NAND3X1 _15859_ (
    .A(_4789_),
    .B(_5476_),
    .C(_5015_),
    .Y(_5477_)
);

NAND2X1 _15860_ (
    .A(\datapath.registers.838[24] [0]),
    .B(_5477__bF$buf7),
    .Y(_5478_)
);

OAI21X1 _15861_ (
    .A(_4786__bF$buf3),
    .B(_5477__bF$buf6),
    .C(_5478_),
    .Y(_4274_)
);

NAND2X1 _15862_ (
    .A(\datapath.registers.838[24] [1]),
    .B(_5477__bF$buf5),
    .Y(_5479_)
);

OAI21X1 _15863_ (
    .A(_4801__bF$buf1),
    .B(_5477__bF$buf4),
    .C(_5479_),
    .Y(_4285_)
);

NAND2X1 _15864_ (
    .A(\datapath.registers.838[24] [2]),
    .B(_5477__bF$buf3),
    .Y(_5480_)
);

OAI21X1 _15865_ (
    .A(_4803__bF$buf3),
    .B(_5477__bF$buf2),
    .C(_5480_),
    .Y(_4296_)
);

NAND2X1 _15866_ (
    .A(\datapath.registers.838[24] [3]),
    .B(_5477__bF$buf1),
    .Y(_5481_)
);

OAI21X1 _15867_ (
    .A(_4805__bF$buf4),
    .B(_5477__bF$buf0),
    .C(_5481_),
    .Y(_4299_)
);

NAND2X1 _15868_ (
    .A(\datapath.registers.838[24] [4]),
    .B(_5477__bF$buf7),
    .Y(_5482_)
);

OAI21X1 _15869_ (
    .A(_4807__bF$buf2),
    .B(_5477__bF$buf6),
    .C(_5482_),
    .Y(_4300_)
);

NAND2X1 _15870_ (
    .A(\datapath.registers.838[24] [5]),
    .B(_5477__bF$buf5),
    .Y(_5483_)
);

OAI21X1 _15871_ (
    .A(_4809__bF$buf2),
    .B(_5477__bF$buf4),
    .C(_5483_),
    .Y(_4301_)
);

NAND2X1 _15872_ (
    .A(\datapath.registers.838[24] [6]),
    .B(_5477__bF$buf3),
    .Y(_5484_)
);

OAI21X1 _15873_ (
    .A(_4811__bF$buf4),
    .B(_5477__bF$buf2),
    .C(_5484_),
    .Y(_4302_)
);

NAND2X1 _15874_ (
    .A(\datapath.registers.838[24] [7]),
    .B(_5477__bF$buf1),
    .Y(_5485_)
);

OAI21X1 _15875_ (
    .A(_4813__bF$buf1),
    .B(_5477__bF$buf0),
    .C(_5485_),
    .Y(_4303_)
);

NAND2X1 _15876_ (
    .A(\datapath.registers.838[24] [8]),
    .B(_5477__bF$buf7),
    .Y(_5486_)
);

OAI21X1 _15877_ (
    .A(_4815__bF$buf1),
    .B(_5477__bF$buf6),
    .C(_5486_),
    .Y(_4304_)
);

NAND2X1 _15878_ (
    .A(\datapath.registers.838[24] [9]),
    .B(_5477__bF$buf5),
    .Y(_5487_)
);

OAI21X1 _15879_ (
    .A(_4817__bF$buf4),
    .B(_5477__bF$buf4),
    .C(_5487_),
    .Y(_4305_)
);

NAND2X1 _15880_ (
    .A(\datapath.registers.838[24] [10]),
    .B(_5477__bF$buf3),
    .Y(_5488_)
);

OAI21X1 _15881_ (
    .A(_4819__bF$buf2),
    .B(_5477__bF$buf2),
    .C(_5488_),
    .Y(_4275_)
);

NAND2X1 _15882_ (
    .A(\datapath.registers.838[24] [11]),
    .B(_5477__bF$buf1),
    .Y(_5489_)
);

OAI21X1 _15883_ (
    .A(_4821__bF$buf1),
    .B(_5477__bF$buf0),
    .C(_5489_),
    .Y(_4276_)
);

NAND2X1 _15884_ (
    .A(\datapath.registers.838[24] [12]),
    .B(_5477__bF$buf7),
    .Y(_5490_)
);

OAI21X1 _15885_ (
    .A(_4823__bF$buf3),
    .B(_5477__bF$buf6),
    .C(_5490_),
    .Y(_4277_)
);

NAND2X1 _15886_ (
    .A(\datapath.registers.838[24] [13]),
    .B(_5477__bF$buf5),
    .Y(_5491_)
);

OAI21X1 _15887_ (
    .A(_4825__bF$buf1),
    .B(_5477__bF$buf4),
    .C(_5491_),
    .Y(_4278_)
);

NAND2X1 _15888_ (
    .A(\datapath.registers.838[24] [14]),
    .B(_5477__bF$buf3),
    .Y(_5492_)
);

OAI21X1 _15889_ (
    .A(_4827__bF$buf1),
    .B(_5477__bF$buf2),
    .C(_5492_),
    .Y(_4279_)
);

NAND2X1 _15890_ (
    .A(\datapath.registers.838[24] [15]),
    .B(_5477__bF$buf1),
    .Y(_5493_)
);

OAI21X1 _15891_ (
    .A(_4829__bF$buf1),
    .B(_5477__bF$buf0),
    .C(_5493_),
    .Y(_4280_)
);

NAND2X1 _15892_ (
    .A(\datapath.registers.838[24] [16]),
    .B(_5477__bF$buf7),
    .Y(_5494_)
);

OAI21X1 _15893_ (
    .A(_4831__bF$buf1),
    .B(_5477__bF$buf6),
    .C(_5494_),
    .Y(_4281_)
);

NAND2X1 _15894_ (
    .A(\datapath.registers.838[24] [17]),
    .B(_5477__bF$buf5),
    .Y(_5495_)
);

OAI21X1 _15895_ (
    .A(_4833__bF$buf3),
    .B(_5477__bF$buf4),
    .C(_5495_),
    .Y(_4282_)
);

NAND2X1 _15896_ (
    .A(\datapath.registers.838[24] [18]),
    .B(_5477__bF$buf3),
    .Y(_5496_)
);

OAI21X1 _15897_ (
    .A(_4835__bF$buf3),
    .B(_5477__bF$buf2),
    .C(_5496_),
    .Y(_4283_)
);

NAND2X1 _15898_ (
    .A(\datapath.registers.838[24] [19]),
    .B(_5477__bF$buf1),
    .Y(_5497_)
);

OAI21X1 _15899_ (
    .A(_4837__bF$buf4),
    .B(_5477__bF$buf0),
    .C(_5497_),
    .Y(_4284_)
);

NAND2X1 _15900_ (
    .A(\datapath.registers.838[24] [20]),
    .B(_5477__bF$buf7),
    .Y(_5498_)
);

OAI21X1 _15901_ (
    .A(_4839__bF$buf1),
    .B(_5477__bF$buf6),
    .C(_5498_),
    .Y(_4286_)
);

NAND2X1 _15902_ (
    .A(\datapath.registers.838[24] [21]),
    .B(_5477__bF$buf5),
    .Y(_5499_)
);

OAI21X1 _15903_ (
    .A(_4841__bF$buf2),
    .B(_5477__bF$buf4),
    .C(_5499_),
    .Y(_4287_)
);

NAND2X1 _15904_ (
    .A(\datapath.registers.838[24] [22]),
    .B(_5477__bF$buf3),
    .Y(_5500_)
);

OAI21X1 _15905_ (
    .A(_4843__bF$buf2),
    .B(_5477__bF$buf2),
    .C(_5500_),
    .Y(_4288_)
);

NAND2X1 _15906_ (
    .A(\datapath.registers.838[24] [23]),
    .B(_5477__bF$buf1),
    .Y(_5501_)
);

OAI21X1 _15907_ (
    .A(_4845__bF$buf2),
    .B(_5477__bF$buf0),
    .C(_5501_),
    .Y(_4289_)
);

NAND2X1 _15908_ (
    .A(\datapath.registers.838[24] [24]),
    .B(_5477__bF$buf7),
    .Y(_5502_)
);

OAI21X1 _15909_ (
    .A(_4847__bF$buf4),
    .B(_5477__bF$buf6),
    .C(_5502_),
    .Y(_4290_)
);

NAND2X1 _15910_ (
    .A(\datapath.registers.838[24] [25]),
    .B(_5477__bF$buf5),
    .Y(_5503_)
);

OAI21X1 _15911_ (
    .A(_4849__bF$buf2),
    .B(_5477__bF$buf4),
    .C(_5503_),
    .Y(_4291_)
);

NAND2X1 _15912_ (
    .A(\datapath.registers.838[24] [26]),
    .B(_5477__bF$buf3),
    .Y(_5504_)
);

OAI21X1 _15913_ (
    .A(_4851__bF$buf1),
    .B(_5477__bF$buf2),
    .C(_5504_),
    .Y(_4292_)
);

NAND2X1 _15914_ (
    .A(\datapath.registers.838[24] [27]),
    .B(_5477__bF$buf1),
    .Y(_5505_)
);

OAI21X1 _15915_ (
    .A(_4853__bF$buf2),
    .B(_5477__bF$buf0),
    .C(_5505_),
    .Y(_4293_)
);

NAND2X1 _15916_ (
    .A(\datapath.registers.838[24] [28]),
    .B(_5477__bF$buf7),
    .Y(_5506_)
);

OAI21X1 _15917_ (
    .A(_4855__bF$buf1),
    .B(_5477__bF$buf6),
    .C(_5506_),
    .Y(_4294_)
);

NAND2X1 _15918_ (
    .A(\datapath.registers.838[24] [29]),
    .B(_5477__bF$buf5),
    .Y(_5507_)
);

OAI21X1 _15919_ (
    .A(_4857__bF$buf1),
    .B(_5477__bF$buf4),
    .C(_5507_),
    .Y(_4295_)
);

NAND2X1 _15920_ (
    .A(\datapath.registers.838[24] [30]),
    .B(_5477__bF$buf3),
    .Y(_5508_)
);

OAI21X1 _15921_ (
    .A(_4859__bF$buf3),
    .B(_5477__bF$buf2),
    .C(_5508_),
    .Y(_4297_)
);

NAND2X1 _15922_ (
    .A(\datapath.registers.838[24] [31]),
    .B(_5477__bF$buf1),
    .Y(_5509_)
);

OAI21X1 _15923_ (
    .A(_4861__bF$buf1),
    .B(_5477__bF$buf0),
    .C(_5509_),
    .Y(_4298_)
);

NOR2X1 _15924_ (
    .A(_4794__bF$buf6),
    .B(_4899__bF$buf7),
    .Y(_5510_)
);

NOR2X1 _15925_ (
    .A(\datapath.registers.838[3] [0]),
    .B(_5510__bF$buf7),
    .Y(_5511_)
);

AOI21X1 _15926_ (
    .A(_4786__bF$buf2),
    .B(_5510__bF$buf6),
    .C(_5511_),
    .Y(_4562_)
);

NOR2X1 _15927_ (
    .A(\datapath.registers.838[3] [1]),
    .B(_5510__bF$buf5),
    .Y(_5512_)
);

AOI21X1 _15928_ (
    .A(_4801__bF$buf0),
    .B(_5510__bF$buf4),
    .C(_5512_),
    .Y(_4573_)
);

NOR2X1 _15929_ (
    .A(\datapath.registers.838[3] [2]),
    .B(_5510__bF$buf3),
    .Y(_5513_)
);

AOI21X1 _15930_ (
    .A(_4803__bF$buf2),
    .B(_5510__bF$buf2),
    .C(_5513_),
    .Y(_4584_)
);

NOR2X1 _15931_ (
    .A(\datapath.registers.838[3] [3]),
    .B(_5510__bF$buf1),
    .Y(_5514_)
);

AOI21X1 _15932_ (
    .A(_4805__bF$buf3),
    .B(_5510__bF$buf0),
    .C(_5514_),
    .Y(_4587_)
);

NOR2X1 _15933_ (
    .A(\datapath.registers.838[3] [4]),
    .B(_5510__bF$buf7),
    .Y(_5515_)
);

AOI21X1 _15934_ (
    .A(_4807__bF$buf1),
    .B(_5510__bF$buf6),
    .C(_5515_),
    .Y(_4588_)
);

NOR2X1 _15935_ (
    .A(\datapath.registers.838[3] [5]),
    .B(_5510__bF$buf5),
    .Y(_5516_)
);

AOI21X1 _15936_ (
    .A(_4809__bF$buf1),
    .B(_5510__bF$buf4),
    .C(_5516_),
    .Y(_4589_)
);

NOR2X1 _15937_ (
    .A(\datapath.registers.838[3] [6]),
    .B(_5510__bF$buf3),
    .Y(_5517_)
);

AOI21X1 _15938_ (
    .A(_4811__bF$buf3),
    .B(_5510__bF$buf2),
    .C(_5517_),
    .Y(_4590_)
);

NOR2X1 _15939_ (
    .A(\datapath.registers.838[3] [7]),
    .B(_5510__bF$buf1),
    .Y(_5518_)
);

AOI21X1 _15940_ (
    .A(_4813__bF$buf0),
    .B(_5510__bF$buf0),
    .C(_5518_),
    .Y(_4591_)
);

INVX1 _15941_ (
    .A(\datapath.registers.838[3] [8]),
    .Y(_5519_)
);

NAND2X1 _15942_ (
    .A(\datapath.rd [8]),
    .B(_5510__bF$buf7),
    .Y(_5520_)
);

OAI21X1 _15943_ (
    .A(_5519_),
    .B(_5510__bF$buf6),
    .C(_5520_),
    .Y(_4592_)
);

INVX1 _15944_ (
    .A(\datapath.registers.838[3] [9]),
    .Y(_5521_)
);

NAND2X1 _15945_ (
    .A(\datapath.rd [9]),
    .B(_5510__bF$buf5),
    .Y(_5522_)
);

OAI21X1 _15946_ (
    .A(_5521_),
    .B(_5510__bF$buf4),
    .C(_5522_),
    .Y(_4593_)
);

INVX1 _15947_ (
    .A(\datapath.registers.838[3] [10]),
    .Y(_5523_)
);

NAND2X1 _15948_ (
    .A(\datapath.rd [10]),
    .B(_5510__bF$buf3),
    .Y(_5524_)
);

OAI21X1 _15949_ (
    .A(_5523_),
    .B(_5510__bF$buf2),
    .C(_5524_),
    .Y(_4563_)
);

NOR2X1 _15950_ (
    .A(\datapath.registers.838[3] [11]),
    .B(_5510__bF$buf1),
    .Y(_5525_)
);

AOI21X1 _15951_ (
    .A(_4821__bF$buf0),
    .B(_5510__bF$buf0),
    .C(_5525_),
    .Y(_4564_)
);

INVX1 _15952_ (
    .A(\datapath.registers.838[3] [12]),
    .Y(_5526_)
);

NAND2X1 _15953_ (
    .A(\datapath.rd [12]),
    .B(_5510__bF$buf7),
    .Y(_5527_)
);

OAI21X1 _15954_ (
    .A(_5526_),
    .B(_5510__bF$buf6),
    .C(_5527_),
    .Y(_4565_)
);

NOR2X1 _15955_ (
    .A(\datapath.registers.838[3] [13]),
    .B(_5510__bF$buf5),
    .Y(_5528_)
);

AOI21X1 _15956_ (
    .A(_4825__bF$buf0),
    .B(_5510__bF$buf4),
    .C(_5528_),
    .Y(_4566_)
);

NOR2X1 _15957_ (
    .A(\datapath.registers.838[3] [14]),
    .B(_5510__bF$buf3),
    .Y(_5529_)
);

AOI21X1 _15958_ (
    .A(_4827__bF$buf0),
    .B(_5510__bF$buf2),
    .C(_5529_),
    .Y(_4567_)
);

NOR2X1 _15959_ (
    .A(\datapath.registers.838[3] [15]),
    .B(_5510__bF$buf1),
    .Y(_5530_)
);

AOI21X1 _15960_ (
    .A(_4829__bF$buf0),
    .B(_5510__bF$buf0),
    .C(_5530_),
    .Y(_4568_)
);

NOR2X1 _15961_ (
    .A(\datapath.registers.838[3] [16]),
    .B(_5510__bF$buf7),
    .Y(_5531_)
);

AOI21X1 _15962_ (
    .A(_4831__bF$buf0),
    .B(_5510__bF$buf6),
    .C(_5531_),
    .Y(_4569_)
);

NOR2X1 _15963_ (
    .A(\datapath.registers.838[3] [17]),
    .B(_5510__bF$buf5),
    .Y(_5532_)
);

AOI21X1 _15964_ (
    .A(_4833__bF$buf2),
    .B(_5510__bF$buf4),
    .C(_5532_),
    .Y(_4570_)
);

NOR2X1 _15965_ (
    .A(\datapath.registers.838[3] [18]),
    .B(_5510__bF$buf3),
    .Y(_5533_)
);

AOI21X1 _15966_ (
    .A(_4835__bF$buf2),
    .B(_5510__bF$buf2),
    .C(_5533_),
    .Y(_4571_)
);

NOR2X1 _15967_ (
    .A(\datapath.registers.838[3] [19]),
    .B(_5510__bF$buf1),
    .Y(_5534_)
);

AOI21X1 _15968_ (
    .A(_4837__bF$buf3),
    .B(_5510__bF$buf0),
    .C(_5534_),
    .Y(_4572_)
);

NOR2X1 _15969_ (
    .A(\datapath.registers.838[3] [20]),
    .B(_5510__bF$buf7),
    .Y(_5535_)
);

AOI21X1 _15970_ (
    .A(_4839__bF$buf0),
    .B(_5510__bF$buf6),
    .C(_5535_),
    .Y(_4574_)
);

INVX1 _15971_ (
    .A(\datapath.registers.838[3] [21]),
    .Y(_5536_)
);

NAND2X1 _15972_ (
    .A(\datapath.rd [21]),
    .B(_5510__bF$buf5),
    .Y(_5537_)
);

OAI21X1 _15973_ (
    .A(_5536_),
    .B(_5510__bF$buf4),
    .C(_5537_),
    .Y(_4575_)
);

NOR2X1 _15974_ (
    .A(\datapath.registers.838[3] [22]),
    .B(_5510__bF$buf3),
    .Y(_5538_)
);

AOI21X1 _15975_ (
    .A(_4843__bF$buf1),
    .B(_5510__bF$buf2),
    .C(_5538_),
    .Y(_4576_)
);

INVX1 _15976_ (
    .A(\datapath.registers.838[3] [23]),
    .Y(_5539_)
);

NAND2X1 _15977_ (
    .A(\datapath.rd [23]),
    .B(_5510__bF$buf1),
    .Y(_5540_)
);

OAI21X1 _15978_ (
    .A(_5539_),
    .B(_5510__bF$buf0),
    .C(_5540_),
    .Y(_4577_)
);

INVX1 _15979_ (
    .A(\datapath.registers.838[3] [24]),
    .Y(_5541_)
);

NAND2X1 _15980_ (
    .A(\datapath.rd [24]),
    .B(_5510__bF$buf7),
    .Y(_5542_)
);

OAI21X1 _15981_ (
    .A(_5541_),
    .B(_5510__bF$buf6),
    .C(_5542_),
    .Y(_4578_)
);

INVX1 _15982_ (
    .A(\datapath.registers.838[3] [25]),
    .Y(_5543_)
);

NAND2X1 _15983_ (
    .A(\datapath.rd [25]),
    .B(_5510__bF$buf5),
    .Y(_5544_)
);

OAI21X1 _15984_ (
    .A(_5543_),
    .B(_5510__bF$buf4),
    .C(_5544_),
    .Y(_4579_)
);

NOR2X1 _15985_ (
    .A(\datapath.registers.838[3] [26]),
    .B(_5510__bF$buf3),
    .Y(_5545_)
);

AOI21X1 _15986_ (
    .A(_4851__bF$buf0),
    .B(_5510__bF$buf2),
    .C(_5545_),
    .Y(_4580_)
);

NOR2X1 _15987_ (
    .A(\datapath.registers.838[3] [27]),
    .B(_5510__bF$buf1),
    .Y(_5546_)
);

AOI21X1 _15988_ (
    .A(_4853__bF$buf1),
    .B(_5510__bF$buf0),
    .C(_5546_),
    .Y(_4581_)
);

NOR2X1 _15989_ (
    .A(\datapath.registers.838[3] [28]),
    .B(_5510__bF$buf7),
    .Y(_5547_)
);

AOI21X1 _15990_ (
    .A(_4855__bF$buf0),
    .B(_5510__bF$buf6),
    .C(_5547_),
    .Y(_4582_)
);

NOR2X1 _15991_ (
    .A(\datapath.registers.838[3] [29]),
    .B(_5510__bF$buf5),
    .Y(_5548_)
);

AOI21X1 _15992_ (
    .A(_4857__bF$buf0),
    .B(_5510__bF$buf4),
    .C(_5548_),
    .Y(_4583_)
);

NOR2X1 _15993_ (
    .A(\datapath.registers.838[3] [30]),
    .B(_5510__bF$buf3),
    .Y(_5549_)
);

AOI21X1 _15994_ (
    .A(_4859__bF$buf2),
    .B(_5510__bF$buf2),
    .C(_5549_),
    .Y(_4585_)
);

NOR2X1 _15995_ (
    .A(\datapath.registers.838[3] [31]),
    .B(_5510__bF$buf1),
    .Y(_5550_)
);

AOI21X1 _15996_ (
    .A(_4861__bF$buf0),
    .B(_5510__bF$buf0),
    .C(_5550_),
    .Y(_4586_)
);

NAND2X1 _15997_ (
    .A(_4898_),
    .B(_4798_),
    .Y(_5551_)
);

NAND2X1 _15998_ (
    .A(\datapath.registers.838[23] [0]),
    .B(_5551__bF$buf7),
    .Y(_5552_)
);

OAI21X1 _15999_ (
    .A(_4786__bF$buf1),
    .B(_5551__bF$buf6),
    .C(_5552_),
    .Y(_4242_)
);

NAND2X1 _16000_ (
    .A(\datapath.registers.838[23] [1]),
    .B(_5551__bF$buf5),
    .Y(_5553_)
);

OAI21X1 _16001_ (
    .A(_4801__bF$buf4),
    .B(_5551__bF$buf4),
    .C(_5553_),
    .Y(_4253_)
);

NAND2X1 _16002_ (
    .A(\datapath.registers.838[23] [2]),
    .B(_5551__bF$buf3),
    .Y(_5554_)
);

OAI21X1 _16003_ (
    .A(_4803__bF$buf1),
    .B(_5551__bF$buf2),
    .C(_5554_),
    .Y(_4264_)
);

NAND2X1 _16004_ (
    .A(\datapath.registers.838[23] [3]),
    .B(_5551__bF$buf1),
    .Y(_5555_)
);

OAI21X1 _16005_ (
    .A(_4805__bF$buf2),
    .B(_5551__bF$buf0),
    .C(_5555_),
    .Y(_4267_)
);

NAND2X1 _16006_ (
    .A(\datapath.registers.838[23] [4]),
    .B(_5551__bF$buf7),
    .Y(_5556_)
);

OAI21X1 _16007_ (
    .A(_4807__bF$buf0),
    .B(_5551__bF$buf6),
    .C(_5556_),
    .Y(_4268_)
);

NAND2X1 _16008_ (
    .A(\datapath.registers.838[23] [5]),
    .B(_5551__bF$buf5),
    .Y(_5557_)
);

OAI21X1 _16009_ (
    .A(_4809__bF$buf0),
    .B(_5551__bF$buf4),
    .C(_5557_),
    .Y(_4269_)
);

NAND2X1 _16010_ (
    .A(\datapath.registers.838[23] [6]),
    .B(_5551__bF$buf3),
    .Y(_5558_)
);

OAI21X1 _16011_ (
    .A(_4811__bF$buf2),
    .B(_5551__bF$buf2),
    .C(_5558_),
    .Y(_4270_)
);

NAND2X1 _16012_ (
    .A(\datapath.registers.838[23] [7]),
    .B(_5551__bF$buf1),
    .Y(_5559_)
);

OAI21X1 _16013_ (
    .A(_4813__bF$buf4),
    .B(_5551__bF$buf0),
    .C(_5559_),
    .Y(_4271_)
);

NAND2X1 _16014_ (
    .A(\datapath.registers.838[23] [8]),
    .B(_5551__bF$buf7),
    .Y(_5560_)
);

OAI21X1 _16015_ (
    .A(_4815__bF$buf0),
    .B(_5551__bF$buf6),
    .C(_5560_),
    .Y(_4272_)
);

NAND2X1 _16016_ (
    .A(\datapath.registers.838[23] [9]),
    .B(_5551__bF$buf5),
    .Y(_5561_)
);

OAI21X1 _16017_ (
    .A(_4817__bF$buf3),
    .B(_5551__bF$buf4),
    .C(_5561_),
    .Y(_4273_)
);

NAND2X1 _16018_ (
    .A(\datapath.registers.838[23] [10]),
    .B(_5551__bF$buf3),
    .Y(_5562_)
);

OAI21X1 _16019_ (
    .A(_4819__bF$buf1),
    .B(_5551__bF$buf2),
    .C(_5562_),
    .Y(_4243_)
);

NAND2X1 _16020_ (
    .A(\datapath.registers.838[23] [11]),
    .B(_5551__bF$buf1),
    .Y(_5563_)
);

OAI21X1 _16021_ (
    .A(_4821__bF$buf4),
    .B(_5551__bF$buf0),
    .C(_5563_),
    .Y(_4244_)
);

NAND2X1 _16022_ (
    .A(\datapath.registers.838[23] [12]),
    .B(_5551__bF$buf7),
    .Y(_5564_)
);

OAI21X1 _16023_ (
    .A(_4823__bF$buf2),
    .B(_5551__bF$buf6),
    .C(_5564_),
    .Y(_4245_)
);

NAND2X1 _16024_ (
    .A(\datapath.registers.838[23] [13]),
    .B(_5551__bF$buf5),
    .Y(_5565_)
);

OAI21X1 _16025_ (
    .A(_4825__bF$buf4),
    .B(_5551__bF$buf4),
    .C(_5565_),
    .Y(_4246_)
);

NAND2X1 _16026_ (
    .A(\datapath.registers.838[23] [14]),
    .B(_5551__bF$buf3),
    .Y(_5566_)
);

OAI21X1 _16027_ (
    .A(_4827__bF$buf4),
    .B(_5551__bF$buf2),
    .C(_5566_),
    .Y(_4247_)
);

NAND2X1 _16028_ (
    .A(\datapath.registers.838[23] [15]),
    .B(_5551__bF$buf1),
    .Y(_5567_)
);

OAI21X1 _16029_ (
    .A(_4829__bF$buf4),
    .B(_5551__bF$buf0),
    .C(_5567_),
    .Y(_4248_)
);

NAND2X1 _16030_ (
    .A(\datapath.registers.838[23] [16]),
    .B(_5551__bF$buf7),
    .Y(_5568_)
);

OAI21X1 _16031_ (
    .A(_4831__bF$buf4),
    .B(_5551__bF$buf6),
    .C(_5568_),
    .Y(_4249_)
);

NAND2X1 _16032_ (
    .A(\datapath.registers.838[23] [17]),
    .B(_5551__bF$buf5),
    .Y(_5569_)
);

OAI21X1 _16033_ (
    .A(_4833__bF$buf1),
    .B(_5551__bF$buf4),
    .C(_5569_),
    .Y(_4250_)
);

NAND2X1 _16034_ (
    .A(\datapath.registers.838[23] [18]),
    .B(_5551__bF$buf3),
    .Y(_5570_)
);

OAI21X1 _16035_ (
    .A(_4835__bF$buf1),
    .B(_5551__bF$buf2),
    .C(_5570_),
    .Y(_4251_)
);

NAND2X1 _16036_ (
    .A(\datapath.registers.838[23] [19]),
    .B(_5551__bF$buf1),
    .Y(_5571_)
);

OAI21X1 _16037_ (
    .A(_4837__bF$buf2),
    .B(_5551__bF$buf0),
    .C(_5571_),
    .Y(_4252_)
);

NAND2X1 _16038_ (
    .A(\datapath.registers.838[23] [20]),
    .B(_5551__bF$buf7),
    .Y(_5572_)
);

OAI21X1 _16039_ (
    .A(_4839__bF$buf4),
    .B(_5551__bF$buf6),
    .C(_5572_),
    .Y(_4254_)
);

NAND2X1 _16040_ (
    .A(\datapath.registers.838[23] [21]),
    .B(_5551__bF$buf5),
    .Y(_5573_)
);

OAI21X1 _16041_ (
    .A(_4841__bF$buf1),
    .B(_5551__bF$buf4),
    .C(_5573_),
    .Y(_4255_)
);

NAND2X1 _16042_ (
    .A(\datapath.registers.838[23] [22]),
    .B(_5551__bF$buf3),
    .Y(_5574_)
);

OAI21X1 _16043_ (
    .A(_4843__bF$buf0),
    .B(_5551__bF$buf2),
    .C(_5574_),
    .Y(_4256_)
);

NAND2X1 _16044_ (
    .A(\datapath.registers.838[23] [23]),
    .B(_5551__bF$buf1),
    .Y(_5575_)
);

OAI21X1 _16045_ (
    .A(_4845__bF$buf1),
    .B(_5551__bF$buf0),
    .C(_5575_),
    .Y(_4257_)
);

NAND2X1 _16046_ (
    .A(\datapath.registers.838[23] [24]),
    .B(_5551__bF$buf7),
    .Y(_5576_)
);

OAI21X1 _16047_ (
    .A(_4847__bF$buf3),
    .B(_5551__bF$buf6),
    .C(_5576_),
    .Y(_4258_)
);

NAND2X1 _16048_ (
    .A(\datapath.registers.838[23] [25]),
    .B(_5551__bF$buf5),
    .Y(_5577_)
);

OAI21X1 _16049_ (
    .A(_4849__bF$buf1),
    .B(_5551__bF$buf4),
    .C(_5577_),
    .Y(_4259_)
);

NAND2X1 _16050_ (
    .A(\datapath.registers.838[23] [26]),
    .B(_5551__bF$buf3),
    .Y(_5578_)
);

OAI21X1 _16051_ (
    .A(_4851__bF$buf4),
    .B(_5551__bF$buf2),
    .C(_5578_),
    .Y(_4260_)
);

NAND2X1 _16052_ (
    .A(\datapath.registers.838[23] [27]),
    .B(_5551__bF$buf1),
    .Y(_5579_)
);

OAI21X1 _16053_ (
    .A(_4853__bF$buf0),
    .B(_5551__bF$buf0),
    .C(_5579_),
    .Y(_4261_)
);

NAND2X1 _16054_ (
    .A(\datapath.registers.838[23] [28]),
    .B(_5551__bF$buf7),
    .Y(_5580_)
);

OAI21X1 _16055_ (
    .A(_4855__bF$buf4),
    .B(_5551__bF$buf6),
    .C(_5580_),
    .Y(_4262_)
);

NAND2X1 _16056_ (
    .A(\datapath.registers.838[23] [29]),
    .B(_5551__bF$buf5),
    .Y(_5581_)
);

OAI21X1 _16057_ (
    .A(_4857__bF$buf4),
    .B(_5551__bF$buf4),
    .C(_5581_),
    .Y(_4263_)
);

NAND2X1 _16058_ (
    .A(\datapath.registers.838[23] [30]),
    .B(_5551__bF$buf3),
    .Y(_5582_)
);

OAI21X1 _16059_ (
    .A(_4859__bF$buf1),
    .B(_5551__bF$buf2),
    .C(_5582_),
    .Y(_4265_)
);

NAND2X1 _16060_ (
    .A(\datapath.registers.838[23] [31]),
    .B(_5551__bF$buf1),
    .Y(_5583_)
);

OAI21X1 _16061_ (
    .A(_4861__bF$buf4),
    .B(_5551__bF$buf0),
    .C(_5583_),
    .Y(_4266_)
);

INVX1 _16062_ (
    .A(_4794__bF$buf5),
    .Y(_5584_)
);

INVX1 _16063_ (
    .A(_4934__bF$buf5),
    .Y(_5585_)
);

NAND2X1 _16064_ (
    .A(_5584_),
    .B(_5585_),
    .Y(_5586_)
);

OAI21X1 _16065_ (
    .A(_4794__bF$buf4),
    .B(_4934__bF$buf4),
    .C(\datapath.registers.838[2] [0]),
    .Y(_5587_)
);

OAI21X1 _16066_ (
    .A(_4786__bF$buf0),
    .B(_5586__bF$buf4),
    .C(_5587_),
    .Y(_4466_)
);

OAI21X1 _16067_ (
    .A(_4794__bF$buf3),
    .B(_4934__bF$buf3),
    .C(\datapath.registers.838[2] [1]),
    .Y(_5588_)
);

OAI21X1 _16068_ (
    .A(_4801__bF$buf3),
    .B(_5586__bF$buf3),
    .C(_5588_),
    .Y(_4477_)
);

OAI21X1 _16069_ (
    .A(_4794__bF$buf2),
    .B(_4934__bF$buf2),
    .C(\datapath.registers.838[2] [2]),
    .Y(_5589_)
);

OAI21X1 _16070_ (
    .A(_4803__bF$buf0),
    .B(_5586__bF$buf2),
    .C(_5589_),
    .Y(_4488_)
);

OAI21X1 _16071_ (
    .A(_4794__bF$buf1),
    .B(_4934__bF$buf1),
    .C(\datapath.registers.838[2] [3]),
    .Y(_5590_)
);

OAI21X1 _16072_ (
    .A(_4805__bF$buf1),
    .B(_5586__bF$buf1),
    .C(_5590_),
    .Y(_4491_)
);

OAI21X1 _16073_ (
    .A(_4794__bF$buf0),
    .B(_4934__bF$buf0),
    .C(\datapath.registers.838[2] [4]),
    .Y(_5591_)
);

OAI21X1 _16074_ (
    .A(_4807__bF$buf4),
    .B(_5586__bF$buf0),
    .C(_5591_),
    .Y(_4492_)
);

OAI21X1 _16075_ (
    .A(_4794__bF$buf7),
    .B(_4934__bF$buf9),
    .C(\datapath.registers.838[2] [5]),
    .Y(_5592_)
);

OAI21X1 _16076_ (
    .A(_4809__bF$buf4),
    .B(_5586__bF$buf4),
    .C(_5592_),
    .Y(_4493_)
);

OAI21X1 _16077_ (
    .A(_4794__bF$buf6),
    .B(_4934__bF$buf8),
    .C(\datapath.registers.838[2] [6]),
    .Y(_5593_)
);

OAI21X1 _16078_ (
    .A(_4811__bF$buf1),
    .B(_5586__bF$buf3),
    .C(_5593_),
    .Y(_4494_)
);

OAI21X1 _16079_ (
    .A(_4794__bF$buf5),
    .B(_4934__bF$buf7),
    .C(\datapath.registers.838[2] [7]),
    .Y(_5594_)
);

OAI21X1 _16080_ (
    .A(_4813__bF$buf3),
    .B(_5586__bF$buf2),
    .C(_5594_),
    .Y(_4495_)
);

OAI21X1 _16081_ (
    .A(_4794__bF$buf4),
    .B(_4934__bF$buf6),
    .C(\datapath.registers.838[2] [8]),
    .Y(_5595_)
);

OAI21X1 _16082_ (
    .A(_4815__bF$buf4),
    .B(_5586__bF$buf1),
    .C(_5595_),
    .Y(_4496_)
);

OAI21X1 _16083_ (
    .A(_4794__bF$buf3),
    .B(_4934__bF$buf5),
    .C(\datapath.registers.838[2] [9]),
    .Y(_5596_)
);

OAI21X1 _16084_ (
    .A(_4817__bF$buf2),
    .B(_5586__bF$buf0),
    .C(_5596_),
    .Y(_4497_)
);

OAI21X1 _16085_ (
    .A(_4794__bF$buf2),
    .B(_4934__bF$buf4),
    .C(\datapath.registers.838[2] [10]),
    .Y(_5597_)
);

OAI21X1 _16086_ (
    .A(_4819__bF$buf0),
    .B(_5586__bF$buf4),
    .C(_5597_),
    .Y(_4467_)
);

OAI21X1 _16087_ (
    .A(_4794__bF$buf1),
    .B(_4934__bF$buf3),
    .C(\datapath.registers.838[2] [11]),
    .Y(_5598_)
);

OAI21X1 _16088_ (
    .A(_4821__bF$buf3),
    .B(_5586__bF$buf3),
    .C(_5598_),
    .Y(_4468_)
);

OAI21X1 _16089_ (
    .A(_4794__bF$buf0),
    .B(_4934__bF$buf2),
    .C(\datapath.registers.838[2] [12]),
    .Y(_5599_)
);

OAI21X1 _16090_ (
    .A(_4823__bF$buf1),
    .B(_5586__bF$buf2),
    .C(_5599_),
    .Y(_4469_)
);

OAI21X1 _16091_ (
    .A(_4794__bF$buf7),
    .B(_4934__bF$buf1),
    .C(\datapath.registers.838[2] [13]),
    .Y(_5600_)
);

OAI21X1 _16092_ (
    .A(_4825__bF$buf3),
    .B(_5586__bF$buf1),
    .C(_5600_),
    .Y(_4470_)
);

OAI21X1 _16093_ (
    .A(_4794__bF$buf6),
    .B(_4934__bF$buf0),
    .C(\datapath.registers.838[2] [14]),
    .Y(_5601_)
);

OAI21X1 _16094_ (
    .A(_4827__bF$buf3),
    .B(_5586__bF$buf0),
    .C(_5601_),
    .Y(_4471_)
);

OAI21X1 _16095_ (
    .A(_4794__bF$buf5),
    .B(_4934__bF$buf9),
    .C(\datapath.registers.838[2] [15]),
    .Y(_5602_)
);

OAI21X1 _16096_ (
    .A(_4829__bF$buf3),
    .B(_5586__bF$buf4),
    .C(_5602_),
    .Y(_4472_)
);

OAI21X1 _16097_ (
    .A(_4794__bF$buf4),
    .B(_4934__bF$buf8),
    .C(\datapath.registers.838[2] [16]),
    .Y(_5603_)
);

OAI21X1 _16098_ (
    .A(_4831__bF$buf3),
    .B(_5586__bF$buf3),
    .C(_5603_),
    .Y(_4473_)
);

OAI21X1 _16099_ (
    .A(_4794__bF$buf3),
    .B(_4934__bF$buf7),
    .C(\datapath.registers.838[2] [17]),
    .Y(_5604_)
);

OAI21X1 _16100_ (
    .A(_4833__bF$buf0),
    .B(_5586__bF$buf2),
    .C(_5604_),
    .Y(_4474_)
);

OAI21X1 _16101_ (
    .A(_4794__bF$buf2),
    .B(_4934__bF$buf6),
    .C(\datapath.registers.838[2] [18]),
    .Y(_5605_)
);

OAI21X1 _16102_ (
    .A(_4835__bF$buf0),
    .B(_5586__bF$buf1),
    .C(_5605_),
    .Y(_4475_)
);

OAI21X1 _16103_ (
    .A(_4794__bF$buf1),
    .B(_4934__bF$buf5),
    .C(\datapath.registers.838[2] [19]),
    .Y(_5606_)
);

OAI21X1 _16104_ (
    .A(_4837__bF$buf1),
    .B(_5586__bF$buf0),
    .C(_5606_),
    .Y(_4476_)
);

OAI21X1 _16105_ (
    .A(_4794__bF$buf0),
    .B(_4934__bF$buf4),
    .C(\datapath.registers.838[2] [20]),
    .Y(_5607_)
);

OAI21X1 _16106_ (
    .A(_4839__bF$buf3),
    .B(_5586__bF$buf4),
    .C(_5607_),
    .Y(_4478_)
);

OAI21X1 _16107_ (
    .A(_4794__bF$buf7),
    .B(_4934__bF$buf3),
    .C(\datapath.registers.838[2] [21]),
    .Y(_5608_)
);

OAI21X1 _16108_ (
    .A(_4841__bF$buf0),
    .B(_5586__bF$buf3),
    .C(_5608_),
    .Y(_4479_)
);

OAI21X1 _16109_ (
    .A(_4794__bF$buf6),
    .B(_4934__bF$buf2),
    .C(\datapath.registers.838[2] [22]),
    .Y(_5609_)
);

OAI21X1 _16110_ (
    .A(_4843__bF$buf4),
    .B(_5586__bF$buf2),
    .C(_5609_),
    .Y(_4480_)
);

OAI21X1 _16111_ (
    .A(_4794__bF$buf5),
    .B(_4934__bF$buf1),
    .C(\datapath.registers.838[2] [23]),
    .Y(_5610_)
);

OAI21X1 _16112_ (
    .A(_4845__bF$buf0),
    .B(_5586__bF$buf1),
    .C(_5610_),
    .Y(_4481_)
);

OAI21X1 _16113_ (
    .A(_4794__bF$buf4),
    .B(_4934__bF$buf0),
    .C(\datapath.registers.838[2] [24]),
    .Y(_5611_)
);

OAI21X1 _16114_ (
    .A(_4847__bF$buf2),
    .B(_5586__bF$buf0),
    .C(_5611_),
    .Y(_4482_)
);

OAI21X1 _16115_ (
    .A(_4794__bF$buf3),
    .B(_4934__bF$buf9),
    .C(\datapath.registers.838[2] [25]),
    .Y(_5612_)
);

OAI21X1 _16116_ (
    .A(_4849__bF$buf0),
    .B(_5586__bF$buf4),
    .C(_5612_),
    .Y(_4483_)
);

OAI21X1 _16117_ (
    .A(_4794__bF$buf2),
    .B(_4934__bF$buf8),
    .C(\datapath.registers.838[2] [26]),
    .Y(_5613_)
);

OAI21X1 _16118_ (
    .A(_4851__bF$buf3),
    .B(_5586__bF$buf3),
    .C(_5613_),
    .Y(_4484_)
);

OAI21X1 _16119_ (
    .A(_4794__bF$buf1),
    .B(_4934__bF$buf7),
    .C(\datapath.registers.838[2] [27]),
    .Y(_5614_)
);

OAI21X1 _16120_ (
    .A(_4853__bF$buf4),
    .B(_5586__bF$buf2),
    .C(_5614_),
    .Y(_4485_)
);

OAI21X1 _16121_ (
    .A(_4794__bF$buf0),
    .B(_4934__bF$buf6),
    .C(\datapath.registers.838[2] [28]),
    .Y(_5615_)
);

OAI21X1 _16122_ (
    .A(_4855__bF$buf3),
    .B(_5586__bF$buf1),
    .C(_5615_),
    .Y(_4486_)
);

OAI21X1 _16123_ (
    .A(_4794__bF$buf7),
    .B(_4934__bF$buf5),
    .C(\datapath.registers.838[2] [29]),
    .Y(_5616_)
);

OAI21X1 _16124_ (
    .A(_4857__bF$buf3),
    .B(_5586__bF$buf0),
    .C(_5616_),
    .Y(_4487_)
);

OAI21X1 _16125_ (
    .A(_4794__bF$buf6),
    .B(_4934__bF$buf4),
    .C(\datapath.registers.838[2] [30]),
    .Y(_5617_)
);

OAI21X1 _16126_ (
    .A(_4859__bF$buf0),
    .B(_5586__bF$buf4),
    .C(_5617_),
    .Y(_4489_)
);

OAI21X1 _16127_ (
    .A(_4794__bF$buf5),
    .B(_4934__bF$buf3),
    .C(\datapath.registers.838[2] [31]),
    .Y(_5618_)
);

OAI21X1 _16128_ (
    .A(_4861__bF$buf3),
    .B(_5586__bF$buf3),
    .C(_5618_),
    .Y(_4490_)
);

INVX1 _16129_ (
    .A(_4968__bF$buf5),
    .Y(_5619_)
);

NAND2X1 _16130_ (
    .A(_5584_),
    .B(_5619_),
    .Y(_5620_)
);

OAI21X1 _16131_ (
    .A(_4794__bF$buf4),
    .B(_4968__bF$buf4),
    .C(\datapath.registers.838[1] [0]),
    .Y(_5621_)
);

OAI21X1 _16132_ (
    .A(_4786__bF$buf4),
    .B(_5620__bF$buf4),
    .C(_5621_),
    .Y(_4114_)
);

OAI21X1 _16133_ (
    .A(_4794__bF$buf3),
    .B(_4968__bF$buf3),
    .C(\datapath.registers.838[1] [1]),
    .Y(_5622_)
);

OAI21X1 _16134_ (
    .A(_4801__bF$buf2),
    .B(_5620__bF$buf3),
    .C(_5622_),
    .Y(_4125_)
);

OAI21X1 _16135_ (
    .A(_4794__bF$buf2),
    .B(_4968__bF$buf2),
    .C(\datapath.registers.838[1] [2]),
    .Y(_5623_)
);

OAI21X1 _16136_ (
    .A(_4803__bF$buf4),
    .B(_5620__bF$buf2),
    .C(_5623_),
    .Y(_4136_)
);

OAI21X1 _16137_ (
    .A(_4794__bF$buf1),
    .B(_4968__bF$buf1),
    .C(\datapath.registers.838[1] [3]),
    .Y(_5624_)
);

OAI21X1 _16138_ (
    .A(_4805__bF$buf0),
    .B(_5620__bF$buf1),
    .C(_5624_),
    .Y(_4139_)
);

OAI21X1 _16139_ (
    .A(_4794__bF$buf0),
    .B(_4968__bF$buf0),
    .C(\datapath.registers.838[1] [4]),
    .Y(_5625_)
);

OAI21X1 _16140_ (
    .A(_4807__bF$buf3),
    .B(_5620__bF$buf0),
    .C(_5625_),
    .Y(_4140_)
);

OAI21X1 _16141_ (
    .A(_4794__bF$buf7),
    .B(_4968__bF$buf9),
    .C(\datapath.registers.838[1] [5]),
    .Y(_5626_)
);

OAI21X1 _16142_ (
    .A(_4809__bF$buf3),
    .B(_5620__bF$buf4),
    .C(_5626_),
    .Y(_4141_)
);

OAI21X1 _16143_ (
    .A(_4794__bF$buf6),
    .B(_4968__bF$buf8),
    .C(\datapath.registers.838[1] [6]),
    .Y(_5627_)
);

OAI21X1 _16144_ (
    .A(_4811__bF$buf0),
    .B(_5620__bF$buf3),
    .C(_5627_),
    .Y(_4142_)
);

OAI21X1 _16145_ (
    .A(_4794__bF$buf5),
    .B(_4968__bF$buf7),
    .C(\datapath.registers.838[1] [7]),
    .Y(_5628_)
);

OAI21X1 _16146_ (
    .A(_4813__bF$buf2),
    .B(_5620__bF$buf2),
    .C(_5628_),
    .Y(_4143_)
);

OAI21X1 _16147_ (
    .A(_4794__bF$buf4),
    .B(_4968__bF$buf6),
    .C(\datapath.registers.838[1] [8]),
    .Y(_5629_)
);

OAI21X1 _16148_ (
    .A(_4815__bF$buf3),
    .B(_5620__bF$buf1),
    .C(_5629_),
    .Y(_4144_)
);

OAI21X1 _16149_ (
    .A(_4794__bF$buf3),
    .B(_4968__bF$buf5),
    .C(\datapath.registers.838[1] [9]),
    .Y(_5630_)
);

OAI21X1 _16150_ (
    .A(_4817__bF$buf1),
    .B(_5620__bF$buf0),
    .C(_5630_),
    .Y(_4145_)
);

OAI21X1 _16151_ (
    .A(_4794__bF$buf2),
    .B(_4968__bF$buf4),
    .C(\datapath.registers.838[1] [10]),
    .Y(_5631_)
);

OAI21X1 _16152_ (
    .A(_4819__bF$buf4),
    .B(_5620__bF$buf4),
    .C(_5631_),
    .Y(_4115_)
);

OAI21X1 _16153_ (
    .A(_4794__bF$buf1),
    .B(_4968__bF$buf3),
    .C(\datapath.registers.838[1] [11]),
    .Y(_5632_)
);

OAI21X1 _16154_ (
    .A(_4821__bF$buf2),
    .B(_5620__bF$buf3),
    .C(_5632_),
    .Y(_4116_)
);

OAI21X1 _16155_ (
    .A(_4794__bF$buf0),
    .B(_4968__bF$buf2),
    .C(\datapath.registers.838[1] [12]),
    .Y(_5633_)
);

OAI21X1 _16156_ (
    .A(_4823__bF$buf0),
    .B(_5620__bF$buf2),
    .C(_5633_),
    .Y(_4117_)
);

OAI21X1 _16157_ (
    .A(_4794__bF$buf7),
    .B(_4968__bF$buf1),
    .C(\datapath.registers.838[1] [13]),
    .Y(_5634_)
);

OAI21X1 _16158_ (
    .A(_4825__bF$buf2),
    .B(_5620__bF$buf1),
    .C(_5634_),
    .Y(_4118_)
);

OAI21X1 _16159_ (
    .A(_4794__bF$buf6),
    .B(_4968__bF$buf0),
    .C(\datapath.registers.838[1] [14]),
    .Y(_5635_)
);

OAI21X1 _16160_ (
    .A(_4827__bF$buf2),
    .B(_5620__bF$buf0),
    .C(_5635_),
    .Y(_4119_)
);

OAI21X1 _16161_ (
    .A(_4794__bF$buf5),
    .B(_4968__bF$buf9),
    .C(\datapath.registers.838[1] [15]),
    .Y(_5636_)
);

OAI21X1 _16162_ (
    .A(_4829__bF$buf2),
    .B(_5620__bF$buf4),
    .C(_5636_),
    .Y(_4120_)
);

OAI21X1 _16163_ (
    .A(_4794__bF$buf4),
    .B(_4968__bF$buf8),
    .C(\datapath.registers.838[1] [16]),
    .Y(_5637_)
);

OAI21X1 _16164_ (
    .A(_4831__bF$buf2),
    .B(_5620__bF$buf3),
    .C(_5637_),
    .Y(_4121_)
);

OAI21X1 _16165_ (
    .A(_4794__bF$buf3),
    .B(_4968__bF$buf7),
    .C(\datapath.registers.838[1] [17]),
    .Y(_5638_)
);

OAI21X1 _16166_ (
    .A(_4833__bF$buf4),
    .B(_5620__bF$buf2),
    .C(_5638_),
    .Y(_4122_)
);

OAI21X1 _16167_ (
    .A(_4794__bF$buf2),
    .B(_4968__bF$buf6),
    .C(\datapath.registers.838[1] [18]),
    .Y(_5639_)
);

OAI21X1 _16168_ (
    .A(_4835__bF$buf4),
    .B(_5620__bF$buf1),
    .C(_5639_),
    .Y(_4123_)
);

OAI21X1 _16169_ (
    .A(_4794__bF$buf1),
    .B(_4968__bF$buf5),
    .C(\datapath.registers.838[1] [19]),
    .Y(_5640_)
);

OAI21X1 _16170_ (
    .A(_4837__bF$buf0),
    .B(_5620__bF$buf0),
    .C(_5640_),
    .Y(_4124_)
);

OAI21X1 _16171_ (
    .A(_4794__bF$buf0),
    .B(_4968__bF$buf4),
    .C(\datapath.registers.838[1] [20]),
    .Y(_5641_)
);

OAI21X1 _16172_ (
    .A(_4839__bF$buf2),
    .B(_5620__bF$buf4),
    .C(_5641_),
    .Y(_4126_)
);

OAI21X1 _16173_ (
    .A(_4794__bF$buf7),
    .B(_4968__bF$buf3),
    .C(\datapath.registers.838[1] [21]),
    .Y(_5642_)
);

OAI21X1 _16174_ (
    .A(_4841__bF$buf4),
    .B(_5620__bF$buf3),
    .C(_5642_),
    .Y(_4127_)
);

OAI21X1 _16175_ (
    .A(_4794__bF$buf6),
    .B(_4968__bF$buf2),
    .C(\datapath.registers.838[1] [22]),
    .Y(_5643_)
);

OAI21X1 _16176_ (
    .A(_4843__bF$buf3),
    .B(_5620__bF$buf2),
    .C(_5643_),
    .Y(_4128_)
);

OAI21X1 _16177_ (
    .A(_4794__bF$buf5),
    .B(_4968__bF$buf1),
    .C(\datapath.registers.838[1] [23]),
    .Y(_5644_)
);

OAI21X1 _16178_ (
    .A(_4845__bF$buf4),
    .B(_5620__bF$buf1),
    .C(_5644_),
    .Y(_4129_)
);

OAI21X1 _16179_ (
    .A(_4794__bF$buf4),
    .B(_4968__bF$buf0),
    .C(\datapath.registers.838[1] [24]),
    .Y(_5645_)
);

OAI21X1 _16180_ (
    .A(_4847__bF$buf1),
    .B(_5620__bF$buf0),
    .C(_5645_),
    .Y(_4130_)
);

OAI21X1 _16181_ (
    .A(_4794__bF$buf3),
    .B(_4968__bF$buf9),
    .C(\datapath.registers.838[1] [25]),
    .Y(_5646_)
);

OAI21X1 _16182_ (
    .A(_4849__bF$buf4),
    .B(_5620__bF$buf4),
    .C(_5646_),
    .Y(_4131_)
);

OAI21X1 _16183_ (
    .A(_4794__bF$buf2),
    .B(_4968__bF$buf8),
    .C(\datapath.registers.838[1] [26]),
    .Y(_5647_)
);

OAI21X1 _16184_ (
    .A(_4851__bF$buf2),
    .B(_5620__bF$buf3),
    .C(_5647_),
    .Y(_4132_)
);

OAI21X1 _16185_ (
    .A(_4794__bF$buf1),
    .B(_4968__bF$buf7),
    .C(\datapath.registers.838[1] [27]),
    .Y(_5648_)
);

OAI21X1 _16186_ (
    .A(_4853__bF$buf3),
    .B(_5620__bF$buf2),
    .C(_5648_),
    .Y(_4133_)
);

OAI21X1 _16187_ (
    .A(_4794__bF$buf0),
    .B(_4968__bF$buf6),
    .C(\datapath.registers.838[1] [28]),
    .Y(_5649_)
);

OAI21X1 _16188_ (
    .A(_4855__bF$buf2),
    .B(_5620__bF$buf1),
    .C(_5649_),
    .Y(_4134_)
);

OAI21X1 _16189_ (
    .A(_4794__bF$buf7),
    .B(_4968__bF$buf5),
    .C(\datapath.registers.838[1] [29]),
    .Y(_5650_)
);

OAI21X1 _16190_ (
    .A(_4857__bF$buf2),
    .B(_5620__bF$buf0),
    .C(_5650_),
    .Y(_4135_)
);

OAI21X1 _16191_ (
    .A(_4794__bF$buf6),
    .B(_4968__bF$buf4),
    .C(\datapath.registers.838[1] [30]),
    .Y(_5651_)
);

OAI21X1 _16192_ (
    .A(_4859__bF$buf4),
    .B(_5620__bF$buf4),
    .C(_5651_),
    .Y(_4137_)
);

OAI21X1 _16193_ (
    .A(_4794__bF$buf5),
    .B(_4968__bF$buf3),
    .C(\datapath.registers.838[1] [31]),
    .Y(_5652_)
);

OAI21X1 _16194_ (
    .A(_4861__bF$buf2),
    .B(_5620__bF$buf3),
    .C(_5652_),
    .Y(_4138_)
);

NAND2X1 _16195_ (
    .A(_4933_),
    .B(_4798_),
    .Y(_5653_)
);

NAND2X1 _16196_ (
    .A(\datapath.registers.838[22] [0]),
    .B(_5653__bF$buf7),
    .Y(_5654_)
);

OAI21X1 _16197_ (
    .A(_4786__bF$buf3),
    .B(_5653__bF$buf6),
    .C(_5654_),
    .Y(_4210_)
);

NAND2X1 _16198_ (
    .A(\datapath.registers.838[22] [1]),
    .B(_5653__bF$buf5),
    .Y(_5655_)
);

OAI21X1 _16199_ (
    .A(_4801__bF$buf1),
    .B(_5653__bF$buf4),
    .C(_5655_),
    .Y(_4221_)
);

NAND2X1 _16200_ (
    .A(\datapath.registers.838[22] [2]),
    .B(_5653__bF$buf3),
    .Y(_5656_)
);

OAI21X1 _16201_ (
    .A(_4803__bF$buf3),
    .B(_5653__bF$buf2),
    .C(_5656_),
    .Y(_4232_)
);

NAND2X1 _16202_ (
    .A(\datapath.registers.838[22] [3]),
    .B(_5653__bF$buf1),
    .Y(_5657_)
);

OAI21X1 _16203_ (
    .A(_4805__bF$buf4),
    .B(_5653__bF$buf0),
    .C(_5657_),
    .Y(_4235_)
);

NAND2X1 _16204_ (
    .A(\datapath.registers.838[22] [4]),
    .B(_5653__bF$buf7),
    .Y(_5658_)
);

OAI21X1 _16205_ (
    .A(_4807__bF$buf2),
    .B(_5653__bF$buf6),
    .C(_5658_),
    .Y(_4236_)
);

NAND2X1 _16206_ (
    .A(\datapath.registers.838[22] [5]),
    .B(_5653__bF$buf5),
    .Y(_5659_)
);

OAI21X1 _16207_ (
    .A(_4809__bF$buf2),
    .B(_5653__bF$buf4),
    .C(_5659_),
    .Y(_4237_)
);

NAND2X1 _16208_ (
    .A(\datapath.registers.838[22] [6]),
    .B(_5653__bF$buf3),
    .Y(_5660_)
);

OAI21X1 _16209_ (
    .A(_4811__bF$buf4),
    .B(_5653__bF$buf2),
    .C(_5660_),
    .Y(_4238_)
);

NAND2X1 _16210_ (
    .A(\datapath.registers.838[22] [7]),
    .B(_5653__bF$buf1),
    .Y(_5661_)
);

OAI21X1 _16211_ (
    .A(_4813__bF$buf1),
    .B(_5653__bF$buf0),
    .C(_5661_),
    .Y(_4239_)
);

NAND2X1 _16212_ (
    .A(\datapath.registers.838[22] [8]),
    .B(_5653__bF$buf7),
    .Y(_5662_)
);

OAI21X1 _16213_ (
    .A(_4815__bF$buf2),
    .B(_5653__bF$buf6),
    .C(_5662_),
    .Y(_4240_)
);

NAND2X1 _16214_ (
    .A(\datapath.registers.838[22] [9]),
    .B(_5653__bF$buf5),
    .Y(_5663_)
);

OAI21X1 _16215_ (
    .A(_4817__bF$buf0),
    .B(_5653__bF$buf4),
    .C(_5663_),
    .Y(_4241_)
);

NAND2X1 _16216_ (
    .A(\datapath.registers.838[22] [10]),
    .B(_5653__bF$buf3),
    .Y(_5664_)
);

OAI21X1 _16217_ (
    .A(_4819__bF$buf3),
    .B(_5653__bF$buf2),
    .C(_5664_),
    .Y(_4211_)
);

NAND2X1 _16218_ (
    .A(\datapath.registers.838[22] [11]),
    .B(_5653__bF$buf1),
    .Y(_5665_)
);

OAI21X1 _16219_ (
    .A(_4821__bF$buf1),
    .B(_5653__bF$buf0),
    .C(_5665_),
    .Y(_4212_)
);

NAND2X1 _16220_ (
    .A(\datapath.registers.838[22] [12]),
    .B(_5653__bF$buf7),
    .Y(_5666_)
);

OAI21X1 _16221_ (
    .A(_4823__bF$buf4),
    .B(_5653__bF$buf6),
    .C(_5666_),
    .Y(_4213_)
);

NAND2X1 _16222_ (
    .A(\datapath.registers.838[22] [13]),
    .B(_5653__bF$buf5),
    .Y(_5667_)
);

OAI21X1 _16223_ (
    .A(_4825__bF$buf1),
    .B(_5653__bF$buf4),
    .C(_5667_),
    .Y(_4214_)
);

NAND2X1 _16224_ (
    .A(\datapath.registers.838[22] [14]),
    .B(_5653__bF$buf3),
    .Y(_5668_)
);

OAI21X1 _16225_ (
    .A(_4827__bF$buf1),
    .B(_5653__bF$buf2),
    .C(_5668_),
    .Y(_4215_)
);

NAND2X1 _16226_ (
    .A(\datapath.registers.838[22] [15]),
    .B(_5653__bF$buf1),
    .Y(_5669_)
);

OAI21X1 _16227_ (
    .A(_4829__bF$buf1),
    .B(_5653__bF$buf0),
    .C(_5669_),
    .Y(_4216_)
);

NAND2X1 _16228_ (
    .A(\datapath.registers.838[22] [16]),
    .B(_5653__bF$buf7),
    .Y(_5670_)
);

OAI21X1 _16229_ (
    .A(_4831__bF$buf1),
    .B(_5653__bF$buf6),
    .C(_5670_),
    .Y(_4217_)
);

NAND2X1 _16230_ (
    .A(\datapath.registers.838[22] [17]),
    .B(_5653__bF$buf5),
    .Y(_5671_)
);

OAI21X1 _16231_ (
    .A(_4833__bF$buf3),
    .B(_5653__bF$buf4),
    .C(_5671_),
    .Y(_4218_)
);

NAND2X1 _16232_ (
    .A(\datapath.registers.838[22] [18]),
    .B(_5653__bF$buf3),
    .Y(_5672_)
);

OAI21X1 _16233_ (
    .A(_4835__bF$buf3),
    .B(_5653__bF$buf2),
    .C(_5672_),
    .Y(_4219_)
);

NAND2X1 _16234_ (
    .A(\datapath.registers.838[22] [19]),
    .B(_5653__bF$buf1),
    .Y(_5673_)
);

OAI21X1 _16235_ (
    .A(_4837__bF$buf4),
    .B(_5653__bF$buf0),
    .C(_5673_),
    .Y(_4220_)
);

NAND2X1 _16236_ (
    .A(\datapath.registers.838[22] [20]),
    .B(_5653__bF$buf7),
    .Y(_5674_)
);

OAI21X1 _16237_ (
    .A(_4839__bF$buf1),
    .B(_5653__bF$buf6),
    .C(_5674_),
    .Y(_4222_)
);

NAND2X1 _16238_ (
    .A(\datapath.registers.838[22] [21]),
    .B(_5653__bF$buf5),
    .Y(_5675_)
);

OAI21X1 _16239_ (
    .A(_4841__bF$buf3),
    .B(_5653__bF$buf4),
    .C(_5675_),
    .Y(_4223_)
);

NAND2X1 _16240_ (
    .A(\datapath.registers.838[22] [22]),
    .B(_5653__bF$buf3),
    .Y(_5676_)
);

OAI21X1 _16241_ (
    .A(_4843__bF$buf2),
    .B(_5653__bF$buf2),
    .C(_5676_),
    .Y(_4224_)
);

NAND2X1 _16242_ (
    .A(\datapath.registers.838[22] [23]),
    .B(_5653__bF$buf1),
    .Y(_5677_)
);

OAI21X1 _16243_ (
    .A(_4845__bF$buf3),
    .B(_5653__bF$buf0),
    .C(_5677_),
    .Y(_4225_)
);

NAND2X1 _16244_ (
    .A(\datapath.registers.838[22] [24]),
    .B(_5653__bF$buf7),
    .Y(_5678_)
);

OAI21X1 _16245_ (
    .A(_4847__bF$buf0),
    .B(_5653__bF$buf6),
    .C(_5678_),
    .Y(_4226_)
);

NAND2X1 _16246_ (
    .A(\datapath.registers.838[22] [25]),
    .B(_5653__bF$buf5),
    .Y(_5679_)
);

OAI21X1 _16247_ (
    .A(_4849__bF$buf3),
    .B(_5653__bF$buf4),
    .C(_5679_),
    .Y(_4227_)
);

NAND2X1 _16248_ (
    .A(\datapath.registers.838[22] [26]),
    .B(_5653__bF$buf3),
    .Y(_5680_)
);

OAI21X1 _16249_ (
    .A(_4851__bF$buf1),
    .B(_5653__bF$buf2),
    .C(_5680_),
    .Y(_4228_)
);

NAND2X1 _16250_ (
    .A(\datapath.registers.838[22] [27]),
    .B(_5653__bF$buf1),
    .Y(_5681_)
);

OAI21X1 _16251_ (
    .A(_4853__bF$buf2),
    .B(_5653__bF$buf0),
    .C(_5681_),
    .Y(_4229_)
);

NAND2X1 _16252_ (
    .A(\datapath.registers.838[22] [28]),
    .B(_5653__bF$buf7),
    .Y(_5682_)
);

OAI21X1 _16253_ (
    .A(_4855__bF$buf1),
    .B(_5653__bF$buf6),
    .C(_5682_),
    .Y(_4230_)
);

NAND2X1 _16254_ (
    .A(\datapath.registers.838[22] [29]),
    .B(_5653__bF$buf5),
    .Y(_5683_)
);

OAI21X1 _16255_ (
    .A(_4857__bF$buf1),
    .B(_5653__bF$buf4),
    .C(_5683_),
    .Y(_4231_)
);

NAND2X1 _16256_ (
    .A(\datapath.registers.838[22] [30]),
    .B(_5653__bF$buf3),
    .Y(_5684_)
);

OAI21X1 _16257_ (
    .A(_4859__bF$buf3),
    .B(_5653__bF$buf2),
    .C(_5684_),
    .Y(_4233_)
);

NAND2X1 _16258_ (
    .A(\datapath.registers.838[22] [31]),
    .B(_5653__bF$buf1),
    .Y(_5685_)
);

OAI21X1 _16259_ (
    .A(_4861__bF$buf1),
    .B(_5653__bF$buf0),
    .C(_5685_),
    .Y(_4234_)
);

INVX1 _16260_ (
    .A(_4899__bF$buf6),
    .Y(_5686_)
);

OR2X2 _16261_ (
    .A(_5475_),
    .B(_4791_),
    .Y(_5687_)
);

INVX1 _16262_ (
    .A(_5687__bF$buf8),
    .Y(_5688_)
);

NAND2X1 _16263_ (
    .A(_5688_),
    .B(_5686_),
    .Y(_5689_)
);

OAI21X1 _16264_ (
    .A(_5687__bF$buf7),
    .B(_4899__bF$buf5),
    .C(\datapath.registers.838[31] [0]),
    .Y(_5690_)
);

OAI21X1 _16265_ (
    .A(_4786__bF$buf2),
    .B(_5689__bF$buf4),
    .C(_5690_),
    .Y(_4530_)
);

OAI21X1 _16266_ (
    .A(_5687__bF$buf6),
    .B(_4899__bF$buf4),
    .C(\datapath.registers.838[31] [1]),
    .Y(_5691_)
);

OAI21X1 _16267_ (
    .A(_4801__bF$buf0),
    .B(_5689__bF$buf3),
    .C(_5691_),
    .Y(_4541_)
);

OAI21X1 _16268_ (
    .A(_5687__bF$buf5),
    .B(_4899__bF$buf3),
    .C(\datapath.registers.838[31] [2]),
    .Y(_5692_)
);

OAI21X1 _16269_ (
    .A(_4803__bF$buf2),
    .B(_5689__bF$buf2),
    .C(_5692_),
    .Y(_4552_)
);

OAI21X1 _16270_ (
    .A(_5687__bF$buf4),
    .B(_4899__bF$buf2),
    .C(\datapath.registers.838[31] [3]),
    .Y(_5693_)
);

OAI21X1 _16271_ (
    .A(_4805__bF$buf3),
    .B(_5689__bF$buf1),
    .C(_5693_),
    .Y(_4555_)
);

OAI21X1 _16272_ (
    .A(_5687__bF$buf3),
    .B(_4899__bF$buf1),
    .C(\datapath.registers.838[31] [4]),
    .Y(_5694_)
);

OAI21X1 _16273_ (
    .A(_4807__bF$buf1),
    .B(_5689__bF$buf0),
    .C(_5694_),
    .Y(_4556_)
);

OAI21X1 _16274_ (
    .A(_5687__bF$buf2),
    .B(_4899__bF$buf0),
    .C(\datapath.registers.838[31] [5]),
    .Y(_5695_)
);

OAI21X1 _16275_ (
    .A(_4809__bF$buf1),
    .B(_5689__bF$buf4),
    .C(_5695_),
    .Y(_4557_)
);

OAI21X1 _16276_ (
    .A(_5687__bF$buf1),
    .B(_4899__bF$buf13),
    .C(\datapath.registers.838[31] [6]),
    .Y(_5696_)
);

OAI21X1 _16277_ (
    .A(_4811__bF$buf3),
    .B(_5689__bF$buf3),
    .C(_5696_),
    .Y(_4558_)
);

OAI21X1 _16278_ (
    .A(_5687__bF$buf0),
    .B(_4899__bF$buf12),
    .C(\datapath.registers.838[31] [7]),
    .Y(_5697_)
);

OAI21X1 _16279_ (
    .A(_4813__bF$buf0),
    .B(_5689__bF$buf2),
    .C(_5697_),
    .Y(_4559_)
);

OAI21X1 _16280_ (
    .A(_5687__bF$buf8),
    .B(_4899__bF$buf11),
    .C(\datapath.registers.838[31] [8]),
    .Y(_5698_)
);

OAI21X1 _16281_ (
    .A(_4815__bF$buf1),
    .B(_5689__bF$buf1),
    .C(_5698_),
    .Y(_4560_)
);

OAI21X1 _16282_ (
    .A(_5687__bF$buf7),
    .B(_4899__bF$buf10),
    .C(\datapath.registers.838[31] [9]),
    .Y(_5699_)
);

OAI21X1 _16283_ (
    .A(_4817__bF$buf4),
    .B(_5689__bF$buf0),
    .C(_5699_),
    .Y(_4561_)
);

OAI21X1 _16284_ (
    .A(_5687__bF$buf6),
    .B(_4899__bF$buf9),
    .C(\datapath.registers.838[31] [10]),
    .Y(_5700_)
);

OAI21X1 _16285_ (
    .A(_4819__bF$buf2),
    .B(_5689__bF$buf4),
    .C(_5700_),
    .Y(_4531_)
);

OAI21X1 _16286_ (
    .A(_5687__bF$buf5),
    .B(_4899__bF$buf8),
    .C(\datapath.registers.838[31] [11]),
    .Y(_5701_)
);

OAI21X1 _16287_ (
    .A(_4821__bF$buf0),
    .B(_5689__bF$buf3),
    .C(_5701_),
    .Y(_4532_)
);

OAI21X1 _16288_ (
    .A(_5687__bF$buf4),
    .B(_4899__bF$buf7),
    .C(\datapath.registers.838[31] [12]),
    .Y(_5702_)
);

OAI21X1 _16289_ (
    .A(_4823__bF$buf3),
    .B(_5689__bF$buf2),
    .C(_5702_),
    .Y(_4533_)
);

OAI21X1 _16290_ (
    .A(_5687__bF$buf3),
    .B(_4899__bF$buf6),
    .C(\datapath.registers.838[31] [13]),
    .Y(_5703_)
);

OAI21X1 _16291_ (
    .A(_4825__bF$buf0),
    .B(_5689__bF$buf1),
    .C(_5703_),
    .Y(_4534_)
);

OAI21X1 _16292_ (
    .A(_5687__bF$buf2),
    .B(_4899__bF$buf5),
    .C(\datapath.registers.838[31] [14]),
    .Y(_5704_)
);

OAI21X1 _16293_ (
    .A(_4827__bF$buf0),
    .B(_5689__bF$buf0),
    .C(_5704_),
    .Y(_4535_)
);

OAI21X1 _16294_ (
    .A(_5687__bF$buf1),
    .B(_4899__bF$buf4),
    .C(\datapath.registers.838[31] [15]),
    .Y(_5705_)
);

OAI21X1 _16295_ (
    .A(_4829__bF$buf0),
    .B(_5689__bF$buf4),
    .C(_5705_),
    .Y(_4536_)
);

OAI21X1 _16296_ (
    .A(_5687__bF$buf0),
    .B(_4899__bF$buf3),
    .C(\datapath.registers.838[31] [16]),
    .Y(_5706_)
);

OAI21X1 _16297_ (
    .A(_4831__bF$buf0),
    .B(_5689__bF$buf3),
    .C(_5706_),
    .Y(_4537_)
);

OAI21X1 _16298_ (
    .A(_5687__bF$buf8),
    .B(_4899__bF$buf2),
    .C(\datapath.registers.838[31] [17]),
    .Y(_5707_)
);

OAI21X1 _16299_ (
    .A(_4833__bF$buf2),
    .B(_5689__bF$buf2),
    .C(_5707_),
    .Y(_4538_)
);

OAI21X1 _16300_ (
    .A(_5687__bF$buf7),
    .B(_4899__bF$buf1),
    .C(\datapath.registers.838[31] [18]),
    .Y(_5708_)
);

OAI21X1 _16301_ (
    .A(_4835__bF$buf2),
    .B(_5689__bF$buf1),
    .C(_5708_),
    .Y(_4539_)
);

OAI21X1 _16302_ (
    .A(_5687__bF$buf6),
    .B(_4899__bF$buf0),
    .C(\datapath.registers.838[31] [19]),
    .Y(_5709_)
);

OAI21X1 _16303_ (
    .A(_4837__bF$buf3),
    .B(_5689__bF$buf0),
    .C(_5709_),
    .Y(_4540_)
);

OAI21X1 _16304_ (
    .A(_5687__bF$buf5),
    .B(_4899__bF$buf13),
    .C(\datapath.registers.838[31] [20]),
    .Y(_5710_)
);

OAI21X1 _16305_ (
    .A(_4839__bF$buf0),
    .B(_5689__bF$buf4),
    .C(_5710_),
    .Y(_4542_)
);

OAI21X1 _16306_ (
    .A(_5687__bF$buf4),
    .B(_4899__bF$buf12),
    .C(\datapath.registers.838[31] [21]),
    .Y(_5711_)
);

OAI21X1 _16307_ (
    .A(_4841__bF$buf2),
    .B(_5689__bF$buf3),
    .C(_5711_),
    .Y(_4543_)
);

OAI21X1 _16308_ (
    .A(_5687__bF$buf3),
    .B(_4899__bF$buf11),
    .C(\datapath.registers.838[31] [22]),
    .Y(_5712_)
);

OAI21X1 _16309_ (
    .A(_4843__bF$buf1),
    .B(_5689__bF$buf2),
    .C(_5712_),
    .Y(_4544_)
);

OAI21X1 _16310_ (
    .A(_5687__bF$buf2),
    .B(_4899__bF$buf10),
    .C(\datapath.registers.838[31] [23]),
    .Y(_5713_)
);

OAI21X1 _16311_ (
    .A(_4845__bF$buf2),
    .B(_5689__bF$buf1),
    .C(_5713_),
    .Y(_4545_)
);

OAI21X1 _16312_ (
    .A(_5687__bF$buf1),
    .B(_4899__bF$buf9),
    .C(\datapath.registers.838[31] [24]),
    .Y(_5714_)
);

OAI21X1 _16313_ (
    .A(_4847__bF$buf4),
    .B(_5689__bF$buf0),
    .C(_5714_),
    .Y(_4546_)
);

OAI21X1 _16314_ (
    .A(_5687__bF$buf0),
    .B(_4899__bF$buf8),
    .C(\datapath.registers.838[31] [25]),
    .Y(_5715_)
);

OAI21X1 _16315_ (
    .A(_4849__bF$buf2),
    .B(_5689__bF$buf4),
    .C(_5715_),
    .Y(_4547_)
);

OAI21X1 _16316_ (
    .A(_5687__bF$buf8),
    .B(_4899__bF$buf7),
    .C(\datapath.registers.838[31] [26]),
    .Y(_5716_)
);

OAI21X1 _16317_ (
    .A(_4851__bF$buf0),
    .B(_5689__bF$buf3),
    .C(_5716_),
    .Y(_4548_)
);

OAI21X1 _16318_ (
    .A(_5687__bF$buf7),
    .B(_4899__bF$buf6),
    .C(\datapath.registers.838[31] [27]),
    .Y(_5717_)
);

OAI21X1 _16319_ (
    .A(_4853__bF$buf1),
    .B(_5689__bF$buf2),
    .C(_5717_),
    .Y(_4549_)
);

OAI21X1 _16320_ (
    .A(_5687__bF$buf6),
    .B(_4899__bF$buf5),
    .C(\datapath.registers.838[31] [28]),
    .Y(_5718_)
);

OAI21X1 _16321_ (
    .A(_4855__bF$buf0),
    .B(_5689__bF$buf1),
    .C(_5718_),
    .Y(_4550_)
);

OAI21X1 _16322_ (
    .A(_5687__bF$buf5),
    .B(_4899__bF$buf4),
    .C(\datapath.registers.838[31] [29]),
    .Y(_5719_)
);

OAI21X1 _16323_ (
    .A(_4857__bF$buf0),
    .B(_5689__bF$buf0),
    .C(_5719_),
    .Y(_4551_)
);

OAI21X1 _16324_ (
    .A(_5687__bF$buf4),
    .B(_4899__bF$buf3),
    .C(\datapath.registers.838[31] [30]),
    .Y(_5720_)
);

OAI21X1 _16325_ (
    .A(_4859__bF$buf2),
    .B(_5689__bF$buf4),
    .C(_5720_),
    .Y(_4553_)
);

OAI21X1 _16326_ (
    .A(_5687__bF$buf3),
    .B(_4899__bF$buf2),
    .C(\datapath.registers.838[31] [31]),
    .Y(_5721_)
);

OAI21X1 _16327_ (
    .A(_4861__bF$buf0),
    .B(_5689__bF$buf3),
    .C(_5721_),
    .Y(_4554_)
);

NAND2X1 _16328_ (
    .A(_5688_),
    .B(_5585_),
    .Y(_5722_)
);

OAI21X1 _16329_ (
    .A(_5687__bF$buf2),
    .B(_4934__bF$buf2),
    .C(\datapath.registers.838[30] [0]),
    .Y(_5723_)
);

OAI21X1 _16330_ (
    .A(_4786__bF$buf1),
    .B(_5722__bF$buf4),
    .C(_5723_),
    .Y(_4498_)
);

OAI21X1 _16331_ (
    .A(_5687__bF$buf1),
    .B(_4934__bF$buf1),
    .C(\datapath.registers.838[30] [1]),
    .Y(_5724_)
);

OAI21X1 _16332_ (
    .A(_4801__bF$buf4),
    .B(_5722__bF$buf3),
    .C(_5724_),
    .Y(_4509_)
);

OAI21X1 _16333_ (
    .A(_5687__bF$buf0),
    .B(_4934__bF$buf0),
    .C(\datapath.registers.838[30] [2]),
    .Y(_5725_)
);

OAI21X1 _16334_ (
    .A(_4803__bF$buf1),
    .B(_5722__bF$buf2),
    .C(_5725_),
    .Y(_4520_)
);

OAI21X1 _16335_ (
    .A(_5687__bF$buf8),
    .B(_4934__bF$buf9),
    .C(\datapath.registers.838[30] [3]),
    .Y(_5726_)
);

OAI21X1 _16336_ (
    .A(_4805__bF$buf2),
    .B(_5722__bF$buf1),
    .C(_5726_),
    .Y(_4523_)
);

OAI21X1 _16337_ (
    .A(_5687__bF$buf7),
    .B(_4934__bF$buf8),
    .C(\datapath.registers.838[30] [4]),
    .Y(_5727_)
);

OAI21X1 _16338_ (
    .A(_4807__bF$buf0),
    .B(_5722__bF$buf0),
    .C(_5727_),
    .Y(_4524_)
);

OAI21X1 _16339_ (
    .A(_5687__bF$buf6),
    .B(_4934__bF$buf7),
    .C(\datapath.registers.838[30] [5]),
    .Y(_5728_)
);

OAI21X1 _16340_ (
    .A(_4809__bF$buf0),
    .B(_5722__bF$buf4),
    .C(_5728_),
    .Y(_4525_)
);

OAI21X1 _16341_ (
    .A(_5687__bF$buf5),
    .B(_4934__bF$buf6),
    .C(\datapath.registers.838[30] [6]),
    .Y(_5729_)
);

OAI21X1 _16342_ (
    .A(_4811__bF$buf2),
    .B(_5722__bF$buf3),
    .C(_5729_),
    .Y(_4526_)
);

OAI21X1 _16343_ (
    .A(_5687__bF$buf4),
    .B(_4934__bF$buf5),
    .C(\datapath.registers.838[30] [7]),
    .Y(_5730_)
);

OAI21X1 _16344_ (
    .A(_4813__bF$buf4),
    .B(_5722__bF$buf2),
    .C(_5730_),
    .Y(_4527_)
);

OAI21X1 _16345_ (
    .A(_5687__bF$buf3),
    .B(_4934__bF$buf4),
    .C(\datapath.registers.838[30] [8]),
    .Y(_5731_)
);

OAI21X1 _16346_ (
    .A(_4815__bF$buf0),
    .B(_5722__bF$buf1),
    .C(_5731_),
    .Y(_4528_)
);

OAI21X1 _16347_ (
    .A(_5687__bF$buf2),
    .B(_4934__bF$buf3),
    .C(\datapath.registers.838[30] [9]),
    .Y(_5732_)
);

OAI21X1 _16348_ (
    .A(_4817__bF$buf3),
    .B(_5722__bF$buf0),
    .C(_5732_),
    .Y(_4529_)
);

OAI21X1 _16349_ (
    .A(_5687__bF$buf1),
    .B(_4934__bF$buf2),
    .C(\datapath.registers.838[30] [10]),
    .Y(_5733_)
);

OAI21X1 _16350_ (
    .A(_4819__bF$buf1),
    .B(_5722__bF$buf4),
    .C(_5733_),
    .Y(_4499_)
);

OAI21X1 _16351_ (
    .A(_5687__bF$buf0),
    .B(_4934__bF$buf1),
    .C(\datapath.registers.838[30] [11]),
    .Y(_5734_)
);

OAI21X1 _16352_ (
    .A(_4821__bF$buf4),
    .B(_5722__bF$buf3),
    .C(_5734_),
    .Y(_4500_)
);

OAI21X1 _16353_ (
    .A(_5687__bF$buf8),
    .B(_4934__bF$buf0),
    .C(\datapath.registers.838[30] [12]),
    .Y(_5735_)
);

OAI21X1 _16354_ (
    .A(_4823__bF$buf2),
    .B(_5722__bF$buf2),
    .C(_5735_),
    .Y(_4501_)
);

OAI21X1 _16355_ (
    .A(_5687__bF$buf7),
    .B(_4934__bF$buf9),
    .C(\datapath.registers.838[30] [13]),
    .Y(_5736_)
);

OAI21X1 _16356_ (
    .A(_4825__bF$buf4),
    .B(_5722__bF$buf1),
    .C(_5736_),
    .Y(_4502_)
);

OAI21X1 _16357_ (
    .A(_5687__bF$buf6),
    .B(_4934__bF$buf8),
    .C(\datapath.registers.838[30] [14]),
    .Y(_5737_)
);

OAI21X1 _16358_ (
    .A(_4827__bF$buf4),
    .B(_5722__bF$buf0),
    .C(_5737_),
    .Y(_4503_)
);

OAI21X1 _16359_ (
    .A(_5687__bF$buf5),
    .B(_4934__bF$buf7),
    .C(\datapath.registers.838[30] [15]),
    .Y(_5738_)
);

OAI21X1 _16360_ (
    .A(_4829__bF$buf4),
    .B(_5722__bF$buf4),
    .C(_5738_),
    .Y(_4504_)
);

OAI21X1 _16361_ (
    .A(_5687__bF$buf4),
    .B(_4934__bF$buf6),
    .C(\datapath.registers.838[30] [16]),
    .Y(_5739_)
);

OAI21X1 _16362_ (
    .A(_4831__bF$buf4),
    .B(_5722__bF$buf3),
    .C(_5739_),
    .Y(_4505_)
);

OAI21X1 _16363_ (
    .A(_5687__bF$buf3),
    .B(_4934__bF$buf5),
    .C(\datapath.registers.838[30] [17]),
    .Y(_5740_)
);

OAI21X1 _16364_ (
    .A(_4833__bF$buf1),
    .B(_5722__bF$buf2),
    .C(_5740_),
    .Y(_4506_)
);

OAI21X1 _16365_ (
    .A(_5687__bF$buf2),
    .B(_4934__bF$buf4),
    .C(\datapath.registers.838[30] [18]),
    .Y(_5741_)
);

OAI21X1 _16366_ (
    .A(_4835__bF$buf1),
    .B(_5722__bF$buf1),
    .C(_5741_),
    .Y(_4507_)
);

OAI21X1 _16367_ (
    .A(_5687__bF$buf1),
    .B(_4934__bF$buf3),
    .C(\datapath.registers.838[30] [19]),
    .Y(_5742_)
);

OAI21X1 _16368_ (
    .A(_4837__bF$buf2),
    .B(_5722__bF$buf0),
    .C(_5742_),
    .Y(_4508_)
);

OAI21X1 _16369_ (
    .A(_5687__bF$buf0),
    .B(_4934__bF$buf2),
    .C(\datapath.registers.838[30] [20]),
    .Y(_5743_)
);

OAI21X1 _16370_ (
    .A(_4839__bF$buf4),
    .B(_5722__bF$buf4),
    .C(_5743_),
    .Y(_4510_)
);

OAI21X1 _16371_ (
    .A(_5687__bF$buf8),
    .B(_4934__bF$buf1),
    .C(\datapath.registers.838[30] [21]),
    .Y(_5744_)
);

OAI21X1 _16372_ (
    .A(_4841__bF$buf1),
    .B(_5722__bF$buf3),
    .C(_5744_),
    .Y(_4511_)
);

OAI21X1 _16373_ (
    .A(_5687__bF$buf7),
    .B(_4934__bF$buf0),
    .C(\datapath.registers.838[30] [22]),
    .Y(_5745_)
);

OAI21X1 _16374_ (
    .A(_4843__bF$buf0),
    .B(_5722__bF$buf2),
    .C(_5745_),
    .Y(_4512_)
);

OAI21X1 _16375_ (
    .A(_5687__bF$buf6),
    .B(_4934__bF$buf9),
    .C(\datapath.registers.838[30] [23]),
    .Y(_5746_)
);

OAI21X1 _16376_ (
    .A(_4845__bF$buf1),
    .B(_5722__bF$buf1),
    .C(_5746_),
    .Y(_4513_)
);

OAI21X1 _16377_ (
    .A(_5687__bF$buf5),
    .B(_4934__bF$buf8),
    .C(\datapath.registers.838[30] [24]),
    .Y(_5747_)
);

OAI21X1 _16378_ (
    .A(_4847__bF$buf3),
    .B(_5722__bF$buf0),
    .C(_5747_),
    .Y(_4514_)
);

OAI21X1 _16379_ (
    .A(_5687__bF$buf4),
    .B(_4934__bF$buf7),
    .C(\datapath.registers.838[30] [25]),
    .Y(_5748_)
);

OAI21X1 _16380_ (
    .A(_4849__bF$buf1),
    .B(_5722__bF$buf4),
    .C(_5748_),
    .Y(_4515_)
);

OAI21X1 _16381_ (
    .A(_5687__bF$buf3),
    .B(_4934__bF$buf6),
    .C(\datapath.registers.838[30] [26]),
    .Y(_5749_)
);

OAI21X1 _16382_ (
    .A(_4851__bF$buf4),
    .B(_5722__bF$buf3),
    .C(_5749_),
    .Y(_4516_)
);

OAI21X1 _16383_ (
    .A(_5687__bF$buf2),
    .B(_4934__bF$buf5),
    .C(\datapath.registers.838[30] [27]),
    .Y(_5750_)
);

OAI21X1 _16384_ (
    .A(_4853__bF$buf0),
    .B(_5722__bF$buf2),
    .C(_5750_),
    .Y(_4517_)
);

OAI21X1 _16385_ (
    .A(_5687__bF$buf1),
    .B(_4934__bF$buf4),
    .C(\datapath.registers.838[30] [28]),
    .Y(_5751_)
);

OAI21X1 _16386_ (
    .A(_4855__bF$buf4),
    .B(_5722__bF$buf1),
    .C(_5751_),
    .Y(_4518_)
);

OAI21X1 _16387_ (
    .A(_5687__bF$buf0),
    .B(_4934__bF$buf3),
    .C(\datapath.registers.838[30] [29]),
    .Y(_5752_)
);

OAI21X1 _16388_ (
    .A(_4857__bF$buf4),
    .B(_5722__bF$buf0),
    .C(_5752_),
    .Y(_4519_)
);

OAI21X1 _16389_ (
    .A(_5687__bF$buf8),
    .B(_4934__bF$buf2),
    .C(\datapath.registers.838[30] [30]),
    .Y(_5753_)
);

OAI21X1 _16390_ (
    .A(_4859__bF$buf1),
    .B(_5722__bF$buf4),
    .C(_5753_),
    .Y(_4521_)
);

OAI21X1 _16391_ (
    .A(_5687__bF$buf7),
    .B(_4934__bF$buf1),
    .C(\datapath.registers.838[30] [31]),
    .Y(_5754_)
);

OAI21X1 _16392_ (
    .A(_4861__bF$buf4),
    .B(_5722__bF$buf3),
    .C(_5754_),
    .Y(_4522_)
);

NOR2X1 _16393_ (
    .A(\datapath.idinstr_19_bF$buf2 ),
    .B(\datapath.idinstr_15_bF$buf51 ),
    .Y(_5755_)
);

INVX8 _16394_ (
    .A(\datapath.idinstr_16_bF$buf48 ),
    .Y(_5756_)
);

INVX8 _16395_ (
    .A(\datapath.idinstr_17_bF$buf12 ),
    .Y(_5757_)
);

NAND2X1 _16396_ (
    .A(_5756__bF$buf9),
    .B(_5757__bF$buf10),
    .Y(_5758_)
);

NOR2X1 _16397_ (
    .A(\datapath.idinstr_18_bF$buf3 ),
    .B(_5758_),
    .Y(_5759_)
);

INVX8 _16398_ (
    .A(\datapath.idinstr_18_bF$buf2 ),
    .Y(_5760_)
);

NAND2X1 _16399_ (
    .A(\datapath.idinstr_15_bF$buf50 ),
    .B(\datapath.registers.838[27] [0]),
    .Y(_5761_)
);

INVX8 _16400_ (
    .A(\datapath.idinstr_15_bF$buf49 ),
    .Y(_5762_)
);

NAND2X1 _16401_ (
    .A(\datapath.registers.838[26] [0]),
    .B(_5762__bF$buf47),
    .Y(_5763_)
);

NAND3X1 _16402_ (
    .A(\datapath.idinstr_16_bF$buf47 ),
    .B(_5761_),
    .C(_5763_),
    .Y(_5764_)
);

NAND2X1 _16403_ (
    .A(\datapath.idinstr_15_bF$buf48 ),
    .B(\datapath.registers.838[25] [0]),
    .Y(_5765_)
);

AOI21X1 _16404_ (
    .A(_5762__bF$buf46),
    .B(\datapath.registers.838[24] [0]),
    .C(\datapath.idinstr_16_bF$buf46 ),
    .Y(_5766_)
);

NAND2X1 _16405_ (
    .A(_5765_),
    .B(_5766_),
    .Y(_5767_)
);

NAND3X1 _16406_ (
    .A(_5757__bF$buf9),
    .B(_5764_),
    .C(_5767_),
    .Y(_5768_)
);

NAND2X1 _16407_ (
    .A(\datapath.registers.838[31] [0]),
    .B(\datapath.idinstr_15_bF$buf47 ),
    .Y(_5769_)
);

AOI21X1 _16408_ (
    .A(_5762__bF$buf45),
    .B(\datapath.registers.838[30] [0]),
    .C(_5756__bF$buf8),
    .Y(_5770_)
);

NAND2X1 _16409_ (
    .A(_5769_),
    .B(_5770_),
    .Y(_5771_)
);

INVX1 _16410_ (
    .A(\datapath.registers.838[28] [0]),
    .Y(_5772_)
);

AOI21X1 _16411_ (
    .A(\datapath.idinstr_15_bF$buf46 ),
    .B(\datapath.registers.838[29] [0]),
    .C(\datapath.idinstr_16_bF$buf45 ),
    .Y(_5773_)
);

OAI21X1 _16412_ (
    .A(\datapath.idinstr_15_bF$buf45 ),
    .B(_5772_),
    .C(_5773_),
    .Y(_5774_)
);

NAND3X1 _16413_ (
    .A(\datapath.idinstr_17_bF$buf11 ),
    .B(_5774_),
    .C(_5771_),
    .Y(_5775_)
);

AOI21X1 _16414_ (
    .A(_5768_),
    .B(_5775_),
    .C(_5760__bF$buf7),
    .Y(_5776_)
);

MUX2X1 _16415_ (
    .A(\datapath.registers.838[18] [0]),
    .B(\datapath.registers.838[16] [0]),
    .S(\datapath.idinstr_16_bF$buf44 ),
    .Y(_5777_)
);

NAND2X1 _16416_ (
    .A(_5762__bF$buf44),
    .B(_5777_),
    .Y(_5778_)
);

MUX2X1 _16417_ (
    .A(\datapath.registers.838[19] [0]),
    .B(\datapath.registers.838[17] [0]),
    .S(\datapath.idinstr_16_bF$buf43 ),
    .Y(_5779_)
);

NAND2X1 _16418_ (
    .A(\datapath.idinstr_15_bF$buf44 ),
    .B(_5779_),
    .Y(_5780_)
);

NAND3X1 _16419_ (
    .A(_5757__bF$buf8),
    .B(_5778_),
    .C(_5780_),
    .Y(_5781_)
);

MUX2X1 _16420_ (
    .A(\datapath.registers.838[22] [0]),
    .B(\datapath.registers.838[20] [0]),
    .S(\datapath.idinstr_16_bF$buf42 ),
    .Y(_5782_)
);

NAND2X1 _16421_ (
    .A(_5762__bF$buf43),
    .B(_5782_),
    .Y(_5783_)
);

MUX2X1 _16422_ (
    .A(\datapath.registers.838[23] [0]),
    .B(\datapath.registers.838[21] [0]),
    .S(\datapath.idinstr_16_bF$buf41 ),
    .Y(_5784_)
);

NAND2X1 _16423_ (
    .A(\datapath.idinstr_15_bF$buf43 ),
    .B(_5784_),
    .Y(_5785_)
);

NAND3X1 _16424_ (
    .A(\datapath.idinstr_17_bF$buf10 ),
    .B(_5783_),
    .C(_5785_),
    .Y(_5786_)
);

AOI21X1 _16425_ (
    .A(_5781_),
    .B(_5786_),
    .C(\datapath.idinstr_18_bF$buf1 ),
    .Y(_5787_)
);

OAI21X1 _16426_ (
    .A(_5787_),
    .B(_5776_),
    .C(\datapath.idinstr_19_bF$buf1 ),
    .Y(_5788_)
);

INVX8 _16427_ (
    .A(\datapath.idinstr_19_bF$buf0 ),
    .Y(_5789_)
);

AOI21X1 _16428_ (
    .A(\datapath.registers.838[13] [0]),
    .B(\datapath.idinstr_17_bF$buf9 ),
    .C(_5762__bF$buf42),
    .Y(_5790_)
);

OAI21X1 _16429_ (
    .A(_5263_),
    .B(\datapath.idinstr_17_bF$buf8 ),
    .C(_5790_),
    .Y(_5791_)
);

INVX1 _16430_ (
    .A(\datapath.registers.838[8] [0]),
    .Y(_5792_)
);

AOI21X1 _16431_ (
    .A(\datapath.registers.838[12] [0]),
    .B(\datapath.idinstr_17_bF$buf7 ),
    .C(\datapath.idinstr_15_bF$buf42 ),
    .Y(_5793_)
);

OAI21X1 _16432_ (
    .A(_5792_),
    .B(\datapath.idinstr_17_bF$buf6 ),
    .C(_5793_),
    .Y(_5794_)
);

NAND3X1 _16433_ (
    .A(_5756__bF$buf7),
    .B(_5794_),
    .C(_5791_),
    .Y(_5795_)
);

INVX1 _16434_ (
    .A(\datapath.registers.838[11] [0]),
    .Y(_5796_)
);

AOI21X1 _16435_ (
    .A(\datapath.registers.838[15] [0]),
    .B(\datapath.idinstr_17_bF$buf5 ),
    .C(_5762__bF$buf41),
    .Y(_5797_)
);

OAI21X1 _16436_ (
    .A(_5796_),
    .B(\datapath.idinstr_17_bF$buf4 ),
    .C(_5797_),
    .Y(_5798_)
);

AOI21X1 _16437_ (
    .A(\datapath.registers.838[14] [0]),
    .B(\datapath.idinstr_17_bF$buf3 ),
    .C(\datapath.idinstr_15_bF$buf41 ),
    .Y(_5799_)
);

OAI21X1 _16438_ (
    .A(_5219_),
    .B(\datapath.idinstr_17_bF$buf2 ),
    .C(_5799_),
    .Y(_5800_)
);

NAND3X1 _16439_ (
    .A(\datapath.idinstr_16_bF$buf40 ),
    .B(_5800_),
    .C(_5798_),
    .Y(_5801_)
);

AOI21X1 _16440_ (
    .A(_5795_),
    .B(_5801_),
    .C(_5760__bF$buf6),
    .Y(_5802_)
);

MUX2X1 _16441_ (
    .A(\datapath.registers.838[1] [0]),
    .B(\datapath.registers.838[0] [0]),
    .S(\datapath.idinstr_15_bF$buf40 ),
    .Y(_5803_)
);

NOR2X1 _16442_ (
    .A(\datapath.registers.838[3] [0]),
    .B(_5762__bF$buf40),
    .Y(_5804_)
);

OAI21X1 _16443_ (
    .A(\datapath.registers.838[2] [0]),
    .B(\datapath.idinstr_15_bF$buf39 ),
    .C(\datapath.idinstr_16_bF$buf39 ),
    .Y(_5805_)
);

OAI22X1 _16444_ (
    .A(_5805_),
    .B(_5804_),
    .C(\datapath.idinstr_16_bF$buf38 ),
    .D(_5803_),
    .Y(_5806_)
);

NAND2X1 _16445_ (
    .A(_5757__bF$buf7),
    .B(_5806_),
    .Y(_5807_)
);

MUX2X1 _16446_ (
    .A(\datapath.registers.838[5] [0]),
    .B(\datapath.registers.838[4] [0]),
    .S(\datapath.idinstr_15_bF$buf38 ),
    .Y(_5808_)
);

NOR2X1 _16447_ (
    .A(\datapath.registers.838[7] [0]),
    .B(_5762__bF$buf39),
    .Y(_5809_)
);

OAI21X1 _16448_ (
    .A(\datapath.registers.838[6] [0]),
    .B(\datapath.idinstr_15_bF$buf37 ),
    .C(\datapath.idinstr_16_bF$buf37 ),
    .Y(_5810_)
);

OAI22X1 _16449_ (
    .A(_5810_),
    .B(_5809_),
    .C(\datapath.idinstr_16_bF$buf36 ),
    .D(_5808_),
    .Y(_5811_)
);

NAND2X1 _16450_ (
    .A(\datapath.idinstr_17_bF$buf1 ),
    .B(_5811_),
    .Y(_5812_)
);

AOI21X1 _16451_ (
    .A(_5807_),
    .B(_5812_),
    .C(\datapath.idinstr_18_bF$buf0 ),
    .Y(_5813_)
);

OAI21X1 _16452_ (
    .A(_5802_),
    .B(_5813_),
    .C(_5789__bF$buf4),
    .Y(_5814_)
);

AOI22X1 _16453_ (
    .A(_5755__bF$buf4),
    .B(_5759__bF$buf4),
    .C(_5788_),
    .D(_5814_),
    .Y(\datapath.registers.rega_data [0])
);

MUX2X1 _16454_ (
    .A(\datapath.registers.838[9] [1]),
    .B(\datapath.registers.838[8] [1]),
    .S(\datapath.idinstr_15_bF$buf36 ),
    .Y(_5815_)
);

NOR2X1 _16455_ (
    .A(\datapath.registers.838[11] [1]),
    .B(_5762__bF$buf38),
    .Y(_5816_)
);

OAI21X1 _16456_ (
    .A(\datapath.registers.838[10] [1]),
    .B(\datapath.idinstr_15_bF$buf35 ),
    .C(\datapath.idinstr_16_bF$buf35 ),
    .Y(_5817_)
);

OAI22X1 _16457_ (
    .A(_5817_),
    .B(_5816_),
    .C(\datapath.idinstr_16_bF$buf34 ),
    .D(_5815_),
    .Y(_5818_)
);

INVX1 _16458_ (
    .A(\datapath.registers.838[15] [1]),
    .Y(_5819_)
);

AOI21X1 _16459_ (
    .A(_5762__bF$buf37),
    .B(\datapath.registers.838[14] [1]),
    .C(_5756__bF$buf6),
    .Y(_5820_)
);

OAI21X1 _16460_ (
    .A(_5819_),
    .B(_5762__bF$buf36),
    .C(_5820_),
    .Y(_5821_)
);

NAND2X1 _16461_ (
    .A(\datapath.registers.838[12] [1]),
    .B(_5762__bF$buf35),
    .Y(_5822_)
);

AOI21X1 _16462_ (
    .A(\datapath.registers.838[13] [1]),
    .B(\datapath.idinstr_15_bF$buf34 ),
    .C(\datapath.idinstr_16_bF$buf33 ),
    .Y(_5823_)
);

AOI21X1 _16463_ (
    .A(_5822_),
    .B(_5823_),
    .C(_5757__bF$buf6),
    .Y(_5824_)
);

AOI22X1 _16464_ (
    .A(_5821_),
    .B(_5824_),
    .C(_5757__bF$buf5),
    .D(_5818_),
    .Y(_5825_)
);

NOR2X1 _16465_ (
    .A(\datapath.registers.838[0] [1]),
    .B(\datapath.idinstr_15_bF$buf33 ),
    .Y(_5826_)
);

OAI21X1 _16466_ (
    .A(\datapath.registers.838[1] [1]),
    .B(_5762__bF$buf34),
    .C(_5756__bF$buf5),
    .Y(_5827_)
);

NOR2X1 _16467_ (
    .A(\datapath.registers.838[3] [1]),
    .B(_5762__bF$buf33),
    .Y(_5828_)
);

OAI21X1 _16468_ (
    .A(\datapath.registers.838[2] [1]),
    .B(\datapath.idinstr_15_bF$buf32 ),
    .C(\datapath.idinstr_16_bF$buf32 ),
    .Y(_5829_)
);

OAI22X1 _16469_ (
    .A(_5828_),
    .B(_5829_),
    .C(_5826_),
    .D(_5827_),
    .Y(_5830_)
);

NOR2X1 _16470_ (
    .A(\datapath.idinstr_17_bF$buf0 ),
    .B(_5830_),
    .Y(_5831_)
);

MUX2X1 _16471_ (
    .A(\datapath.registers.838[5] [1]),
    .B(\datapath.registers.838[4] [1]),
    .S(\datapath.idinstr_15_bF$buf31 ),
    .Y(_5832_)
);

NOR2X1 _16472_ (
    .A(\datapath.registers.838[7] [1]),
    .B(_5762__bF$buf32),
    .Y(_5833_)
);

OAI21X1 _16473_ (
    .A(\datapath.registers.838[6] [1]),
    .B(\datapath.idinstr_15_bF$buf30 ),
    .C(\datapath.idinstr_16_bF$buf31 ),
    .Y(_5834_)
);

OAI22X1 _16474_ (
    .A(_5834_),
    .B(_5833_),
    .C(\datapath.idinstr_16_bF$buf30 ),
    .D(_5832_),
    .Y(_5835_)
);

OAI21X1 _16475_ (
    .A(_5757__bF$buf4),
    .B(_5835_),
    .C(_5760__bF$buf5),
    .Y(_5836_)
);

OAI22X1 _16476_ (
    .A(_5760__bF$buf4),
    .B(_5825_),
    .C(_5831_),
    .D(_5836_),
    .Y(_5837_)
);

NAND2X1 _16477_ (
    .A(_5789__bF$buf3),
    .B(_5837_),
    .Y(_5838_)
);

INVX1 _16478_ (
    .A(\datapath.registers.838[27] [1]),
    .Y(_5839_)
);

AOI21X1 _16479_ (
    .A(\datapath.registers.838[31] [1]),
    .B(\datapath.idinstr_17_bF$buf15 ),
    .C(_5762__bF$buf31),
    .Y(_5840_)
);

OAI21X1 _16480_ (
    .A(\datapath.idinstr_17_bF$buf14 ),
    .B(_5839_),
    .C(_5840_),
    .Y(_5841_)
);

INVX1 _16481_ (
    .A(\datapath.registers.838[26] [1]),
    .Y(_5842_)
);

AOI21X1 _16482_ (
    .A(\datapath.registers.838[30] [1]),
    .B(\datapath.idinstr_17_bF$buf13 ),
    .C(\datapath.idinstr_15_bF$buf29 ),
    .Y(_5843_)
);

OAI21X1 _16483_ (
    .A(\datapath.idinstr_17_bF$buf12 ),
    .B(_5842_),
    .C(_5843_),
    .Y(_5844_)
);

NAND3X1 _16484_ (
    .A(\datapath.idinstr_16_bF$buf29 ),
    .B(_5844_),
    .C(_5841_),
    .Y(_5845_)
);

INVX1 _16485_ (
    .A(\datapath.registers.838[25] [1]),
    .Y(_5846_)
);

AOI21X1 _16486_ (
    .A(\datapath.idinstr_17_bF$buf11 ),
    .B(\datapath.registers.838[29] [1]),
    .C(_5762__bF$buf30),
    .Y(_5847_)
);

OAI21X1 _16487_ (
    .A(\datapath.idinstr_17_bF$buf10 ),
    .B(_5846_),
    .C(_5847_),
    .Y(_5848_)
);

INVX1 _16488_ (
    .A(\datapath.registers.838[24] [1]),
    .Y(_5849_)
);

AOI21X1 _16489_ (
    .A(\datapath.idinstr_17_bF$buf9 ),
    .B(\datapath.registers.838[28] [1]),
    .C(\datapath.idinstr_15_bF$buf28 ),
    .Y(_5850_)
);

OAI21X1 _16490_ (
    .A(_5849_),
    .B(\datapath.idinstr_17_bF$buf8 ),
    .C(_5850_),
    .Y(_5851_)
);

NAND3X1 _16491_ (
    .A(_5756__bF$buf4),
    .B(_5851_),
    .C(_5848_),
    .Y(_5852_)
);

AOI21X1 _16492_ (
    .A(_5845_),
    .B(_5852_),
    .C(_5760__bF$buf3),
    .Y(_5853_)
);

MUX2X1 _16493_ (
    .A(\datapath.registers.838[18] [1]),
    .B(\datapath.registers.838[16] [1]),
    .S(\datapath.idinstr_16_bF$buf28 ),
    .Y(_5854_)
);

NAND2X1 _16494_ (
    .A(_5762__bF$buf29),
    .B(_5854_),
    .Y(_5855_)
);

MUX2X1 _16495_ (
    .A(\datapath.registers.838[19] [1]),
    .B(\datapath.registers.838[17] [1]),
    .S(\datapath.idinstr_16_bF$buf27 ),
    .Y(_5856_)
);

NAND2X1 _16496_ (
    .A(\datapath.idinstr_15_bF$buf27 ),
    .B(_5856_),
    .Y(_5857_)
);

NAND3X1 _16497_ (
    .A(_5757__bF$buf3),
    .B(_5855_),
    .C(_5857_),
    .Y(_5858_)
);

MUX2X1 _16498_ (
    .A(\datapath.registers.838[22] [1]),
    .B(\datapath.registers.838[20] [1]),
    .S(\datapath.idinstr_16_bF$buf26 ),
    .Y(_5859_)
);

NAND2X1 _16499_ (
    .A(_5762__bF$buf28),
    .B(_5859_),
    .Y(_5860_)
);

MUX2X1 _16500_ (
    .A(\datapath.registers.838[23] [1]),
    .B(\datapath.registers.838[21] [1]),
    .S(\datapath.idinstr_16_bF$buf25 ),
    .Y(_5861_)
);

NAND2X1 _16501_ (
    .A(\datapath.idinstr_15_bF$buf26 ),
    .B(_5861_),
    .Y(_5862_)
);

NAND3X1 _16502_ (
    .A(\datapath.idinstr_17_bF$buf7 ),
    .B(_5860_),
    .C(_5862_),
    .Y(_5863_)
);

AOI21X1 _16503_ (
    .A(_5858_),
    .B(_5863_),
    .C(\datapath.idinstr_18_bF$buf6 ),
    .Y(_5864_)
);

OAI21X1 _16504_ (
    .A(_5853_),
    .B(_5864_),
    .C(\datapath.idinstr_19_bF$buf5 ),
    .Y(_5865_)
);

AOI22X1 _16505_ (
    .A(_5755__bF$buf3),
    .B(_5759__bF$buf3),
    .C(_5865_),
    .D(_5838_),
    .Y(\datapath.registers.rega_data [1])
);

NAND2X1 _16506_ (
    .A(\datapath.idinstr_15_bF$buf25 ),
    .B(\datapath.registers.838[27] [2]),
    .Y(_5866_)
);

NAND2X1 _16507_ (
    .A(\datapath.registers.838[26] [2]),
    .B(_5762__bF$buf27),
    .Y(_5867_)
);

NAND3X1 _16508_ (
    .A(\datapath.idinstr_16_bF$buf24 ),
    .B(_5866_),
    .C(_5867_),
    .Y(_5868_)
);

NAND2X1 _16509_ (
    .A(\datapath.idinstr_15_bF$buf24 ),
    .B(\datapath.registers.838[25] [2]),
    .Y(_5869_)
);

AOI21X1 _16510_ (
    .A(_5762__bF$buf26),
    .B(\datapath.registers.838[24] [2]),
    .C(\datapath.idinstr_16_bF$buf23 ),
    .Y(_5870_)
);

NAND2X1 _16511_ (
    .A(_5869_),
    .B(_5870_),
    .Y(_5871_)
);

NAND3X1 _16512_ (
    .A(_5757__bF$buf2),
    .B(_5868_),
    .C(_5871_),
    .Y(_5872_)
);

NAND2X1 _16513_ (
    .A(\datapath.registers.838[31] [2]),
    .B(\datapath.idinstr_15_bF$buf23 ),
    .Y(_5873_)
);

AOI21X1 _16514_ (
    .A(_5762__bF$buf25),
    .B(\datapath.registers.838[30] [2]),
    .C(_5756__bF$buf3),
    .Y(_5874_)
);

NAND2X1 _16515_ (
    .A(_5873_),
    .B(_5874_),
    .Y(_5875_)
);

INVX1 _16516_ (
    .A(\datapath.registers.838[28] [2]),
    .Y(_5876_)
);

AOI21X1 _16517_ (
    .A(\datapath.idinstr_15_bF$buf22 ),
    .B(\datapath.registers.838[29] [2]),
    .C(\datapath.idinstr_16_bF$buf22 ),
    .Y(_5877_)
);

OAI21X1 _16518_ (
    .A(\datapath.idinstr_15_bF$buf21 ),
    .B(_5876_),
    .C(_5877_),
    .Y(_5878_)
);

NAND3X1 _16519_ (
    .A(\datapath.idinstr_17_bF$buf6 ),
    .B(_5878_),
    .C(_5875_),
    .Y(_5879_)
);

AOI21X1 _16520_ (
    .A(_5872_),
    .B(_5879_),
    .C(_5760__bF$buf2),
    .Y(_5880_)
);

MUX2X1 _16521_ (
    .A(\datapath.registers.838[18] [2]),
    .B(\datapath.registers.838[16] [2]),
    .S(\datapath.idinstr_16_bF$buf21 ),
    .Y(_5881_)
);

NAND2X1 _16522_ (
    .A(_5762__bF$buf24),
    .B(_5881_),
    .Y(_5882_)
);

MUX2X1 _16523_ (
    .A(\datapath.registers.838[19] [2]),
    .B(\datapath.registers.838[17] [2]),
    .S(\datapath.idinstr_16_bF$buf20 ),
    .Y(_5883_)
);

NAND2X1 _16524_ (
    .A(\datapath.idinstr_15_bF$buf20 ),
    .B(_5883_),
    .Y(_5884_)
);

NAND3X1 _16525_ (
    .A(_5757__bF$buf1),
    .B(_5882_),
    .C(_5884_),
    .Y(_5885_)
);

MUX2X1 _16526_ (
    .A(\datapath.registers.838[22] [2]),
    .B(\datapath.registers.838[20] [2]),
    .S(\datapath.idinstr_16_bF$buf19 ),
    .Y(_5886_)
);

NAND2X1 _16527_ (
    .A(_5762__bF$buf23),
    .B(_5886_),
    .Y(_5887_)
);

MUX2X1 _16528_ (
    .A(\datapath.registers.838[23] [2]),
    .B(\datapath.registers.838[21] [2]),
    .S(\datapath.idinstr_16_bF$buf18 ),
    .Y(_5888_)
);

NAND2X1 _16529_ (
    .A(\datapath.idinstr_15_bF$buf19 ),
    .B(_5888_),
    .Y(_5889_)
);

NAND3X1 _16530_ (
    .A(\datapath.idinstr_17_bF$buf5 ),
    .B(_5887_),
    .C(_5889_),
    .Y(_5890_)
);

AOI21X1 _16531_ (
    .A(_5885_),
    .B(_5890_),
    .C(\datapath.idinstr_18_bF$buf5 ),
    .Y(_5891_)
);

OAI21X1 _16532_ (
    .A(_5891_),
    .B(_5880_),
    .C(\datapath.idinstr_19_bF$buf4 ),
    .Y(_5892_)
);

MUX2X1 _16533_ (
    .A(\datapath.registers.838[9] [2]),
    .B(\datapath.registers.838[8] [2]),
    .S(\datapath.idinstr_15_bF$buf18 ),
    .Y(_5893_)
);

NOR2X1 _16534_ (
    .A(\datapath.registers.838[11] [2]),
    .B(_5762__bF$buf22),
    .Y(_5894_)
);

OAI21X1 _16535_ (
    .A(\datapath.registers.838[10] [2]),
    .B(\datapath.idinstr_15_bF$buf17 ),
    .C(\datapath.idinstr_16_bF$buf17 ),
    .Y(_5895_)
);

OAI22X1 _16536_ (
    .A(_5895_),
    .B(_5894_),
    .C(\datapath.idinstr_16_bF$buf16 ),
    .D(_5893_),
    .Y(_5896_)
);

INVX1 _16537_ (
    .A(\datapath.registers.838[15] [2]),
    .Y(_5897_)
);

AOI21X1 _16538_ (
    .A(_5762__bF$buf21),
    .B(\datapath.registers.838[14] [2]),
    .C(_5756__bF$buf2),
    .Y(_5898_)
);

OAI21X1 _16539_ (
    .A(_5897_),
    .B(_5762__bF$buf20),
    .C(_5898_),
    .Y(_5899_)
);

NAND2X1 _16540_ (
    .A(\datapath.registers.838[12] [2]),
    .B(_5762__bF$buf19),
    .Y(_5900_)
);

AOI21X1 _16541_ (
    .A(\datapath.registers.838[13] [2]),
    .B(\datapath.idinstr_15_bF$buf16 ),
    .C(\datapath.idinstr_16_bF$buf15 ),
    .Y(_5901_)
);

AOI21X1 _16542_ (
    .A(_5900_),
    .B(_5901_),
    .C(_5757__bF$buf0),
    .Y(_5902_)
);

AOI22X1 _16543_ (
    .A(_5899_),
    .B(_5902_),
    .C(_5757__bF$buf10),
    .D(_5896_),
    .Y(_5903_)
);

NOR2X1 _16544_ (
    .A(\datapath.registers.838[0] [2]),
    .B(\datapath.idinstr_15_bF$buf15 ),
    .Y(_5904_)
);

OAI21X1 _16545_ (
    .A(\datapath.registers.838[1] [2]),
    .B(_5762__bF$buf18),
    .C(_5756__bF$buf1),
    .Y(_5905_)
);

NOR2X1 _16546_ (
    .A(\datapath.registers.838[3] [2]),
    .B(_5762__bF$buf17),
    .Y(_5906_)
);

OAI21X1 _16547_ (
    .A(\datapath.registers.838[2] [2]),
    .B(\datapath.idinstr_15_bF$buf14 ),
    .C(\datapath.idinstr_16_bF$buf14 ),
    .Y(_5907_)
);

OAI22X1 _16548_ (
    .A(_5906_),
    .B(_5907_),
    .C(_5904_),
    .D(_5905_),
    .Y(_5908_)
);

NOR2X1 _16549_ (
    .A(\datapath.idinstr_17_bF$buf4 ),
    .B(_5908_),
    .Y(_5909_)
);

MUX2X1 _16550_ (
    .A(\datapath.registers.838[5] [2]),
    .B(\datapath.registers.838[4] [2]),
    .S(\datapath.idinstr_15_bF$buf13 ),
    .Y(_5910_)
);

NOR2X1 _16551_ (
    .A(\datapath.registers.838[7] [2]),
    .B(_5762__bF$buf16),
    .Y(_5911_)
);

OAI21X1 _16552_ (
    .A(\datapath.registers.838[6] [2]),
    .B(\datapath.idinstr_15_bF$buf12 ),
    .C(\datapath.idinstr_16_bF$buf13 ),
    .Y(_5912_)
);

OAI22X1 _16553_ (
    .A(_5912_),
    .B(_5911_),
    .C(\datapath.idinstr_16_bF$buf12 ),
    .D(_5910_),
    .Y(_5913_)
);

OAI21X1 _16554_ (
    .A(_5757__bF$buf9),
    .B(_5913_),
    .C(_5760__bF$buf1),
    .Y(_5914_)
);

OAI22X1 _16555_ (
    .A(_5760__bF$buf0),
    .B(_5903_),
    .C(_5909_),
    .D(_5914_),
    .Y(_5915_)
);

NAND2X1 _16556_ (
    .A(_5789__bF$buf2),
    .B(_5915_),
    .Y(_5916_)
);

AOI22X1 _16557_ (
    .A(_5755__bF$buf2),
    .B(_5759__bF$buf2),
    .C(_5892_),
    .D(_5916_),
    .Y(\datapath.registers.rega_data [2])
);

MUX2X1 _16558_ (
    .A(\datapath.registers.838[2] [3]),
    .B(\datapath.registers.838[0] [3]),
    .S(\datapath.idinstr_16_bF$buf11 ),
    .Y(_5917_)
);

NAND2X1 _16559_ (
    .A(_5762__bF$buf15),
    .B(_5917_),
    .Y(_5918_)
);

MUX2X1 _16560_ (
    .A(\datapath.registers.838[3] [3]),
    .B(\datapath.registers.838[1] [3]),
    .S(\datapath.idinstr_16_bF$buf10 ),
    .Y(_5919_)
);

NAND2X1 _16561_ (
    .A(\datapath.idinstr_15_bF$buf11 ),
    .B(_5919_),
    .Y(_5920_)
);

NAND3X1 _16562_ (
    .A(_5757__bF$buf8),
    .B(_5918_),
    .C(_5920_),
    .Y(_5921_)
);

MUX2X1 _16563_ (
    .A(\datapath.registers.838[6] [3]),
    .B(\datapath.registers.838[4] [3]),
    .S(\datapath.idinstr_16_bF$buf9 ),
    .Y(_5922_)
);

NAND2X1 _16564_ (
    .A(_5762__bF$buf14),
    .B(_5922_),
    .Y(_5923_)
);

MUX2X1 _16565_ (
    .A(\datapath.registers.838[7] [3]),
    .B(\datapath.registers.838[5] [3]),
    .S(\datapath.idinstr_16_bF$buf8 ),
    .Y(_5924_)
);

NAND2X1 _16566_ (
    .A(\datapath.idinstr_15_bF$buf10 ),
    .B(_5924_),
    .Y(_5925_)
);

NAND3X1 _16567_ (
    .A(\datapath.idinstr_17_bF$buf3 ),
    .B(_5923_),
    .C(_5925_),
    .Y(_5926_)
);

AOI21X1 _16568_ (
    .A(_5921_),
    .B(_5926_),
    .C(\datapath.idinstr_18_bF$buf4 ),
    .Y(_5927_)
);

AOI21X1 _16569_ (
    .A(\datapath.registers.838[13] [3]),
    .B(\datapath.idinstr_17_bF$buf2 ),
    .C(_5762__bF$buf13),
    .Y(_5928_)
);

OAI21X1 _16570_ (
    .A(_5269_),
    .B(\datapath.idinstr_17_bF$buf1 ),
    .C(_5928_),
    .Y(_5929_)
);

INVX1 _16571_ (
    .A(\datapath.registers.838[8] [3]),
    .Y(_5930_)
);

AOI21X1 _16572_ (
    .A(\datapath.registers.838[12] [3]),
    .B(\datapath.idinstr_17_bF$buf0 ),
    .C(\datapath.idinstr_15_bF$buf9 ),
    .Y(_5931_)
);

OAI21X1 _16573_ (
    .A(_5930_),
    .B(\datapath.idinstr_17_bF$buf15 ),
    .C(_5931_),
    .Y(_5932_)
);

NAND3X1 _16574_ (
    .A(_5756__bF$buf0),
    .B(_5932_),
    .C(_5929_),
    .Y(_5933_)
);

INVX1 _16575_ (
    .A(\datapath.registers.838[11] [3]),
    .Y(_5934_)
);

AOI21X1 _16576_ (
    .A(\datapath.registers.838[15] [3]),
    .B(\datapath.idinstr_17_bF$buf14 ),
    .C(_5762__bF$buf12),
    .Y(_5935_)
);

OAI21X1 _16577_ (
    .A(_5934_),
    .B(\datapath.idinstr_17_bF$buf13 ),
    .C(_5935_),
    .Y(_5936_)
);

AOI21X1 _16578_ (
    .A(\datapath.registers.838[14] [3]),
    .B(\datapath.idinstr_17_bF$buf12 ),
    .C(\datapath.idinstr_15_bF$buf8 ),
    .Y(_5937_)
);

OAI21X1 _16579_ (
    .A(_5225_),
    .B(\datapath.idinstr_17_bF$buf11 ),
    .C(_5937_),
    .Y(_5938_)
);

NAND3X1 _16580_ (
    .A(\datapath.idinstr_16_bF$buf7 ),
    .B(_5938_),
    .C(_5936_),
    .Y(_5939_)
);

AOI21X1 _16581_ (
    .A(_5933_),
    .B(_5939_),
    .C(_5760__bF$buf7),
    .Y(_5940_)
);

OAI21X1 _16582_ (
    .A(_5940_),
    .B(_5927_),
    .C(_5789__bF$buf1),
    .Y(_5941_)
);

NOR2X1 _16583_ (
    .A(\datapath.registers.838[24] [3]),
    .B(\datapath.idinstr_15_bF$buf7 ),
    .Y(_5942_)
);

OAI21X1 _16584_ (
    .A(\datapath.registers.838[25] [3]),
    .B(_5762__bF$buf11),
    .C(_5756__bF$buf9),
    .Y(_5943_)
);

NOR2X1 _16585_ (
    .A(\datapath.registers.838[27] [3]),
    .B(_5762__bF$buf10),
    .Y(_5944_)
);

OAI21X1 _16586_ (
    .A(\datapath.idinstr_15_bF$buf6 ),
    .B(\datapath.registers.838[26] [3]),
    .C(\datapath.idinstr_16_bF$buf6 ),
    .Y(_5945_)
);

OAI22X1 _16587_ (
    .A(_5944_),
    .B(_5945_),
    .C(_5942_),
    .D(_5943_),
    .Y(_5946_)
);

NOR2X1 _16588_ (
    .A(\datapath.idinstr_17_bF$buf10 ),
    .B(_5946_),
    .Y(_5947_)
);

MUX2X1 _16589_ (
    .A(\datapath.registers.838[29] [3]),
    .B(\datapath.registers.838[28] [3]),
    .S(\datapath.idinstr_15_bF$buf5 ),
    .Y(_5948_)
);

NOR2X1 _16590_ (
    .A(\datapath.registers.838[31] [3]),
    .B(_5762__bF$buf9),
    .Y(_5949_)
);

OAI21X1 _16591_ (
    .A(\datapath.registers.838[30] [3]),
    .B(\datapath.idinstr_15_bF$buf4 ),
    .C(\datapath.idinstr_16_bF$buf5 ),
    .Y(_5950_)
);

OAI22X1 _16592_ (
    .A(_5950_),
    .B(_5949_),
    .C(\datapath.idinstr_16_bF$buf4 ),
    .D(_5948_),
    .Y(_5951_)
);

OAI21X1 _16593_ (
    .A(_5757__bF$buf7),
    .B(_5951_),
    .C(\datapath.idinstr_18_bF$buf3 ),
    .Y(_5952_)
);

INVX1 _16594_ (
    .A(\datapath.registers.838[19] [3]),
    .Y(_5953_)
);

AOI21X1 _16595_ (
    .A(\datapath.registers.838[23] [3]),
    .B(\datapath.idinstr_17_bF$buf9 ),
    .C(_5762__bF$buf8),
    .Y(_5954_)
);

OAI21X1 _16596_ (
    .A(_5953_),
    .B(\datapath.idinstr_17_bF$buf8 ),
    .C(_5954_),
    .Y(_5955_)
);

NAND2X1 _16597_ (
    .A(\datapath.registers.838[18] [3]),
    .B(_5757__bF$buf6),
    .Y(_5956_)
);

AOI21X1 _16598_ (
    .A(\datapath.registers.838[22] [3]),
    .B(\datapath.idinstr_17_bF$buf7 ),
    .C(\datapath.idinstr_15_bF$buf3 ),
    .Y(_5957_)
);

AOI21X1 _16599_ (
    .A(_5956_),
    .B(_5957_),
    .C(_5756__bF$buf8),
    .Y(_5958_)
);

AOI21X1 _16600_ (
    .A(\datapath.registers.838[21] [3]),
    .B(\datapath.idinstr_17_bF$buf6 ),
    .C(_5762__bF$buf7),
    .Y(_5959_)
);

OAI21X1 _16601_ (
    .A(_4973_),
    .B(\datapath.idinstr_17_bF$buf5 ),
    .C(_5959_),
    .Y(_5960_)
);

NAND2X1 _16602_ (
    .A(\datapath.registers.838[16] [3]),
    .B(_5757__bF$buf5),
    .Y(_5961_)
);

AOI21X1 _16603_ (
    .A(\datapath.registers.838[20] [3]),
    .B(\datapath.idinstr_17_bF$buf4 ),
    .C(\datapath.idinstr_15_bF$buf2 ),
    .Y(_5962_)
);

AOI21X1 _16604_ (
    .A(_5961_),
    .B(_5962_),
    .C(\datapath.idinstr_16_bF$buf3 ),
    .Y(_5963_)
);

AOI22X1 _16605_ (
    .A(_5958_),
    .B(_5955_),
    .C(_5960_),
    .D(_5963_),
    .Y(_5964_)
);

OAI22X1 _16606_ (
    .A(\datapath.idinstr_18_bF$buf2 ),
    .B(_5964_),
    .C(_5947_),
    .D(_5952_),
    .Y(_5965_)
);

NAND2X1 _16607_ (
    .A(\datapath.idinstr_19_bF$buf3 ),
    .B(_5965_),
    .Y(_5966_)
);

AOI22X1 _16608_ (
    .A(_5755__bF$buf1),
    .B(_5759__bF$buf1),
    .C(_5941_),
    .D(_5966_),
    .Y(\datapath.registers.rega_data [3])
);

NAND2X1 _16609_ (
    .A(\datapath.idinstr_15_bF$buf1 ),
    .B(\datapath.registers.838[27] [4]),
    .Y(_5967_)
);

NAND2X1 _16610_ (
    .A(\datapath.registers.838[26] [4]),
    .B(_5762__bF$buf6),
    .Y(_5968_)
);

NAND3X1 _16611_ (
    .A(\datapath.idinstr_16_bF$buf2 ),
    .B(_5967_),
    .C(_5968_),
    .Y(_5969_)
);

NAND2X1 _16612_ (
    .A(\datapath.idinstr_15_bF$buf0 ),
    .B(\datapath.registers.838[25] [4]),
    .Y(_5970_)
);

AOI21X1 _16613_ (
    .A(_5762__bF$buf5),
    .B(\datapath.registers.838[24] [4]),
    .C(\datapath.idinstr_16_bF$buf1 ),
    .Y(_5971_)
);

NAND2X1 _16614_ (
    .A(_5970_),
    .B(_5971_),
    .Y(_5972_)
);

NAND3X1 _16615_ (
    .A(_5757__bF$buf4),
    .B(_5969_),
    .C(_5972_),
    .Y(_5973_)
);

NAND2X1 _16616_ (
    .A(\datapath.registers.838[31] [4]),
    .B(\datapath.idinstr_15_bF$buf54 ),
    .Y(_5974_)
);

AOI21X1 _16617_ (
    .A(_5762__bF$buf4),
    .B(\datapath.registers.838[30] [4]),
    .C(_5756__bF$buf7),
    .Y(_5975_)
);

NAND2X1 _16618_ (
    .A(_5974_),
    .B(_5975_),
    .Y(_5976_)
);

INVX1 _16619_ (
    .A(\datapath.registers.838[28] [4]),
    .Y(_5977_)
);

AOI21X1 _16620_ (
    .A(\datapath.idinstr_15_bF$buf53 ),
    .B(\datapath.registers.838[29] [4]),
    .C(\datapath.idinstr_16_bF$buf0 ),
    .Y(_5978_)
);

OAI21X1 _16621_ (
    .A(\datapath.idinstr_15_bF$buf52 ),
    .B(_5977_),
    .C(_5978_),
    .Y(_5979_)
);

NAND3X1 _16622_ (
    .A(\datapath.idinstr_17_bF$buf3 ),
    .B(_5979_),
    .C(_5976_),
    .Y(_5980_)
);

AOI21X1 _16623_ (
    .A(_5973_),
    .B(_5980_),
    .C(_5760__bF$buf6),
    .Y(_5981_)
);

MUX2X1 _16624_ (
    .A(\datapath.registers.838[18] [4]),
    .B(\datapath.registers.838[16] [4]),
    .S(\datapath.idinstr_16_bF$buf51 ),
    .Y(_5982_)
);

NAND2X1 _16625_ (
    .A(_5762__bF$buf3),
    .B(_5982_),
    .Y(_5983_)
);

MUX2X1 _16626_ (
    .A(\datapath.registers.838[19] [4]),
    .B(\datapath.registers.838[17] [4]),
    .S(\datapath.idinstr_16_bF$buf50 ),
    .Y(_5984_)
);

NAND2X1 _16627_ (
    .A(\datapath.idinstr_15_bF$buf51 ),
    .B(_5984_),
    .Y(_5985_)
);

NAND3X1 _16628_ (
    .A(_5757__bF$buf3),
    .B(_5983_),
    .C(_5985_),
    .Y(_5986_)
);

MUX2X1 _16629_ (
    .A(\datapath.registers.838[22] [4]),
    .B(\datapath.registers.838[20] [4]),
    .S(\datapath.idinstr_16_bF$buf49 ),
    .Y(_5987_)
);

NAND2X1 _16630_ (
    .A(_5762__bF$buf2),
    .B(_5987_),
    .Y(_5988_)
);

MUX2X1 _16631_ (
    .A(\datapath.registers.838[23] [4]),
    .B(\datapath.registers.838[21] [4]),
    .S(\datapath.idinstr_16_bF$buf48 ),
    .Y(_5989_)
);

NAND2X1 _16632_ (
    .A(\datapath.idinstr_15_bF$buf50 ),
    .B(_5989_),
    .Y(_5990_)
);

NAND3X1 _16633_ (
    .A(\datapath.idinstr_17_bF$buf2 ),
    .B(_5988_),
    .C(_5990_),
    .Y(_5991_)
);

AOI21X1 _16634_ (
    .A(_5986_),
    .B(_5991_),
    .C(\datapath.idinstr_18_bF$buf1 ),
    .Y(_5992_)
);

OAI21X1 _16635_ (
    .A(_5992_),
    .B(_5981_),
    .C(\datapath.idinstr_19_bF$buf2 ),
    .Y(_5993_)
);

MUX2X1 _16636_ (
    .A(\datapath.registers.838[9] [4]),
    .B(\datapath.registers.838[8] [4]),
    .S(\datapath.idinstr_15_bF$buf49 ),
    .Y(_5994_)
);

NOR2X1 _16637_ (
    .A(\datapath.registers.838[11] [4]),
    .B(_5762__bF$buf1),
    .Y(_5995_)
);

OAI21X1 _16638_ (
    .A(\datapath.registers.838[10] [4]),
    .B(\datapath.idinstr_15_bF$buf48 ),
    .C(\datapath.idinstr_16_bF$buf47 ),
    .Y(_5996_)
);

OAI22X1 _16639_ (
    .A(_5996_),
    .B(_5995_),
    .C(\datapath.idinstr_16_bF$buf46 ),
    .D(_5994_),
    .Y(_5997_)
);

INVX1 _16640_ (
    .A(\datapath.registers.838[15] [4]),
    .Y(_5998_)
);

AOI21X1 _16641_ (
    .A(_5762__bF$buf0),
    .B(\datapath.registers.838[14] [4]),
    .C(_5756__bF$buf6),
    .Y(_5999_)
);

OAI21X1 _16642_ (
    .A(_5998_),
    .B(_5762__bF$buf47),
    .C(_5999_),
    .Y(_6000_)
);

NAND2X1 _16643_ (
    .A(\datapath.registers.838[12] [4]),
    .B(_5762__bF$buf46),
    .Y(_6001_)
);

AOI21X1 _16644_ (
    .A(\datapath.registers.838[13] [4]),
    .B(\datapath.idinstr_15_bF$buf47 ),
    .C(\datapath.idinstr_16_bF$buf45 ),
    .Y(_6002_)
);

AOI21X1 _16645_ (
    .A(_6001_),
    .B(_6002_),
    .C(_5757__bF$buf2),
    .Y(_6003_)
);

AOI22X1 _16646_ (
    .A(_6000_),
    .B(_6003_),
    .C(_5757__bF$buf1),
    .D(_5997_),
    .Y(_6004_)
);

NOR2X1 _16647_ (
    .A(\datapath.registers.838[0] [4]),
    .B(\datapath.idinstr_15_bF$buf46 ),
    .Y(_6005_)
);

OAI21X1 _16648_ (
    .A(\datapath.registers.838[1] [4]),
    .B(_5762__bF$buf45),
    .C(_5756__bF$buf5),
    .Y(_6006_)
);

NOR2X1 _16649_ (
    .A(\datapath.registers.838[3] [4]),
    .B(_5762__bF$buf44),
    .Y(_6007_)
);

OAI21X1 _16650_ (
    .A(\datapath.registers.838[2] [4]),
    .B(\datapath.idinstr_15_bF$buf45 ),
    .C(\datapath.idinstr_16_bF$buf44 ),
    .Y(_6008_)
);

OAI22X1 _16651_ (
    .A(_6007_),
    .B(_6008_),
    .C(_6005_),
    .D(_6006_),
    .Y(_6009_)
);

NOR2X1 _16652_ (
    .A(\datapath.idinstr_17_bF$buf1 ),
    .B(_6009_),
    .Y(_6010_)
);

MUX2X1 _16653_ (
    .A(\datapath.registers.838[5] [4]),
    .B(\datapath.registers.838[4] [4]),
    .S(\datapath.idinstr_15_bF$buf44 ),
    .Y(_6011_)
);

NOR2X1 _16654_ (
    .A(\datapath.registers.838[7] [4]),
    .B(_5762__bF$buf43),
    .Y(_6012_)
);

OAI21X1 _16655_ (
    .A(\datapath.registers.838[6] [4]),
    .B(\datapath.idinstr_15_bF$buf43 ),
    .C(\datapath.idinstr_16_bF$buf43 ),
    .Y(_6013_)
);

OAI22X1 _16656_ (
    .A(_6013_),
    .B(_6012_),
    .C(\datapath.idinstr_16_bF$buf42 ),
    .D(_6011_),
    .Y(_6014_)
);

OAI21X1 _16657_ (
    .A(_5757__bF$buf0),
    .B(_6014_),
    .C(_5760__bF$buf5),
    .Y(_6015_)
);

OAI22X1 _16658_ (
    .A(_5760__bF$buf4),
    .B(_6004_),
    .C(_6010_),
    .D(_6015_),
    .Y(_6016_)
);

NAND2X1 _16659_ (
    .A(_5789__bF$buf0),
    .B(_6016_),
    .Y(_6017_)
);

AOI22X1 _16660_ (
    .A(_5755__bF$buf0),
    .B(_5759__bF$buf0),
    .C(_5993_),
    .D(_6017_),
    .Y(\datapath.registers.rega_data [4])
);

MUX2X1 _16661_ (
    .A(\datapath.registers.838[9] [5]),
    .B(\datapath.registers.838[8] [5]),
    .S(\datapath.idinstr_15_bF$buf42 ),
    .Y(_6018_)
);

NOR2X1 _16662_ (
    .A(\datapath.registers.838[11] [5]),
    .B(_5762__bF$buf42),
    .Y(_6019_)
);

OAI21X1 _16663_ (
    .A(\datapath.registers.838[10] [5]),
    .B(\datapath.idinstr_15_bF$buf41 ),
    .C(\datapath.idinstr_16_bF$buf41 ),
    .Y(_6020_)
);

OAI22X1 _16664_ (
    .A(_6020_),
    .B(_6019_),
    .C(\datapath.idinstr_16_bF$buf40 ),
    .D(_6018_),
    .Y(_6021_)
);

INVX1 _16665_ (
    .A(\datapath.registers.838[15] [5]),
    .Y(_6022_)
);

AOI21X1 _16666_ (
    .A(_5762__bF$buf41),
    .B(\datapath.registers.838[14] [5]),
    .C(_5756__bF$buf4),
    .Y(_6023_)
);

OAI21X1 _16667_ (
    .A(_6022_),
    .B(_5762__bF$buf40),
    .C(_6023_),
    .Y(_6024_)
);

NAND2X1 _16668_ (
    .A(\datapath.registers.838[12] [5]),
    .B(_5762__bF$buf39),
    .Y(_6025_)
);

AOI21X1 _16669_ (
    .A(\datapath.registers.838[13] [5]),
    .B(\datapath.idinstr_15_bF$buf40 ),
    .C(\datapath.idinstr_16_bF$buf39 ),
    .Y(_6026_)
);

AOI21X1 _16670_ (
    .A(_6025_),
    .B(_6026_),
    .C(_5757__bF$buf10),
    .Y(_6027_)
);

AOI22X1 _16671_ (
    .A(_6024_),
    .B(_6027_),
    .C(_5757__bF$buf9),
    .D(_6021_),
    .Y(_6028_)
);

NOR2X1 _16672_ (
    .A(\datapath.registers.838[0] [5]),
    .B(\datapath.idinstr_15_bF$buf39 ),
    .Y(_6029_)
);

OAI21X1 _16673_ (
    .A(\datapath.registers.838[1] [5]),
    .B(_5762__bF$buf38),
    .C(_5756__bF$buf3),
    .Y(_6030_)
);

NOR2X1 _16674_ (
    .A(\datapath.registers.838[3] [5]),
    .B(_5762__bF$buf37),
    .Y(_6031_)
);

OAI21X1 _16675_ (
    .A(\datapath.registers.838[2] [5]),
    .B(\datapath.idinstr_15_bF$buf38 ),
    .C(\datapath.idinstr_16_bF$buf38 ),
    .Y(_6032_)
);

OAI22X1 _16676_ (
    .A(_6031_),
    .B(_6032_),
    .C(_6029_),
    .D(_6030_),
    .Y(_6033_)
);

NOR2X1 _16677_ (
    .A(\datapath.idinstr_17_bF$buf0 ),
    .B(_6033_),
    .Y(_6034_)
);

MUX2X1 _16678_ (
    .A(\datapath.registers.838[5] [5]),
    .B(\datapath.registers.838[4] [5]),
    .S(\datapath.idinstr_15_bF$buf37 ),
    .Y(_6035_)
);

NOR2X1 _16679_ (
    .A(\datapath.registers.838[7] [5]),
    .B(_5762__bF$buf36),
    .Y(_6036_)
);

OAI21X1 _16680_ (
    .A(\datapath.registers.838[6] [5]),
    .B(\datapath.idinstr_15_bF$buf36 ),
    .C(\datapath.idinstr_16_bF$buf37 ),
    .Y(_6037_)
);

OAI22X1 _16681_ (
    .A(_6037_),
    .B(_6036_),
    .C(\datapath.idinstr_16_bF$buf36 ),
    .D(_6035_),
    .Y(_6038_)
);

OAI21X1 _16682_ (
    .A(_5757__bF$buf8),
    .B(_6038_),
    .C(_5760__bF$buf3),
    .Y(_6039_)
);

OAI22X1 _16683_ (
    .A(_5760__bF$buf2),
    .B(_6028_),
    .C(_6034_),
    .D(_6039_),
    .Y(_6040_)
);

NAND2X1 _16684_ (
    .A(_5789__bF$buf4),
    .B(_6040_),
    .Y(_6041_)
);

INVX1 _16685_ (
    .A(\datapath.registers.838[27] [5]),
    .Y(_6042_)
);

AOI21X1 _16686_ (
    .A(\datapath.registers.838[31] [5]),
    .B(\datapath.idinstr_17_bF$buf15 ),
    .C(_5762__bF$buf35),
    .Y(_6043_)
);

OAI21X1 _16687_ (
    .A(\datapath.idinstr_17_bF$buf14 ),
    .B(_6042_),
    .C(_6043_),
    .Y(_6044_)
);

INVX1 _16688_ (
    .A(\datapath.registers.838[26] [5]),
    .Y(_6045_)
);

AOI21X1 _16689_ (
    .A(\datapath.registers.838[30] [5]),
    .B(\datapath.idinstr_17_bF$buf13 ),
    .C(\datapath.idinstr_15_bF$buf35 ),
    .Y(_6046_)
);

OAI21X1 _16690_ (
    .A(\datapath.idinstr_17_bF$buf12 ),
    .B(_6045_),
    .C(_6046_),
    .Y(_6047_)
);

NAND3X1 _16691_ (
    .A(\datapath.idinstr_16_bF$buf35 ),
    .B(_6047_),
    .C(_6044_),
    .Y(_6048_)
);

INVX1 _16692_ (
    .A(\datapath.registers.838[25] [5]),
    .Y(_6049_)
);

AOI21X1 _16693_ (
    .A(\datapath.idinstr_17_bF$buf11 ),
    .B(\datapath.registers.838[29] [5]),
    .C(_5762__bF$buf34),
    .Y(_6050_)
);

OAI21X1 _16694_ (
    .A(\datapath.idinstr_17_bF$buf10 ),
    .B(_6049_),
    .C(_6050_),
    .Y(_6051_)
);

INVX1 _16695_ (
    .A(\datapath.registers.838[24] [5]),
    .Y(_6052_)
);

AOI21X1 _16696_ (
    .A(\datapath.idinstr_17_bF$buf9 ),
    .B(\datapath.registers.838[28] [5]),
    .C(\datapath.idinstr_15_bF$buf34 ),
    .Y(_6053_)
);

OAI21X1 _16697_ (
    .A(_6052_),
    .B(\datapath.idinstr_17_bF$buf8 ),
    .C(_6053_),
    .Y(_6054_)
);

NAND3X1 _16698_ (
    .A(_5756__bF$buf2),
    .B(_6054_),
    .C(_6051_),
    .Y(_6055_)
);

AOI21X1 _16699_ (
    .A(_6048_),
    .B(_6055_),
    .C(_5760__bF$buf1),
    .Y(_6056_)
);

MUX2X1 _16700_ (
    .A(\datapath.registers.838[18] [5]),
    .B(\datapath.registers.838[16] [5]),
    .S(\datapath.idinstr_16_bF$buf34 ),
    .Y(_6057_)
);

NAND2X1 _16701_ (
    .A(_5762__bF$buf33),
    .B(_6057_),
    .Y(_6058_)
);

MUX2X1 _16702_ (
    .A(\datapath.registers.838[19] [5]),
    .B(\datapath.registers.838[17] [5]),
    .S(\datapath.idinstr_16_bF$buf33 ),
    .Y(_6059_)
);

NAND2X1 _16703_ (
    .A(\datapath.idinstr_15_bF$buf33 ),
    .B(_6059_),
    .Y(_6060_)
);

NAND3X1 _16704_ (
    .A(_5757__bF$buf7),
    .B(_6058_),
    .C(_6060_),
    .Y(_6061_)
);

MUX2X1 _16705_ (
    .A(\datapath.registers.838[22] [5]),
    .B(\datapath.registers.838[20] [5]),
    .S(\datapath.idinstr_16_bF$buf32 ),
    .Y(_6062_)
);

NAND2X1 _16706_ (
    .A(_5762__bF$buf32),
    .B(_6062_),
    .Y(_6063_)
);

MUX2X1 _16707_ (
    .A(\datapath.registers.838[23] [5]),
    .B(\datapath.registers.838[21] [5]),
    .S(\datapath.idinstr_16_bF$buf31 ),
    .Y(_6064_)
);

NAND2X1 _16708_ (
    .A(\datapath.idinstr_15_bF$buf32 ),
    .B(_6064_),
    .Y(_6065_)
);

NAND3X1 _16709_ (
    .A(\datapath.idinstr_17_bF$buf7 ),
    .B(_6063_),
    .C(_6065_),
    .Y(_6066_)
);

AOI21X1 _16710_ (
    .A(_6061_),
    .B(_6066_),
    .C(\datapath.idinstr_18_bF$buf0 ),
    .Y(_6067_)
);

OAI21X1 _16711_ (
    .A(_6056_),
    .B(_6067_),
    .C(\datapath.idinstr_19_bF$buf1 ),
    .Y(_6068_)
);

AOI22X1 _16712_ (
    .A(_5755__bF$buf4),
    .B(_5759__bF$buf4),
    .C(_6068_),
    .D(_6041_),
    .Y(\datapath.registers.rega_data [5])
);

MUX2X1 _16713_ (
    .A(\datapath.registers.838[2] [6]),
    .B(\datapath.registers.838[0] [6]),
    .S(\datapath.idinstr_16_bF$buf30 ),
    .Y(_6069_)
);

NAND2X1 _16714_ (
    .A(_5762__bF$buf31),
    .B(_6069_),
    .Y(_6070_)
);

MUX2X1 _16715_ (
    .A(\datapath.registers.838[3] [6]),
    .B(\datapath.registers.838[1] [6]),
    .S(\datapath.idinstr_16_bF$buf29 ),
    .Y(_6071_)
);

NAND2X1 _16716_ (
    .A(\datapath.idinstr_15_bF$buf31 ),
    .B(_6071_),
    .Y(_6072_)
);

NAND3X1 _16717_ (
    .A(_5757__bF$buf6),
    .B(_6070_),
    .C(_6072_),
    .Y(_6073_)
);

MUX2X1 _16718_ (
    .A(\datapath.registers.838[6] [6]),
    .B(\datapath.registers.838[4] [6]),
    .S(\datapath.idinstr_16_bF$buf28 ),
    .Y(_6074_)
);

NAND2X1 _16719_ (
    .A(_5762__bF$buf30),
    .B(_6074_),
    .Y(_6075_)
);

MUX2X1 _16720_ (
    .A(\datapath.registers.838[7] [6]),
    .B(\datapath.registers.838[5] [6]),
    .S(\datapath.idinstr_16_bF$buf27 ),
    .Y(_6076_)
);

NAND2X1 _16721_ (
    .A(\datapath.idinstr_15_bF$buf30 ),
    .B(_6076_),
    .Y(_6077_)
);

NAND3X1 _16722_ (
    .A(\datapath.idinstr_17_bF$buf6 ),
    .B(_6075_),
    .C(_6077_),
    .Y(_6078_)
);

AOI21X1 _16723_ (
    .A(_6073_),
    .B(_6078_),
    .C(\datapath.idinstr_18_bF$buf6 ),
    .Y(_6079_)
);

AOI21X1 _16724_ (
    .A(\datapath.registers.838[13] [6]),
    .B(\datapath.idinstr_17_bF$buf5 ),
    .C(_5762__bF$buf29),
    .Y(_6080_)
);

OAI21X1 _16725_ (
    .A(_5273_),
    .B(\datapath.idinstr_17_bF$buf4 ),
    .C(_6080_),
    .Y(_6081_)
);

INVX1 _16726_ (
    .A(\datapath.registers.838[8] [6]),
    .Y(_6082_)
);

AOI21X1 _16727_ (
    .A(\datapath.registers.838[12] [6]),
    .B(\datapath.idinstr_17_bF$buf3 ),
    .C(\datapath.idinstr_15_bF$buf29 ),
    .Y(_6083_)
);

OAI21X1 _16728_ (
    .A(_6082_),
    .B(\datapath.idinstr_17_bF$buf2 ),
    .C(_6083_),
    .Y(_6084_)
);

NAND3X1 _16729_ (
    .A(_5756__bF$buf1),
    .B(_6084_),
    .C(_6081_),
    .Y(_6085_)
);

INVX1 _16730_ (
    .A(\datapath.registers.838[11] [6]),
    .Y(_6086_)
);

AOI21X1 _16731_ (
    .A(\datapath.registers.838[15] [6]),
    .B(\datapath.idinstr_17_bF$buf1 ),
    .C(_5762__bF$buf28),
    .Y(_6087_)
);

OAI21X1 _16732_ (
    .A(_6086_),
    .B(\datapath.idinstr_17_bF$buf0 ),
    .C(_6087_),
    .Y(_6088_)
);

AOI21X1 _16733_ (
    .A(\datapath.registers.838[14] [6]),
    .B(\datapath.idinstr_17_bF$buf15 ),
    .C(\datapath.idinstr_15_bF$buf28 ),
    .Y(_6089_)
);

OAI21X1 _16734_ (
    .A(_5229_),
    .B(\datapath.idinstr_17_bF$buf14 ),
    .C(_6089_),
    .Y(_6090_)
);

NAND3X1 _16735_ (
    .A(\datapath.idinstr_16_bF$buf26 ),
    .B(_6090_),
    .C(_6088_),
    .Y(_6091_)
);

AOI21X1 _16736_ (
    .A(_6085_),
    .B(_6091_),
    .C(_5760__bF$buf0),
    .Y(_6092_)
);

OAI21X1 _16737_ (
    .A(_6092_),
    .B(_6079_),
    .C(_5789__bF$buf3),
    .Y(_6093_)
);

NOR2X1 _16738_ (
    .A(\datapath.registers.838[24] [6]),
    .B(\datapath.idinstr_15_bF$buf27 ),
    .Y(_6094_)
);

OAI21X1 _16739_ (
    .A(\datapath.registers.838[25] [6]),
    .B(_5762__bF$buf27),
    .C(_5756__bF$buf0),
    .Y(_6095_)
);

NOR2X1 _16740_ (
    .A(\datapath.registers.838[27] [6]),
    .B(_5762__bF$buf26),
    .Y(_6096_)
);

OAI21X1 _16741_ (
    .A(\datapath.idinstr_15_bF$buf26 ),
    .B(\datapath.registers.838[26] [6]),
    .C(\datapath.idinstr_16_bF$buf25 ),
    .Y(_6097_)
);

OAI22X1 _16742_ (
    .A(_6096_),
    .B(_6097_),
    .C(_6094_),
    .D(_6095_),
    .Y(_6098_)
);

NOR2X1 _16743_ (
    .A(\datapath.idinstr_17_bF$buf13 ),
    .B(_6098_),
    .Y(_6099_)
);

MUX2X1 _16744_ (
    .A(\datapath.registers.838[29] [6]),
    .B(\datapath.registers.838[28] [6]),
    .S(\datapath.idinstr_15_bF$buf25 ),
    .Y(_6100_)
);

NOR2X1 _16745_ (
    .A(\datapath.registers.838[31] [6]),
    .B(_5762__bF$buf25),
    .Y(_6101_)
);

OAI21X1 _16746_ (
    .A(\datapath.registers.838[30] [6]),
    .B(\datapath.idinstr_15_bF$buf24 ),
    .C(\datapath.idinstr_16_bF$buf24 ),
    .Y(_6102_)
);

OAI22X1 _16747_ (
    .A(_6102_),
    .B(_6101_),
    .C(\datapath.idinstr_16_bF$buf23 ),
    .D(_6100_),
    .Y(_6103_)
);

OAI21X1 _16748_ (
    .A(_5757__bF$buf5),
    .B(_6103_),
    .C(\datapath.idinstr_18_bF$buf5 ),
    .Y(_6104_)
);

INVX1 _16749_ (
    .A(\datapath.registers.838[19] [6]),
    .Y(_6105_)
);

AOI21X1 _16750_ (
    .A(\datapath.registers.838[23] [6]),
    .B(\datapath.idinstr_17_bF$buf12 ),
    .C(_5762__bF$buf24),
    .Y(_6106_)
);

OAI21X1 _16751_ (
    .A(_6105_),
    .B(\datapath.idinstr_17_bF$buf11 ),
    .C(_6106_),
    .Y(_6107_)
);

NAND2X1 _16752_ (
    .A(\datapath.registers.838[18] [6]),
    .B(_5757__bF$buf4),
    .Y(_6108_)
);

AOI21X1 _16753_ (
    .A(\datapath.registers.838[22] [6]),
    .B(\datapath.idinstr_17_bF$buf10 ),
    .C(\datapath.idinstr_15_bF$buf23 ),
    .Y(_6109_)
);

AOI21X1 _16754_ (
    .A(_6108_),
    .B(_6109_),
    .C(_5756__bF$buf9),
    .Y(_6110_)
);

AOI21X1 _16755_ (
    .A(\datapath.registers.838[21] [6]),
    .B(\datapath.idinstr_17_bF$buf9 ),
    .C(_5762__bF$buf23),
    .Y(_6111_)
);

OAI21X1 _16756_ (
    .A(_4979_),
    .B(\datapath.idinstr_17_bF$buf8 ),
    .C(_6111_),
    .Y(_6112_)
);

NAND2X1 _16757_ (
    .A(\datapath.registers.838[16] [6]),
    .B(_5757__bF$buf3),
    .Y(_6113_)
);

AOI21X1 _16758_ (
    .A(\datapath.registers.838[20] [6]),
    .B(\datapath.idinstr_17_bF$buf7 ),
    .C(\datapath.idinstr_15_bF$buf22 ),
    .Y(_6114_)
);

AOI21X1 _16759_ (
    .A(_6113_),
    .B(_6114_),
    .C(\datapath.idinstr_16_bF$buf22 ),
    .Y(_6115_)
);

AOI22X1 _16760_ (
    .A(_6110_),
    .B(_6107_),
    .C(_6112_),
    .D(_6115_),
    .Y(_6116_)
);

OAI22X1 _16761_ (
    .A(\datapath.idinstr_18_bF$buf4 ),
    .B(_6116_),
    .C(_6099_),
    .D(_6104_),
    .Y(_6117_)
);

NAND2X1 _16762_ (
    .A(\datapath.idinstr_19_bF$buf0 ),
    .B(_6117_),
    .Y(_6118_)
);

AOI22X1 _16763_ (
    .A(_5755__bF$buf3),
    .B(_5759__bF$buf3),
    .C(_6093_),
    .D(_6118_),
    .Y(\datapath.registers.rega_data [6])
);

MUX2X1 _16764_ (
    .A(\datapath.registers.838[9] [7]),
    .B(\datapath.registers.838[8] [7]),
    .S(\datapath.idinstr_15_bF$buf21 ),
    .Y(_6119_)
);

NOR2X1 _16765_ (
    .A(\datapath.registers.838[11] [7]),
    .B(_5762__bF$buf22),
    .Y(_6120_)
);

OAI21X1 _16766_ (
    .A(\datapath.registers.838[10] [7]),
    .B(\datapath.idinstr_15_bF$buf20 ),
    .C(\datapath.idinstr_16_bF$buf21 ),
    .Y(_6121_)
);

OAI22X1 _16767_ (
    .A(_6121_),
    .B(_6120_),
    .C(\datapath.idinstr_16_bF$buf20 ),
    .D(_6119_),
    .Y(_6122_)
);

INVX1 _16768_ (
    .A(\datapath.registers.838[15] [7]),
    .Y(_6123_)
);

AOI21X1 _16769_ (
    .A(_5762__bF$buf21),
    .B(\datapath.registers.838[14] [7]),
    .C(_5756__bF$buf8),
    .Y(_6124_)
);

OAI21X1 _16770_ (
    .A(_6123_),
    .B(_5762__bF$buf20),
    .C(_6124_),
    .Y(_6125_)
);

NAND2X1 _16771_ (
    .A(\datapath.registers.838[12] [7]),
    .B(_5762__bF$buf19),
    .Y(_6126_)
);

AOI21X1 _16772_ (
    .A(\datapath.registers.838[13] [7]),
    .B(\datapath.idinstr_15_bF$buf19 ),
    .C(\datapath.idinstr_16_bF$buf19 ),
    .Y(_6127_)
);

AOI21X1 _16773_ (
    .A(_6126_),
    .B(_6127_),
    .C(_5757__bF$buf2),
    .Y(_6128_)
);

AOI22X1 _16774_ (
    .A(_6125_),
    .B(_6128_),
    .C(_5757__bF$buf1),
    .D(_6122_),
    .Y(_6129_)
);

NOR2X1 _16775_ (
    .A(\datapath.registers.838[0] [7]),
    .B(\datapath.idinstr_15_bF$buf18 ),
    .Y(_6130_)
);

OAI21X1 _16776_ (
    .A(\datapath.registers.838[1] [7]),
    .B(_5762__bF$buf18),
    .C(_5756__bF$buf7),
    .Y(_6131_)
);

NOR2X1 _16777_ (
    .A(\datapath.registers.838[3] [7]),
    .B(_5762__bF$buf17),
    .Y(_6132_)
);

OAI21X1 _16778_ (
    .A(\datapath.registers.838[2] [7]),
    .B(\datapath.idinstr_15_bF$buf17 ),
    .C(\datapath.idinstr_16_bF$buf18 ),
    .Y(_6133_)
);

OAI22X1 _16779_ (
    .A(_6132_),
    .B(_6133_),
    .C(_6130_),
    .D(_6131_),
    .Y(_6134_)
);

NOR2X1 _16780_ (
    .A(\datapath.idinstr_17_bF$buf6 ),
    .B(_6134_),
    .Y(_6135_)
);

MUX2X1 _16781_ (
    .A(\datapath.registers.838[5] [7]),
    .B(\datapath.registers.838[4] [7]),
    .S(\datapath.idinstr_15_bF$buf16 ),
    .Y(_6136_)
);

NOR2X1 _16782_ (
    .A(\datapath.registers.838[7] [7]),
    .B(_5762__bF$buf16),
    .Y(_6137_)
);

OAI21X1 _16783_ (
    .A(\datapath.registers.838[6] [7]),
    .B(\datapath.idinstr_15_bF$buf15 ),
    .C(\datapath.idinstr_16_bF$buf17 ),
    .Y(_6138_)
);

OAI22X1 _16784_ (
    .A(_6138_),
    .B(_6137_),
    .C(\datapath.idinstr_16_bF$buf16 ),
    .D(_6136_),
    .Y(_6139_)
);

OAI21X1 _16785_ (
    .A(_5757__bF$buf0),
    .B(_6139_),
    .C(_5760__bF$buf7),
    .Y(_6140_)
);

OAI22X1 _16786_ (
    .A(_5760__bF$buf6),
    .B(_6129_),
    .C(_6135_),
    .D(_6140_),
    .Y(_6141_)
);

NAND2X1 _16787_ (
    .A(_5789__bF$buf2),
    .B(_6141_),
    .Y(_6142_)
);

INVX1 _16788_ (
    .A(\datapath.registers.838[27] [7]),
    .Y(_6143_)
);

AOI21X1 _16789_ (
    .A(\datapath.registers.838[31] [7]),
    .B(\datapath.idinstr_17_bF$buf5 ),
    .C(_5762__bF$buf15),
    .Y(_6144_)
);

OAI21X1 _16790_ (
    .A(\datapath.idinstr_17_bF$buf4 ),
    .B(_6143_),
    .C(_6144_),
    .Y(_6145_)
);

INVX1 _16791_ (
    .A(\datapath.registers.838[26] [7]),
    .Y(_6146_)
);

AOI21X1 _16792_ (
    .A(\datapath.registers.838[30] [7]),
    .B(\datapath.idinstr_17_bF$buf3 ),
    .C(\datapath.idinstr_15_bF$buf14 ),
    .Y(_6147_)
);

OAI21X1 _16793_ (
    .A(\datapath.idinstr_17_bF$buf2 ),
    .B(_6146_),
    .C(_6147_),
    .Y(_6148_)
);

NAND3X1 _16794_ (
    .A(\datapath.idinstr_16_bF$buf15 ),
    .B(_6148_),
    .C(_6145_),
    .Y(_6149_)
);

INVX1 _16795_ (
    .A(\datapath.registers.838[25] [7]),
    .Y(_6150_)
);

AOI21X1 _16796_ (
    .A(\datapath.idinstr_17_bF$buf1 ),
    .B(\datapath.registers.838[29] [7]),
    .C(_5762__bF$buf14),
    .Y(_6151_)
);

OAI21X1 _16797_ (
    .A(\datapath.idinstr_17_bF$buf0 ),
    .B(_6150_),
    .C(_6151_),
    .Y(_6152_)
);

INVX1 _16798_ (
    .A(\datapath.registers.838[24] [7]),
    .Y(_6153_)
);

AOI21X1 _16799_ (
    .A(\datapath.idinstr_17_bF$buf15 ),
    .B(\datapath.registers.838[28] [7]),
    .C(\datapath.idinstr_15_bF$buf13 ),
    .Y(_6154_)
);

OAI21X1 _16800_ (
    .A(_6153_),
    .B(\datapath.idinstr_17_bF$buf14 ),
    .C(_6154_),
    .Y(_6155_)
);

NAND3X1 _16801_ (
    .A(_5756__bF$buf6),
    .B(_6155_),
    .C(_6152_),
    .Y(_6156_)
);

AOI21X1 _16802_ (
    .A(_6149_),
    .B(_6156_),
    .C(_5760__bF$buf5),
    .Y(_6157_)
);

MUX2X1 _16803_ (
    .A(\datapath.registers.838[18] [7]),
    .B(\datapath.registers.838[16] [7]),
    .S(\datapath.idinstr_16_bF$buf14 ),
    .Y(_6158_)
);

NAND2X1 _16804_ (
    .A(_5762__bF$buf13),
    .B(_6158_),
    .Y(_6159_)
);

MUX2X1 _16805_ (
    .A(\datapath.registers.838[19] [7]),
    .B(\datapath.registers.838[17] [7]),
    .S(\datapath.idinstr_16_bF$buf13 ),
    .Y(_6160_)
);

NAND2X1 _16806_ (
    .A(\datapath.idinstr_15_bF$buf12 ),
    .B(_6160_),
    .Y(_6161_)
);

NAND3X1 _16807_ (
    .A(_5757__bF$buf10),
    .B(_6159_),
    .C(_6161_),
    .Y(_6162_)
);

MUX2X1 _16808_ (
    .A(\datapath.registers.838[22] [7]),
    .B(\datapath.registers.838[20] [7]),
    .S(\datapath.idinstr_16_bF$buf12 ),
    .Y(_6163_)
);

NAND2X1 _16809_ (
    .A(_5762__bF$buf12),
    .B(_6163_),
    .Y(_6164_)
);

MUX2X1 _16810_ (
    .A(\datapath.registers.838[23] [7]),
    .B(\datapath.registers.838[21] [7]),
    .S(\datapath.idinstr_16_bF$buf11 ),
    .Y(_6165_)
);

NAND2X1 _16811_ (
    .A(\datapath.idinstr_15_bF$buf11 ),
    .B(_6165_),
    .Y(_6166_)
);

NAND3X1 _16812_ (
    .A(\datapath.idinstr_17_bF$buf13 ),
    .B(_6164_),
    .C(_6166_),
    .Y(_6167_)
);

AOI21X1 _16813_ (
    .A(_6162_),
    .B(_6167_),
    .C(\datapath.idinstr_18_bF$buf3 ),
    .Y(_6168_)
);

OAI21X1 _16814_ (
    .A(_6157_),
    .B(_6168_),
    .C(\datapath.idinstr_19_bF$buf5 ),
    .Y(_6169_)
);

AOI22X1 _16815_ (
    .A(_5755__bF$buf2),
    .B(_5759__bF$buf2),
    .C(_6169_),
    .D(_6142_),
    .Y(\datapath.registers.rega_data [7])
);

NAND2X1 _16816_ (
    .A(\datapath.idinstr_15_bF$buf10 ),
    .B(\datapath.registers.838[27] [8]),
    .Y(_6170_)
);

NAND2X1 _16817_ (
    .A(\datapath.registers.838[26] [8]),
    .B(_5762__bF$buf11),
    .Y(_6171_)
);

NAND3X1 _16818_ (
    .A(\datapath.idinstr_16_bF$buf10 ),
    .B(_6170_),
    .C(_6171_),
    .Y(_6172_)
);

NAND2X1 _16819_ (
    .A(\datapath.idinstr_15_bF$buf9 ),
    .B(\datapath.registers.838[25] [8]),
    .Y(_6173_)
);

AOI21X1 _16820_ (
    .A(_5762__bF$buf10),
    .B(\datapath.registers.838[24] [8]),
    .C(\datapath.idinstr_16_bF$buf9 ),
    .Y(_6174_)
);

NAND2X1 _16821_ (
    .A(_6173_),
    .B(_6174_),
    .Y(_6175_)
);

NAND3X1 _16822_ (
    .A(_5757__bF$buf9),
    .B(_6172_),
    .C(_6175_),
    .Y(_6176_)
);

NAND2X1 _16823_ (
    .A(\datapath.registers.838[31] [8]),
    .B(\datapath.idinstr_15_bF$buf8 ),
    .Y(_6177_)
);

AOI21X1 _16824_ (
    .A(_5762__bF$buf9),
    .B(\datapath.registers.838[30] [8]),
    .C(_5756__bF$buf5),
    .Y(_6178_)
);

NAND2X1 _16825_ (
    .A(_6177_),
    .B(_6178_),
    .Y(_6179_)
);

INVX1 _16826_ (
    .A(\datapath.registers.838[28] [8]),
    .Y(_6180_)
);

AOI21X1 _16827_ (
    .A(\datapath.idinstr_15_bF$buf7 ),
    .B(\datapath.registers.838[29] [8]),
    .C(\datapath.idinstr_16_bF$buf8 ),
    .Y(_6181_)
);

OAI21X1 _16828_ (
    .A(\datapath.idinstr_15_bF$buf6 ),
    .B(_6180_),
    .C(_6181_),
    .Y(_6182_)
);

NAND3X1 _16829_ (
    .A(\datapath.idinstr_17_bF$buf12 ),
    .B(_6182_),
    .C(_6179_),
    .Y(_6183_)
);

AOI21X1 _16830_ (
    .A(_6176_),
    .B(_6183_),
    .C(_5760__bF$buf4),
    .Y(_6184_)
);

MUX2X1 _16831_ (
    .A(\datapath.registers.838[17] [8]),
    .B(\datapath.registers.838[16] [8]),
    .S(\datapath.idinstr_15_bF$buf5 ),
    .Y(_6185_)
);

NOR2X1 _16832_ (
    .A(\datapath.registers.838[19] [8]),
    .B(_5762__bF$buf8),
    .Y(_6186_)
);

OAI21X1 _16833_ (
    .A(\datapath.registers.838[18] [8]),
    .B(\datapath.idinstr_15_bF$buf4 ),
    .C(\datapath.idinstr_16_bF$buf7 ),
    .Y(_6187_)
);

OAI22X1 _16834_ (
    .A(_6187_),
    .B(_6186_),
    .C(\datapath.idinstr_16_bF$buf6 ),
    .D(_6185_),
    .Y(_6188_)
);

NAND2X1 _16835_ (
    .A(_5757__bF$buf8),
    .B(_6188_),
    .Y(_6189_)
);

MUX2X1 _16836_ (
    .A(\datapath.registers.838[21] [8]),
    .B(\datapath.registers.838[20] [8]),
    .S(\datapath.idinstr_15_bF$buf3 ),
    .Y(_6190_)
);

NOR2X1 _16837_ (
    .A(\datapath.registers.838[23] [8]),
    .B(_5762__bF$buf7),
    .Y(_6191_)
);

OAI21X1 _16838_ (
    .A(\datapath.registers.838[22] [8]),
    .B(\datapath.idinstr_15_bF$buf2 ),
    .C(\datapath.idinstr_16_bF$buf5 ),
    .Y(_6192_)
);

OAI22X1 _16839_ (
    .A(_6192_),
    .B(_6191_),
    .C(\datapath.idinstr_16_bF$buf4 ),
    .D(_6190_),
    .Y(_6193_)
);

NAND2X1 _16840_ (
    .A(\datapath.idinstr_17_bF$buf11 ),
    .B(_6193_),
    .Y(_6194_)
);

AOI21X1 _16841_ (
    .A(_6189_),
    .B(_6194_),
    .C(\datapath.idinstr_18_bF$buf2 ),
    .Y(_6195_)
);

OAI21X1 _16842_ (
    .A(_6184_),
    .B(_6195_),
    .C(\datapath.idinstr_19_bF$buf4 ),
    .Y(_6196_)
);

NAND2X1 _16843_ (
    .A(\datapath.registers.838[11] [8]),
    .B(\datapath.idinstr_16_bF$buf3 ),
    .Y(_6197_)
);

NAND2X1 _16844_ (
    .A(\datapath.registers.838[9] [8]),
    .B(_5756__bF$buf4),
    .Y(_6198_)
);

NAND3X1 _16845_ (
    .A(\datapath.idinstr_15_bF$buf1 ),
    .B(_6197_),
    .C(_6198_),
    .Y(_6199_)
);

NAND2X1 _16846_ (
    .A(\datapath.registers.838[10] [8]),
    .B(\datapath.idinstr_16_bF$buf2 ),
    .Y(_6200_)
);

AOI21X1 _16847_ (
    .A(_5756__bF$buf3),
    .B(\datapath.registers.838[8] [8]),
    .C(\datapath.idinstr_15_bF$buf0 ),
    .Y(_6201_)
);

NAND2X1 _16848_ (
    .A(_6200_),
    .B(_6201_),
    .Y(_6202_)
);

NAND3X1 _16849_ (
    .A(_5757__bF$buf7),
    .B(_6199_),
    .C(_6202_),
    .Y(_6203_)
);

NAND2X1 _16850_ (
    .A(\datapath.registers.838[15] [8]),
    .B(\datapath.idinstr_16_bF$buf1 ),
    .Y(_6204_)
);

NAND2X1 _16851_ (
    .A(\datapath.registers.838[13] [8]),
    .B(_5756__bF$buf2),
    .Y(_6205_)
);

NAND3X1 _16852_ (
    .A(\datapath.idinstr_15_bF$buf54 ),
    .B(_6204_),
    .C(_6205_),
    .Y(_6206_)
);

NAND2X1 _16853_ (
    .A(\datapath.registers.838[14] [8]),
    .B(\datapath.idinstr_16_bF$buf0 ),
    .Y(_6207_)
);

AOI21X1 _16854_ (
    .A(_5756__bF$buf1),
    .B(\datapath.registers.838[12] [8]),
    .C(\datapath.idinstr_15_bF$buf53 ),
    .Y(_6208_)
);

NAND2X1 _16855_ (
    .A(_6207_),
    .B(_6208_),
    .Y(_6209_)
);

NAND3X1 _16856_ (
    .A(\datapath.idinstr_17_bF$buf10 ),
    .B(_6206_),
    .C(_6209_),
    .Y(_6210_)
);

AOI21X1 _16857_ (
    .A(_6203_),
    .B(_6210_),
    .C(_5760__bF$buf3),
    .Y(_6211_)
);

INVX1 _16858_ (
    .A(\datapath.registers.838[1] [8]),
    .Y(_6212_)
);

AOI21X1 _16859_ (
    .A(\datapath.registers.838[5] [8]),
    .B(\datapath.idinstr_17_bF$buf9 ),
    .C(_5762__bF$buf6),
    .Y(_6213_)
);

OAI21X1 _16860_ (
    .A(_6212_),
    .B(\datapath.idinstr_17_bF$buf8 ),
    .C(_6213_),
    .Y(_6214_)
);

INVX1 _16861_ (
    .A(\datapath.registers.838[0] [8]),
    .Y(_6215_)
);

AOI21X1 _16862_ (
    .A(\datapath.registers.838[4] [8]),
    .B(\datapath.idinstr_17_bF$buf7 ),
    .C(\datapath.idinstr_15_bF$buf52 ),
    .Y(_6216_)
);

OAI21X1 _16863_ (
    .A(_6215_),
    .B(\datapath.idinstr_17_bF$buf6 ),
    .C(_6216_),
    .Y(_6217_)
);

NAND3X1 _16864_ (
    .A(_5756__bF$buf0),
    .B(_6217_),
    .C(_6214_),
    .Y(_6218_)
);

AOI21X1 _16865_ (
    .A(\datapath.registers.838[7] [8]),
    .B(\datapath.idinstr_17_bF$buf5 ),
    .C(_5762__bF$buf5),
    .Y(_6219_)
);

OAI21X1 _16866_ (
    .A(_5519_),
    .B(\datapath.idinstr_17_bF$buf4 ),
    .C(_6219_),
    .Y(_6220_)
);

INVX1 _16867_ (
    .A(\datapath.registers.838[2] [8]),
    .Y(_6221_)
);

AOI21X1 _16868_ (
    .A(\datapath.registers.838[6] [8]),
    .B(\datapath.idinstr_17_bF$buf3 ),
    .C(\datapath.idinstr_15_bF$buf51 ),
    .Y(_6222_)
);

OAI21X1 _16869_ (
    .A(_6221_),
    .B(\datapath.idinstr_17_bF$buf2 ),
    .C(_6222_),
    .Y(_6223_)
);

NAND3X1 _16870_ (
    .A(\datapath.idinstr_16_bF$buf51 ),
    .B(_6223_),
    .C(_6220_),
    .Y(_6224_)
);

AOI21X1 _16871_ (
    .A(_6218_),
    .B(_6224_),
    .C(\datapath.idinstr_18_bF$buf1 ),
    .Y(_6225_)
);

OAI21X1 _16872_ (
    .A(_6225_),
    .B(_6211_),
    .C(_5789__bF$buf1),
    .Y(_6226_)
);

AOI22X1 _16873_ (
    .A(_5755__bF$buf1),
    .B(_5759__bF$buf1),
    .C(_6226_),
    .D(_6196_),
    .Y(\datapath.registers.rega_data [8])
);

NAND2X1 _16874_ (
    .A(\datapath.idinstr_15_bF$buf50 ),
    .B(\datapath.registers.838[27] [9]),
    .Y(_6227_)
);

NAND2X1 _16875_ (
    .A(\datapath.registers.838[26] [9]),
    .B(_5762__bF$buf4),
    .Y(_6228_)
);

NAND3X1 _16876_ (
    .A(\datapath.idinstr_16_bF$buf50 ),
    .B(_6227_),
    .C(_6228_),
    .Y(_6229_)
);

NAND2X1 _16877_ (
    .A(\datapath.idinstr_15_bF$buf49 ),
    .B(\datapath.registers.838[25] [9]),
    .Y(_6230_)
);

AOI21X1 _16878_ (
    .A(_5762__bF$buf3),
    .B(\datapath.registers.838[24] [9]),
    .C(\datapath.idinstr_16_bF$buf49 ),
    .Y(_6231_)
);

NAND2X1 _16879_ (
    .A(_6230_),
    .B(_6231_),
    .Y(_6232_)
);

NAND3X1 _16880_ (
    .A(_5757__bF$buf6),
    .B(_6229_),
    .C(_6232_),
    .Y(_6233_)
);

NAND2X1 _16881_ (
    .A(\datapath.registers.838[31] [9]),
    .B(\datapath.idinstr_15_bF$buf48 ),
    .Y(_6234_)
);

AOI21X1 _16882_ (
    .A(_5762__bF$buf2),
    .B(\datapath.registers.838[30] [9]),
    .C(_5756__bF$buf9),
    .Y(_6235_)
);

NAND2X1 _16883_ (
    .A(_6234_),
    .B(_6235_),
    .Y(_6236_)
);

INVX1 _16884_ (
    .A(\datapath.registers.838[28] [9]),
    .Y(_6237_)
);

AOI21X1 _16885_ (
    .A(\datapath.idinstr_15_bF$buf47 ),
    .B(\datapath.registers.838[29] [9]),
    .C(\datapath.idinstr_16_bF$buf48 ),
    .Y(_6238_)
);

OAI21X1 _16886_ (
    .A(\datapath.idinstr_15_bF$buf46 ),
    .B(_6237_),
    .C(_6238_),
    .Y(_6239_)
);

NAND3X1 _16887_ (
    .A(\datapath.idinstr_17_bF$buf1 ),
    .B(_6239_),
    .C(_6236_),
    .Y(_6240_)
);

AOI21X1 _16888_ (
    .A(_6233_),
    .B(_6240_),
    .C(_5760__bF$buf2),
    .Y(_6241_)
);

MUX2X1 _16889_ (
    .A(\datapath.registers.838[18] [9]),
    .B(\datapath.registers.838[16] [9]),
    .S(\datapath.idinstr_16_bF$buf47 ),
    .Y(_6242_)
);

NAND2X1 _16890_ (
    .A(_5762__bF$buf1),
    .B(_6242_),
    .Y(_6243_)
);

MUX2X1 _16891_ (
    .A(\datapath.registers.838[19] [9]),
    .B(\datapath.registers.838[17] [9]),
    .S(\datapath.idinstr_16_bF$buf46 ),
    .Y(_6244_)
);

NAND2X1 _16892_ (
    .A(\datapath.idinstr_15_bF$buf45 ),
    .B(_6244_),
    .Y(_6245_)
);

NAND3X1 _16893_ (
    .A(_5757__bF$buf5),
    .B(_6243_),
    .C(_6245_),
    .Y(_6246_)
);

MUX2X1 _16894_ (
    .A(\datapath.registers.838[22] [9]),
    .B(\datapath.registers.838[20] [9]),
    .S(\datapath.idinstr_16_bF$buf45 ),
    .Y(_6247_)
);

NAND2X1 _16895_ (
    .A(_5762__bF$buf0),
    .B(_6247_),
    .Y(_6248_)
);

MUX2X1 _16896_ (
    .A(\datapath.registers.838[23] [9]),
    .B(\datapath.registers.838[21] [9]),
    .S(\datapath.idinstr_16_bF$buf44 ),
    .Y(_6249_)
);

NAND2X1 _16897_ (
    .A(\datapath.idinstr_15_bF$buf44 ),
    .B(_6249_),
    .Y(_6250_)
);

NAND3X1 _16898_ (
    .A(\datapath.idinstr_17_bF$buf0 ),
    .B(_6248_),
    .C(_6250_),
    .Y(_6251_)
);

AOI21X1 _16899_ (
    .A(_6246_),
    .B(_6251_),
    .C(\datapath.idinstr_18_bF$buf0 ),
    .Y(_6252_)
);

OAI21X1 _16900_ (
    .A(_6252_),
    .B(_6241_),
    .C(\datapath.idinstr_19_bF$buf3 ),
    .Y(_6253_)
);

AOI21X1 _16901_ (
    .A(\datapath.registers.838[13] [9]),
    .B(\datapath.idinstr_17_bF$buf15 ),
    .C(_5762__bF$buf47),
    .Y(_6254_)
);

OAI21X1 _16902_ (
    .A(_5277_),
    .B(\datapath.idinstr_17_bF$buf14 ),
    .C(_6254_),
    .Y(_6255_)
);

INVX1 _16903_ (
    .A(\datapath.registers.838[8] [9]),
    .Y(_6256_)
);

AOI21X1 _16904_ (
    .A(\datapath.registers.838[12] [9]),
    .B(\datapath.idinstr_17_bF$buf13 ),
    .C(\datapath.idinstr_15_bF$buf43 ),
    .Y(_6257_)
);

OAI21X1 _16905_ (
    .A(_6256_),
    .B(\datapath.idinstr_17_bF$buf12 ),
    .C(_6257_),
    .Y(_6258_)
);

NAND3X1 _16906_ (
    .A(_5756__bF$buf8),
    .B(_6258_),
    .C(_6255_),
    .Y(_6259_)
);

INVX1 _16907_ (
    .A(\datapath.registers.838[11] [9]),
    .Y(_6260_)
);

AOI21X1 _16908_ (
    .A(\datapath.registers.838[15] [9]),
    .B(\datapath.idinstr_17_bF$buf11 ),
    .C(_5762__bF$buf46),
    .Y(_6261_)
);

OAI21X1 _16909_ (
    .A(_6260_),
    .B(\datapath.idinstr_17_bF$buf10 ),
    .C(_6261_),
    .Y(_6262_)
);

AOI21X1 _16910_ (
    .A(\datapath.registers.838[14] [9]),
    .B(\datapath.idinstr_17_bF$buf9 ),
    .C(\datapath.idinstr_15_bF$buf42 ),
    .Y(_6263_)
);

OAI21X1 _16911_ (
    .A(_5233_),
    .B(\datapath.idinstr_17_bF$buf8 ),
    .C(_6263_),
    .Y(_6264_)
);

NAND3X1 _16912_ (
    .A(\datapath.idinstr_16_bF$buf43 ),
    .B(_6264_),
    .C(_6262_),
    .Y(_6265_)
);

AOI21X1 _16913_ (
    .A(_6259_),
    .B(_6265_),
    .C(_5760__bF$buf1),
    .Y(_6266_)
);

MUX2X1 _16914_ (
    .A(\datapath.registers.838[1] [9]),
    .B(\datapath.registers.838[0] [9]),
    .S(\datapath.idinstr_15_bF$buf41 ),
    .Y(_6267_)
);

NOR2X1 _16915_ (
    .A(\datapath.registers.838[3] [9]),
    .B(_5762__bF$buf45),
    .Y(_6268_)
);

OAI21X1 _16916_ (
    .A(\datapath.registers.838[2] [9]),
    .B(\datapath.idinstr_15_bF$buf40 ),
    .C(\datapath.idinstr_16_bF$buf42 ),
    .Y(_6269_)
);

OAI22X1 _16917_ (
    .A(_6269_),
    .B(_6268_),
    .C(\datapath.idinstr_16_bF$buf41 ),
    .D(_6267_),
    .Y(_6270_)
);

NAND2X1 _16918_ (
    .A(_5757__bF$buf4),
    .B(_6270_),
    .Y(_6271_)
);

MUX2X1 _16919_ (
    .A(\datapath.registers.838[5] [9]),
    .B(\datapath.registers.838[4] [9]),
    .S(\datapath.idinstr_15_bF$buf39 ),
    .Y(_6272_)
);

NOR2X1 _16920_ (
    .A(\datapath.registers.838[7] [9]),
    .B(_5762__bF$buf44),
    .Y(_6273_)
);

OAI21X1 _16921_ (
    .A(\datapath.registers.838[6] [9]),
    .B(\datapath.idinstr_15_bF$buf38 ),
    .C(\datapath.idinstr_16_bF$buf40 ),
    .Y(_6274_)
);

OAI22X1 _16922_ (
    .A(_6274_),
    .B(_6273_),
    .C(\datapath.idinstr_16_bF$buf39 ),
    .D(_6272_),
    .Y(_6275_)
);

NAND2X1 _16923_ (
    .A(\datapath.idinstr_17_bF$buf7 ),
    .B(_6275_),
    .Y(_6276_)
);

AOI21X1 _16924_ (
    .A(_6271_),
    .B(_6276_),
    .C(\datapath.idinstr_18_bF$buf6 ),
    .Y(_6277_)
);

OAI21X1 _16925_ (
    .A(_6266_),
    .B(_6277_),
    .C(_5789__bF$buf0),
    .Y(_6278_)
);

AOI22X1 _16926_ (
    .A(_5755__bF$buf0),
    .B(_5759__bF$buf0),
    .C(_6253_),
    .D(_6278_),
    .Y(\datapath.registers.rega_data [9])
);

NAND2X1 _16927_ (
    .A(\datapath.registers.838[11] [10]),
    .B(\datapath.idinstr_16_bF$buf38 ),
    .Y(_6279_)
);

NAND2X1 _16928_ (
    .A(\datapath.registers.838[9] [10]),
    .B(_5756__bF$buf7),
    .Y(_6280_)
);

NAND3X1 _16929_ (
    .A(\datapath.idinstr_15_bF$buf37 ),
    .B(_6279_),
    .C(_6280_),
    .Y(_6281_)
);

NAND2X1 _16930_ (
    .A(\datapath.registers.838[10] [10]),
    .B(\datapath.idinstr_16_bF$buf37 ),
    .Y(_6282_)
);

AOI21X1 _16931_ (
    .A(_5756__bF$buf6),
    .B(\datapath.registers.838[8] [10]),
    .C(\datapath.idinstr_15_bF$buf36 ),
    .Y(_6283_)
);

NAND2X1 _16932_ (
    .A(_6282_),
    .B(_6283_),
    .Y(_6284_)
);

NAND3X1 _16933_ (
    .A(_5757__bF$buf3),
    .B(_6281_),
    .C(_6284_),
    .Y(_6285_)
);

NAND2X1 _16934_ (
    .A(\datapath.registers.838[15] [10]),
    .B(\datapath.idinstr_16_bF$buf36 ),
    .Y(_6286_)
);

NAND2X1 _16935_ (
    .A(\datapath.registers.838[13] [10]),
    .B(_5756__bF$buf5),
    .Y(_6287_)
);

NAND3X1 _16936_ (
    .A(\datapath.idinstr_15_bF$buf35 ),
    .B(_6286_),
    .C(_6287_),
    .Y(_6288_)
);

NAND2X1 _16937_ (
    .A(\datapath.registers.838[14] [10]),
    .B(\datapath.idinstr_16_bF$buf35 ),
    .Y(_6289_)
);

AOI21X1 _16938_ (
    .A(_5756__bF$buf4),
    .B(\datapath.registers.838[12] [10]),
    .C(\datapath.idinstr_15_bF$buf34 ),
    .Y(_6290_)
);

NAND2X1 _16939_ (
    .A(_6289_),
    .B(_6290_),
    .Y(_6291_)
);

NAND3X1 _16940_ (
    .A(\datapath.idinstr_17_bF$buf6 ),
    .B(_6288_),
    .C(_6291_),
    .Y(_6292_)
);

AOI21X1 _16941_ (
    .A(_6285_),
    .B(_6292_),
    .C(_5760__bF$buf0),
    .Y(_6293_)
);

INVX1 _16942_ (
    .A(\datapath.registers.838[1] [10]),
    .Y(_6294_)
);

AOI21X1 _16943_ (
    .A(\datapath.registers.838[5] [10]),
    .B(\datapath.idinstr_17_bF$buf5 ),
    .C(_5762__bF$buf43),
    .Y(_6295_)
);

OAI21X1 _16944_ (
    .A(_6294_),
    .B(\datapath.idinstr_17_bF$buf4 ),
    .C(_6295_),
    .Y(_6296_)
);

INVX1 _16945_ (
    .A(\datapath.registers.838[0] [10]),
    .Y(_6297_)
);

AOI21X1 _16946_ (
    .A(\datapath.registers.838[4] [10]),
    .B(\datapath.idinstr_17_bF$buf3 ),
    .C(\datapath.idinstr_15_bF$buf33 ),
    .Y(_6298_)
);

OAI21X1 _16947_ (
    .A(_6297_),
    .B(\datapath.idinstr_17_bF$buf2 ),
    .C(_6298_),
    .Y(_6299_)
);

NAND3X1 _16948_ (
    .A(_5756__bF$buf3),
    .B(_6299_),
    .C(_6296_),
    .Y(_6300_)
);

AOI21X1 _16949_ (
    .A(\datapath.registers.838[7] [10]),
    .B(\datapath.idinstr_17_bF$buf1 ),
    .C(_5762__bF$buf42),
    .Y(_6301_)
);

OAI21X1 _16950_ (
    .A(_5523_),
    .B(\datapath.idinstr_17_bF$buf0 ),
    .C(_6301_),
    .Y(_6302_)
);

INVX1 _16951_ (
    .A(\datapath.registers.838[2] [10]),
    .Y(_6303_)
);

AOI21X1 _16952_ (
    .A(\datapath.registers.838[6] [10]),
    .B(\datapath.idinstr_17_bF$buf15 ),
    .C(\datapath.idinstr_15_bF$buf32 ),
    .Y(_6304_)
);

OAI21X1 _16953_ (
    .A(_6303_),
    .B(\datapath.idinstr_17_bF$buf14 ),
    .C(_6304_),
    .Y(_6305_)
);

NAND3X1 _16954_ (
    .A(\datapath.idinstr_16_bF$buf34 ),
    .B(_6305_),
    .C(_6302_),
    .Y(_6306_)
);

AOI21X1 _16955_ (
    .A(_6300_),
    .B(_6306_),
    .C(\datapath.idinstr_18_bF$buf5 ),
    .Y(_6307_)
);

OAI21X1 _16956_ (
    .A(_6307_),
    .B(_6293_),
    .C(_5789__bF$buf4),
    .Y(_6308_)
);

INVX1 _16957_ (
    .A(\datapath.registers.838[19] [10]),
    .Y(_6309_)
);

AOI21X1 _16958_ (
    .A(\datapath.registers.838[23] [10]),
    .B(\datapath.idinstr_17_bF$buf13 ),
    .C(_5762__bF$buf41),
    .Y(_6310_)
);

OAI21X1 _16959_ (
    .A(_6309_),
    .B(\datapath.idinstr_17_bF$buf12 ),
    .C(_6310_),
    .Y(_6311_)
);

NAND2X1 _16960_ (
    .A(\datapath.registers.838[18] [10]),
    .B(_5757__bF$buf2),
    .Y(_6312_)
);

AOI21X1 _16961_ (
    .A(\datapath.registers.838[22] [10]),
    .B(\datapath.idinstr_17_bF$buf11 ),
    .C(\datapath.idinstr_15_bF$buf31 ),
    .Y(_6313_)
);

AOI21X1 _16962_ (
    .A(_6312_),
    .B(_6313_),
    .C(_5756__bF$buf2),
    .Y(_6314_)
);

AOI21X1 _16963_ (
    .A(\datapath.registers.838[21] [10]),
    .B(\datapath.idinstr_17_bF$buf10 ),
    .C(_5762__bF$buf40),
    .Y(_6315_)
);

OAI21X1 _16964_ (
    .A(_4985_),
    .B(\datapath.idinstr_17_bF$buf9 ),
    .C(_6315_),
    .Y(_6316_)
);

NAND2X1 _16965_ (
    .A(\datapath.registers.838[16] [10]),
    .B(_5757__bF$buf1),
    .Y(_6317_)
);

AOI21X1 _16966_ (
    .A(\datapath.registers.838[20] [10]),
    .B(\datapath.idinstr_17_bF$buf8 ),
    .C(\datapath.idinstr_15_bF$buf30 ),
    .Y(_6318_)
);

AOI21X1 _16967_ (
    .A(_6317_),
    .B(_6318_),
    .C(\datapath.idinstr_16_bF$buf33 ),
    .Y(_6319_)
);

AOI22X1 _16968_ (
    .A(_6314_),
    .B(_6311_),
    .C(_6316_),
    .D(_6319_),
    .Y(_6320_)
);

NOR2X1 _16969_ (
    .A(\datapath.registers.838[24] [10]),
    .B(\datapath.idinstr_15_bF$buf29 ),
    .Y(_6321_)
);

OAI21X1 _16970_ (
    .A(\datapath.registers.838[25] [10]),
    .B(_5762__bF$buf39),
    .C(_5756__bF$buf1),
    .Y(_6322_)
);

NOR2X1 _16971_ (
    .A(\datapath.registers.838[27] [10]),
    .B(_5762__bF$buf38),
    .Y(_6323_)
);

OAI21X1 _16972_ (
    .A(\datapath.idinstr_15_bF$buf28 ),
    .B(\datapath.registers.838[26] [10]),
    .C(\datapath.idinstr_16_bF$buf32 ),
    .Y(_6324_)
);

OAI22X1 _16973_ (
    .A(_6323_),
    .B(_6324_),
    .C(_6321_),
    .D(_6322_),
    .Y(_6325_)
);

NOR2X1 _16974_ (
    .A(\datapath.idinstr_17_bF$buf7 ),
    .B(_6325_),
    .Y(_6326_)
);

MUX2X1 _16975_ (
    .A(\datapath.registers.838[29] [10]),
    .B(\datapath.registers.838[28] [10]),
    .S(\datapath.idinstr_15_bF$buf27 ),
    .Y(_6327_)
);

NOR2X1 _16976_ (
    .A(\datapath.registers.838[31] [10]),
    .B(_5762__bF$buf37),
    .Y(_6328_)
);

OAI21X1 _16977_ (
    .A(\datapath.registers.838[30] [10]),
    .B(\datapath.idinstr_15_bF$buf26 ),
    .C(\datapath.idinstr_16_bF$buf31 ),
    .Y(_6329_)
);

OAI22X1 _16978_ (
    .A(_6329_),
    .B(_6328_),
    .C(\datapath.idinstr_16_bF$buf30 ),
    .D(_6327_),
    .Y(_6330_)
);

OAI21X1 _16979_ (
    .A(_5757__bF$buf0),
    .B(_6330_),
    .C(\datapath.idinstr_18_bF$buf4 ),
    .Y(_6331_)
);

OAI22X1 _16980_ (
    .A(\datapath.idinstr_18_bF$buf3 ),
    .B(_6320_),
    .C(_6326_),
    .D(_6331_),
    .Y(_6332_)
);

NAND2X1 _16981_ (
    .A(\datapath.idinstr_19_bF$buf2 ),
    .B(_6332_),
    .Y(_6333_)
);

AOI22X1 _16982_ (
    .A(_5755__bF$buf4),
    .B(_5759__bF$buf4),
    .C(_6308_),
    .D(_6333_),
    .Y(\datapath.registers.rega_data [10])
);

NAND2X1 _16983_ (
    .A(\datapath.idinstr_15_bF$buf25 ),
    .B(\datapath.registers.838[27] [11]),
    .Y(_6334_)
);

NAND2X1 _16984_ (
    .A(\datapath.registers.838[26] [11]),
    .B(_5762__bF$buf36),
    .Y(_6335_)
);

NAND3X1 _16985_ (
    .A(\datapath.idinstr_16_bF$buf29 ),
    .B(_6334_),
    .C(_6335_),
    .Y(_6336_)
);

NAND2X1 _16986_ (
    .A(\datapath.idinstr_15_bF$buf24 ),
    .B(\datapath.registers.838[25] [11]),
    .Y(_6337_)
);

AOI21X1 _16987_ (
    .A(_5762__bF$buf35),
    .B(\datapath.registers.838[24] [11]),
    .C(\datapath.idinstr_16_bF$buf28 ),
    .Y(_6338_)
);

NAND2X1 _16988_ (
    .A(_6337_),
    .B(_6338_),
    .Y(_6339_)
);

NAND3X1 _16989_ (
    .A(_5757__bF$buf10),
    .B(_6336_),
    .C(_6339_),
    .Y(_6340_)
);

NAND2X1 _16990_ (
    .A(\datapath.registers.838[31] [11]),
    .B(\datapath.idinstr_15_bF$buf23 ),
    .Y(_6341_)
);

AOI21X1 _16991_ (
    .A(_5762__bF$buf34),
    .B(\datapath.registers.838[30] [11]),
    .C(_5756__bF$buf0),
    .Y(_6342_)
);

NAND2X1 _16992_ (
    .A(_6341_),
    .B(_6342_),
    .Y(_6343_)
);

INVX1 _16993_ (
    .A(\datapath.registers.838[28] [11]),
    .Y(_6344_)
);

AOI21X1 _16994_ (
    .A(\datapath.idinstr_15_bF$buf22 ),
    .B(\datapath.registers.838[29] [11]),
    .C(\datapath.idinstr_16_bF$buf27 ),
    .Y(_6345_)
);

OAI21X1 _16995_ (
    .A(\datapath.idinstr_15_bF$buf21 ),
    .B(_6344_),
    .C(_6345_),
    .Y(_6346_)
);

NAND3X1 _16996_ (
    .A(\datapath.idinstr_17_bF$buf6 ),
    .B(_6346_),
    .C(_6343_),
    .Y(_6347_)
);

AOI21X1 _16997_ (
    .A(_6340_),
    .B(_6347_),
    .C(_5760__bF$buf7),
    .Y(_6348_)
);

MUX2X1 _16998_ (
    .A(\datapath.registers.838[18] [11]),
    .B(\datapath.registers.838[16] [11]),
    .S(\datapath.idinstr_16_bF$buf26 ),
    .Y(_6349_)
);

NAND2X1 _16999_ (
    .A(_5762__bF$buf33),
    .B(_6349_),
    .Y(_6350_)
);

MUX2X1 _17000_ (
    .A(\datapath.registers.838[19] [11]),
    .B(\datapath.registers.838[17] [11]),
    .S(\datapath.idinstr_16_bF$buf25 ),
    .Y(_6351_)
);

NAND2X1 _17001_ (
    .A(\datapath.idinstr_15_bF$buf20 ),
    .B(_6351_),
    .Y(_6352_)
);

NAND3X1 _17002_ (
    .A(_5757__bF$buf9),
    .B(_6350_),
    .C(_6352_),
    .Y(_6353_)
);

MUX2X1 _17003_ (
    .A(\datapath.registers.838[22] [11]),
    .B(\datapath.registers.838[20] [11]),
    .S(\datapath.idinstr_16_bF$buf24 ),
    .Y(_6354_)
);

NAND2X1 _17004_ (
    .A(_5762__bF$buf32),
    .B(_6354_),
    .Y(_6355_)
);

MUX2X1 _17005_ (
    .A(\datapath.registers.838[23] [11]),
    .B(\datapath.registers.838[21] [11]),
    .S(\datapath.idinstr_16_bF$buf23 ),
    .Y(_6356_)
);

NAND2X1 _17006_ (
    .A(\datapath.idinstr_15_bF$buf19 ),
    .B(_6356_),
    .Y(_6357_)
);

NAND3X1 _17007_ (
    .A(\datapath.idinstr_17_bF$buf5 ),
    .B(_6355_),
    .C(_6357_),
    .Y(_6358_)
);

AOI21X1 _17008_ (
    .A(_6353_),
    .B(_6358_),
    .C(\datapath.idinstr_18_bF$buf2 ),
    .Y(_6359_)
);

OAI21X1 _17009_ (
    .A(_6359_),
    .B(_6348_),
    .C(\datapath.idinstr_19_bF$buf1 ),
    .Y(_6360_)
);

MUX2X1 _17010_ (
    .A(\datapath.registers.838[9] [11]),
    .B(\datapath.registers.838[8] [11]),
    .S(\datapath.idinstr_15_bF$buf18 ),
    .Y(_6361_)
);

NOR2X1 _17011_ (
    .A(\datapath.registers.838[11] [11]),
    .B(_5762__bF$buf31),
    .Y(_6362_)
);

OAI21X1 _17012_ (
    .A(\datapath.registers.838[10] [11]),
    .B(\datapath.idinstr_15_bF$buf17 ),
    .C(\datapath.idinstr_16_bF$buf22 ),
    .Y(_6363_)
);

OAI22X1 _17013_ (
    .A(_6363_),
    .B(_6362_),
    .C(\datapath.idinstr_16_bF$buf21 ),
    .D(_6361_),
    .Y(_6364_)
);

INVX1 _17014_ (
    .A(\datapath.registers.838[15] [11]),
    .Y(_6365_)
);

AOI21X1 _17015_ (
    .A(_5762__bF$buf30),
    .B(\datapath.registers.838[14] [11]),
    .C(_5756__bF$buf9),
    .Y(_6366_)
);

OAI21X1 _17016_ (
    .A(_6365_),
    .B(_5762__bF$buf29),
    .C(_6366_),
    .Y(_6367_)
);

NAND2X1 _17017_ (
    .A(\datapath.registers.838[12] [11]),
    .B(_5762__bF$buf28),
    .Y(_6368_)
);

AOI21X1 _17018_ (
    .A(\datapath.registers.838[13] [11]),
    .B(\datapath.idinstr_15_bF$buf16 ),
    .C(\datapath.idinstr_16_bF$buf20 ),
    .Y(_6369_)
);

AOI21X1 _17019_ (
    .A(_6368_),
    .B(_6369_),
    .C(_5757__bF$buf8),
    .Y(_6370_)
);

AOI22X1 _17020_ (
    .A(_6367_),
    .B(_6370_),
    .C(_5757__bF$buf7),
    .D(_6364_),
    .Y(_6371_)
);

NOR2X1 _17021_ (
    .A(\datapath.registers.838[0] [11]),
    .B(\datapath.idinstr_15_bF$buf15 ),
    .Y(_6372_)
);

OAI21X1 _17022_ (
    .A(\datapath.registers.838[1] [11]),
    .B(_5762__bF$buf27),
    .C(_5756__bF$buf8),
    .Y(_6373_)
);

NOR2X1 _17023_ (
    .A(\datapath.registers.838[3] [11]),
    .B(_5762__bF$buf26),
    .Y(_6374_)
);

OAI21X1 _17024_ (
    .A(\datapath.registers.838[2] [11]),
    .B(\datapath.idinstr_15_bF$buf14 ),
    .C(\datapath.idinstr_16_bF$buf19 ),
    .Y(_6375_)
);

OAI22X1 _17025_ (
    .A(_6374_),
    .B(_6375_),
    .C(_6372_),
    .D(_6373_),
    .Y(_6376_)
);

NOR2X1 _17026_ (
    .A(\datapath.idinstr_17_bF$buf4 ),
    .B(_6376_),
    .Y(_6377_)
);

MUX2X1 _17027_ (
    .A(\datapath.registers.838[5] [11]),
    .B(\datapath.registers.838[4] [11]),
    .S(\datapath.idinstr_15_bF$buf13 ),
    .Y(_6378_)
);

NOR2X1 _17028_ (
    .A(\datapath.registers.838[7] [11]),
    .B(_5762__bF$buf25),
    .Y(_6379_)
);

OAI21X1 _17029_ (
    .A(\datapath.registers.838[6] [11]),
    .B(\datapath.idinstr_15_bF$buf12 ),
    .C(\datapath.idinstr_16_bF$buf18 ),
    .Y(_6380_)
);

OAI22X1 _17030_ (
    .A(_6380_),
    .B(_6379_),
    .C(\datapath.idinstr_16_bF$buf17 ),
    .D(_6378_),
    .Y(_6381_)
);

OAI21X1 _17031_ (
    .A(_5757__bF$buf6),
    .B(_6381_),
    .C(_5760__bF$buf6),
    .Y(_6382_)
);

OAI22X1 _17032_ (
    .A(_5760__bF$buf5),
    .B(_6371_),
    .C(_6377_),
    .D(_6382_),
    .Y(_6383_)
);

NAND2X1 _17033_ (
    .A(_5789__bF$buf3),
    .B(_6383_),
    .Y(_6384_)
);

AOI22X1 _17034_ (
    .A(_5755__bF$buf3),
    .B(_5759__bF$buf3),
    .C(_6360_),
    .D(_6384_),
    .Y(\datapath.registers.rega_data [11])
);

NAND2X1 _17035_ (
    .A(\datapath.idinstr_15_bF$buf11 ),
    .B(\datapath.registers.838[27] [12]),
    .Y(_6385_)
);

NAND2X1 _17036_ (
    .A(\datapath.registers.838[26] [12]),
    .B(_5762__bF$buf24),
    .Y(_6386_)
);

NAND3X1 _17037_ (
    .A(\datapath.idinstr_16_bF$buf16 ),
    .B(_6385_),
    .C(_6386_),
    .Y(_6387_)
);

NAND2X1 _17038_ (
    .A(\datapath.idinstr_15_bF$buf10 ),
    .B(\datapath.registers.838[25] [12]),
    .Y(_6388_)
);

AOI21X1 _17039_ (
    .A(_5762__bF$buf23),
    .B(\datapath.registers.838[24] [12]),
    .C(\datapath.idinstr_16_bF$buf15 ),
    .Y(_6389_)
);

NAND2X1 _17040_ (
    .A(_6388_),
    .B(_6389_),
    .Y(_6390_)
);

NAND3X1 _17041_ (
    .A(_5757__bF$buf5),
    .B(_6387_),
    .C(_6390_),
    .Y(_6391_)
);

NAND2X1 _17042_ (
    .A(\datapath.registers.838[31] [12]),
    .B(\datapath.idinstr_15_bF$buf9 ),
    .Y(_6392_)
);

AOI21X1 _17043_ (
    .A(_5762__bF$buf22),
    .B(\datapath.registers.838[30] [12]),
    .C(_5756__bF$buf7),
    .Y(_6393_)
);

NAND2X1 _17044_ (
    .A(_6392_),
    .B(_6393_),
    .Y(_6394_)
);

INVX1 _17045_ (
    .A(\datapath.registers.838[28] [12]),
    .Y(_6395_)
);

AOI21X1 _17046_ (
    .A(\datapath.idinstr_15_bF$buf8 ),
    .B(\datapath.registers.838[29] [12]),
    .C(\datapath.idinstr_16_bF$buf14 ),
    .Y(_6396_)
);

OAI21X1 _17047_ (
    .A(\datapath.idinstr_15_bF$buf7 ),
    .B(_6395_),
    .C(_6396_),
    .Y(_6397_)
);

NAND3X1 _17048_ (
    .A(\datapath.idinstr_17_bF$buf3 ),
    .B(_6397_),
    .C(_6394_),
    .Y(_6398_)
);

AOI21X1 _17049_ (
    .A(_6391_),
    .B(_6398_),
    .C(_5760__bF$buf4),
    .Y(_6399_)
);

MUX2X1 _17050_ (
    .A(\datapath.registers.838[17] [12]),
    .B(\datapath.registers.838[16] [12]),
    .S(\datapath.idinstr_15_bF$buf6 ),
    .Y(_6400_)
);

NOR2X1 _17051_ (
    .A(\datapath.registers.838[19] [12]),
    .B(_5762__bF$buf21),
    .Y(_6401_)
);

OAI21X1 _17052_ (
    .A(\datapath.registers.838[18] [12]),
    .B(\datapath.idinstr_15_bF$buf5 ),
    .C(\datapath.idinstr_16_bF$buf13 ),
    .Y(_6402_)
);

OAI22X1 _17053_ (
    .A(_6402_),
    .B(_6401_),
    .C(\datapath.idinstr_16_bF$buf12 ),
    .D(_6400_),
    .Y(_6403_)
);

NAND2X1 _17054_ (
    .A(_5757__bF$buf4),
    .B(_6403_),
    .Y(_6404_)
);

MUX2X1 _17055_ (
    .A(\datapath.registers.838[21] [12]),
    .B(\datapath.registers.838[20] [12]),
    .S(\datapath.idinstr_15_bF$buf4 ),
    .Y(_6405_)
);

NOR2X1 _17056_ (
    .A(\datapath.registers.838[23] [12]),
    .B(_5762__bF$buf20),
    .Y(_6406_)
);

OAI21X1 _17057_ (
    .A(\datapath.registers.838[22] [12]),
    .B(\datapath.idinstr_15_bF$buf3 ),
    .C(\datapath.idinstr_16_bF$buf11 ),
    .Y(_6407_)
);

OAI22X1 _17058_ (
    .A(_6407_),
    .B(_6406_),
    .C(\datapath.idinstr_16_bF$buf10 ),
    .D(_6405_),
    .Y(_6408_)
);

NAND2X1 _17059_ (
    .A(\datapath.idinstr_17_bF$buf2 ),
    .B(_6408_),
    .Y(_6409_)
);

AOI21X1 _17060_ (
    .A(_6404_),
    .B(_6409_),
    .C(\datapath.idinstr_18_bF$buf1 ),
    .Y(_6410_)
);

OAI21X1 _17061_ (
    .A(_6399_),
    .B(_6410_),
    .C(\datapath.idinstr_19_bF$buf0 ),
    .Y(_6411_)
);

NAND2X1 _17062_ (
    .A(\datapath.registers.838[11] [12]),
    .B(\datapath.idinstr_16_bF$buf9 ),
    .Y(_6412_)
);

NAND2X1 _17063_ (
    .A(\datapath.registers.838[9] [12]),
    .B(_5756__bF$buf6),
    .Y(_6413_)
);

NAND3X1 _17064_ (
    .A(\datapath.idinstr_15_bF$buf2 ),
    .B(_6412_),
    .C(_6413_),
    .Y(_6414_)
);

NAND2X1 _17065_ (
    .A(\datapath.registers.838[10] [12]),
    .B(\datapath.idinstr_16_bF$buf8 ),
    .Y(_6415_)
);

AOI21X1 _17066_ (
    .A(_5756__bF$buf5),
    .B(\datapath.registers.838[8] [12]),
    .C(\datapath.idinstr_15_bF$buf1 ),
    .Y(_6416_)
);

NAND2X1 _17067_ (
    .A(_6415_),
    .B(_6416_),
    .Y(_6417_)
);

NAND3X1 _17068_ (
    .A(_5757__bF$buf3),
    .B(_6414_),
    .C(_6417_),
    .Y(_6418_)
);

NAND2X1 _17069_ (
    .A(\datapath.registers.838[15] [12]),
    .B(\datapath.idinstr_16_bF$buf7 ),
    .Y(_6419_)
);

NAND2X1 _17070_ (
    .A(\datapath.registers.838[13] [12]),
    .B(_5756__bF$buf4),
    .Y(_6420_)
);

NAND3X1 _17071_ (
    .A(\datapath.idinstr_15_bF$buf0 ),
    .B(_6419_),
    .C(_6420_),
    .Y(_6421_)
);

NAND2X1 _17072_ (
    .A(\datapath.registers.838[14] [12]),
    .B(\datapath.idinstr_16_bF$buf6 ),
    .Y(_6422_)
);

AOI21X1 _17073_ (
    .A(_5756__bF$buf3),
    .B(\datapath.registers.838[12] [12]),
    .C(\datapath.idinstr_15_bF$buf54 ),
    .Y(_6423_)
);

NAND2X1 _17074_ (
    .A(_6422_),
    .B(_6423_),
    .Y(_6424_)
);

NAND3X1 _17075_ (
    .A(\datapath.idinstr_17_bF$buf1 ),
    .B(_6421_),
    .C(_6424_),
    .Y(_6425_)
);

AOI21X1 _17076_ (
    .A(_6418_),
    .B(_6425_),
    .C(_5760__bF$buf3),
    .Y(_6426_)
);

INVX1 _17077_ (
    .A(\datapath.registers.838[1] [12]),
    .Y(_6427_)
);

AOI21X1 _17078_ (
    .A(\datapath.registers.838[5] [12]),
    .B(\datapath.idinstr_17_bF$buf0 ),
    .C(_5762__bF$buf19),
    .Y(_6428_)
);

OAI21X1 _17079_ (
    .A(_6427_),
    .B(\datapath.idinstr_17_bF$buf15 ),
    .C(_6428_),
    .Y(_6429_)
);

INVX1 _17080_ (
    .A(\datapath.registers.838[0] [12]),
    .Y(_6430_)
);

AOI21X1 _17081_ (
    .A(\datapath.registers.838[4] [12]),
    .B(\datapath.idinstr_17_bF$buf14 ),
    .C(\datapath.idinstr_15_bF$buf53 ),
    .Y(_6431_)
);

OAI21X1 _17082_ (
    .A(_6430_),
    .B(\datapath.idinstr_17_bF$buf13 ),
    .C(_6431_),
    .Y(_6432_)
);

NAND3X1 _17083_ (
    .A(_5756__bF$buf2),
    .B(_6432_),
    .C(_6429_),
    .Y(_6433_)
);

AOI21X1 _17084_ (
    .A(\datapath.registers.838[7] [12]),
    .B(\datapath.idinstr_17_bF$buf12 ),
    .C(_5762__bF$buf18),
    .Y(_6434_)
);

OAI21X1 _17085_ (
    .A(_5526_),
    .B(\datapath.idinstr_17_bF$buf11 ),
    .C(_6434_),
    .Y(_6435_)
);

INVX1 _17086_ (
    .A(\datapath.registers.838[2] [12]),
    .Y(_6436_)
);

AOI21X1 _17087_ (
    .A(\datapath.registers.838[6] [12]),
    .B(\datapath.idinstr_17_bF$buf10 ),
    .C(\datapath.idinstr_15_bF$buf52 ),
    .Y(_6437_)
);

OAI21X1 _17088_ (
    .A(_6436_),
    .B(\datapath.idinstr_17_bF$buf9 ),
    .C(_6437_),
    .Y(_6438_)
);

NAND3X1 _17089_ (
    .A(\datapath.idinstr_16_bF$buf5 ),
    .B(_6438_),
    .C(_6435_),
    .Y(_6439_)
);

AOI21X1 _17090_ (
    .A(_6433_),
    .B(_6439_),
    .C(\datapath.idinstr_18_bF$buf0 ),
    .Y(_6440_)
);

OAI21X1 _17091_ (
    .A(_6440_),
    .B(_6426_),
    .C(_5789__bF$buf2),
    .Y(_6441_)
);

AOI22X1 _17092_ (
    .A(_5755__bF$buf2),
    .B(_5759__bF$buf2),
    .C(_6441_),
    .D(_6411_),
    .Y(\datapath.registers.rega_data [12])
);

NAND2X1 _17093_ (
    .A(\datapath.idinstr_15_bF$buf51 ),
    .B(\datapath.registers.838[27] [13]),
    .Y(_6442_)
);

NAND2X1 _17094_ (
    .A(\datapath.registers.838[26] [13]),
    .B(_5762__bF$buf17),
    .Y(_6443_)
);

NAND3X1 _17095_ (
    .A(\datapath.idinstr_16_bF$buf4 ),
    .B(_6442_),
    .C(_6443_),
    .Y(_6444_)
);

NAND2X1 _17096_ (
    .A(\datapath.idinstr_15_bF$buf50 ),
    .B(\datapath.registers.838[25] [13]),
    .Y(_6445_)
);

AOI21X1 _17097_ (
    .A(_5762__bF$buf16),
    .B(\datapath.registers.838[24] [13]),
    .C(\datapath.idinstr_16_bF$buf3 ),
    .Y(_6446_)
);

NAND2X1 _17098_ (
    .A(_6445_),
    .B(_6446_),
    .Y(_6447_)
);

NAND3X1 _17099_ (
    .A(_5757__bF$buf2),
    .B(_6444_),
    .C(_6447_),
    .Y(_6448_)
);

NAND2X1 _17100_ (
    .A(\datapath.registers.838[31] [13]),
    .B(\datapath.idinstr_15_bF$buf49 ),
    .Y(_6449_)
);

AOI21X1 _17101_ (
    .A(_5762__bF$buf15),
    .B(\datapath.registers.838[30] [13]),
    .C(_5756__bF$buf1),
    .Y(_6450_)
);

NAND2X1 _17102_ (
    .A(_6449_),
    .B(_6450_),
    .Y(_6451_)
);

INVX1 _17103_ (
    .A(\datapath.registers.838[28] [13]),
    .Y(_6452_)
);

AOI21X1 _17104_ (
    .A(\datapath.idinstr_15_bF$buf48 ),
    .B(\datapath.registers.838[29] [13]),
    .C(\datapath.idinstr_16_bF$buf2 ),
    .Y(_6453_)
);

OAI21X1 _17105_ (
    .A(\datapath.idinstr_15_bF$buf47 ),
    .B(_6452_),
    .C(_6453_),
    .Y(_6454_)
);

NAND3X1 _17106_ (
    .A(\datapath.idinstr_17_bF$buf8 ),
    .B(_6454_),
    .C(_6451_),
    .Y(_6455_)
);

AOI21X1 _17107_ (
    .A(_6448_),
    .B(_6455_),
    .C(_5760__bF$buf2),
    .Y(_6456_)
);

MUX2X1 _17108_ (
    .A(\datapath.registers.838[18] [13]),
    .B(\datapath.registers.838[16] [13]),
    .S(\datapath.idinstr_16_bF$buf1 ),
    .Y(_6457_)
);

NAND2X1 _17109_ (
    .A(_5762__bF$buf14),
    .B(_6457_),
    .Y(_6458_)
);

MUX2X1 _17110_ (
    .A(\datapath.registers.838[19] [13]),
    .B(\datapath.registers.838[17] [13]),
    .S(\datapath.idinstr_16_bF$buf0 ),
    .Y(_6459_)
);

NAND2X1 _17111_ (
    .A(\datapath.idinstr_15_bF$buf46 ),
    .B(_6459_),
    .Y(_6460_)
);

NAND3X1 _17112_ (
    .A(_5757__bF$buf1),
    .B(_6458_),
    .C(_6460_),
    .Y(_6461_)
);

MUX2X1 _17113_ (
    .A(\datapath.registers.838[22] [13]),
    .B(\datapath.registers.838[20] [13]),
    .S(\datapath.idinstr_16_bF$buf51 ),
    .Y(_6462_)
);

NAND2X1 _17114_ (
    .A(_5762__bF$buf13),
    .B(_6462_),
    .Y(_6463_)
);

MUX2X1 _17115_ (
    .A(\datapath.registers.838[23] [13]),
    .B(\datapath.registers.838[21] [13]),
    .S(\datapath.idinstr_16_bF$buf50 ),
    .Y(_6464_)
);

NAND2X1 _17116_ (
    .A(\datapath.idinstr_15_bF$buf45 ),
    .B(_6464_),
    .Y(_6465_)
);

NAND3X1 _17117_ (
    .A(\datapath.idinstr_17_bF$buf7 ),
    .B(_6463_),
    .C(_6465_),
    .Y(_6466_)
);

AOI21X1 _17118_ (
    .A(_6461_),
    .B(_6466_),
    .C(\datapath.idinstr_18_bF$buf6 ),
    .Y(_6467_)
);

OAI21X1 _17119_ (
    .A(_6467_),
    .B(_6456_),
    .C(\datapath.idinstr_19_bF$buf5 ),
    .Y(_6468_)
);

MUX2X1 _17120_ (
    .A(\datapath.registers.838[9] [13]),
    .B(\datapath.registers.838[8] [13]),
    .S(\datapath.idinstr_15_bF$buf44 ),
    .Y(_6469_)
);

NOR2X1 _17121_ (
    .A(\datapath.registers.838[11] [13]),
    .B(_5762__bF$buf12),
    .Y(_6470_)
);

OAI21X1 _17122_ (
    .A(\datapath.registers.838[10] [13]),
    .B(\datapath.idinstr_15_bF$buf43 ),
    .C(\datapath.idinstr_16_bF$buf49 ),
    .Y(_6471_)
);

OAI22X1 _17123_ (
    .A(_6471_),
    .B(_6470_),
    .C(\datapath.idinstr_16_bF$buf48 ),
    .D(_6469_),
    .Y(_6472_)
);

INVX1 _17124_ (
    .A(\datapath.registers.838[15] [13]),
    .Y(_6473_)
);

AOI21X1 _17125_ (
    .A(_5762__bF$buf11),
    .B(\datapath.registers.838[14] [13]),
    .C(_5756__bF$buf0),
    .Y(_6474_)
);

OAI21X1 _17126_ (
    .A(_6473_),
    .B(_5762__bF$buf10),
    .C(_6474_),
    .Y(_6475_)
);

NAND2X1 _17127_ (
    .A(\datapath.registers.838[12] [13]),
    .B(_5762__bF$buf9),
    .Y(_6476_)
);

AOI21X1 _17128_ (
    .A(\datapath.registers.838[13] [13]),
    .B(\datapath.idinstr_15_bF$buf42 ),
    .C(\datapath.idinstr_16_bF$buf47 ),
    .Y(_6477_)
);

AOI21X1 _17129_ (
    .A(_6476_),
    .B(_6477_),
    .C(_5757__bF$buf0),
    .Y(_6478_)
);

AOI22X1 _17130_ (
    .A(_6475_),
    .B(_6478_),
    .C(_5757__bF$buf10),
    .D(_6472_),
    .Y(_6479_)
);

NOR2X1 _17131_ (
    .A(\datapath.registers.838[0] [13]),
    .B(\datapath.idinstr_15_bF$buf41 ),
    .Y(_6480_)
);

OAI21X1 _17132_ (
    .A(\datapath.registers.838[1] [13]),
    .B(_5762__bF$buf8),
    .C(_5756__bF$buf9),
    .Y(_6481_)
);

NOR2X1 _17133_ (
    .A(\datapath.registers.838[3] [13]),
    .B(_5762__bF$buf7),
    .Y(_6482_)
);

OAI21X1 _17134_ (
    .A(\datapath.registers.838[2] [13]),
    .B(\datapath.idinstr_15_bF$buf40 ),
    .C(\datapath.idinstr_16_bF$buf46 ),
    .Y(_6483_)
);

OAI22X1 _17135_ (
    .A(_6482_),
    .B(_6483_),
    .C(_6480_),
    .D(_6481_),
    .Y(_6484_)
);

NOR2X1 _17136_ (
    .A(\datapath.idinstr_17_bF$buf6 ),
    .B(_6484_),
    .Y(_6485_)
);

MUX2X1 _17137_ (
    .A(\datapath.registers.838[5] [13]),
    .B(\datapath.registers.838[4] [13]),
    .S(\datapath.idinstr_15_bF$buf39 ),
    .Y(_6486_)
);

NOR2X1 _17138_ (
    .A(\datapath.registers.838[7] [13]),
    .B(_5762__bF$buf6),
    .Y(_6487_)
);

OAI21X1 _17139_ (
    .A(\datapath.registers.838[6] [13]),
    .B(\datapath.idinstr_15_bF$buf38 ),
    .C(\datapath.idinstr_16_bF$buf45 ),
    .Y(_6488_)
);

OAI22X1 _17140_ (
    .A(_6488_),
    .B(_6487_),
    .C(\datapath.idinstr_16_bF$buf44 ),
    .D(_6486_),
    .Y(_6489_)
);

OAI21X1 _17141_ (
    .A(_5757__bF$buf9),
    .B(_6489_),
    .C(_5760__bF$buf1),
    .Y(_6490_)
);

OAI22X1 _17142_ (
    .A(_5760__bF$buf0),
    .B(_6479_),
    .C(_6485_),
    .D(_6490_),
    .Y(_6491_)
);

NAND2X1 _17143_ (
    .A(_5789__bF$buf1),
    .B(_6491_),
    .Y(_6492_)
);

AOI22X1 _17144_ (
    .A(_5755__bF$buf1),
    .B(_5759__bF$buf1),
    .C(_6468_),
    .D(_6492_),
    .Y(\datapath.registers.rega_data [13])
);

NAND2X1 _17145_ (
    .A(\datapath.idinstr_15_bF$buf37 ),
    .B(\datapath.registers.838[27] [14]),
    .Y(_6493_)
);

NAND2X1 _17146_ (
    .A(\datapath.registers.838[26] [14]),
    .B(_5762__bF$buf5),
    .Y(_6494_)
);

NAND3X1 _17147_ (
    .A(\datapath.idinstr_16_bF$buf43 ),
    .B(_6493_),
    .C(_6494_),
    .Y(_6495_)
);

NAND2X1 _17148_ (
    .A(\datapath.idinstr_15_bF$buf36 ),
    .B(\datapath.registers.838[25] [14]),
    .Y(_6496_)
);

AOI21X1 _17149_ (
    .A(_5762__bF$buf4),
    .B(\datapath.registers.838[24] [14]),
    .C(\datapath.idinstr_16_bF$buf42 ),
    .Y(_6497_)
);

NAND2X1 _17150_ (
    .A(_6496_),
    .B(_6497_),
    .Y(_6498_)
);

NAND3X1 _17151_ (
    .A(_5757__bF$buf8),
    .B(_6495_),
    .C(_6498_),
    .Y(_6499_)
);

NAND2X1 _17152_ (
    .A(\datapath.registers.838[31] [14]),
    .B(\datapath.idinstr_15_bF$buf35 ),
    .Y(_6500_)
);

AOI21X1 _17153_ (
    .A(_5762__bF$buf3),
    .B(\datapath.registers.838[30] [14]),
    .C(_5756__bF$buf8),
    .Y(_6501_)
);

NAND2X1 _17154_ (
    .A(_6500_),
    .B(_6501_),
    .Y(_6502_)
);

INVX1 _17155_ (
    .A(\datapath.registers.838[28] [14]),
    .Y(_6503_)
);

AOI21X1 _17156_ (
    .A(\datapath.idinstr_15_bF$buf34 ),
    .B(\datapath.registers.838[29] [14]),
    .C(\datapath.idinstr_16_bF$buf41 ),
    .Y(_6504_)
);

OAI21X1 _17157_ (
    .A(\datapath.idinstr_15_bF$buf33 ),
    .B(_6503_),
    .C(_6504_),
    .Y(_6505_)
);

NAND3X1 _17158_ (
    .A(\datapath.idinstr_17_bF$buf5 ),
    .B(_6505_),
    .C(_6502_),
    .Y(_6506_)
);

AOI21X1 _17159_ (
    .A(_6499_),
    .B(_6506_),
    .C(_5760__bF$buf7),
    .Y(_6507_)
);

MUX2X1 _17160_ (
    .A(\datapath.registers.838[18] [14]),
    .B(\datapath.registers.838[16] [14]),
    .S(\datapath.idinstr_16_bF$buf40 ),
    .Y(_6508_)
);

NAND2X1 _17161_ (
    .A(_5762__bF$buf2),
    .B(_6508_),
    .Y(_6509_)
);

MUX2X1 _17162_ (
    .A(\datapath.registers.838[19] [14]),
    .B(\datapath.registers.838[17] [14]),
    .S(\datapath.idinstr_16_bF$buf39 ),
    .Y(_6510_)
);

NAND2X1 _17163_ (
    .A(\datapath.idinstr_15_bF$buf32 ),
    .B(_6510_),
    .Y(_6511_)
);

NAND3X1 _17164_ (
    .A(_5757__bF$buf7),
    .B(_6509_),
    .C(_6511_),
    .Y(_6512_)
);

MUX2X1 _17165_ (
    .A(\datapath.registers.838[22] [14]),
    .B(\datapath.registers.838[20] [14]),
    .S(\datapath.idinstr_16_bF$buf38 ),
    .Y(_6513_)
);

NAND2X1 _17166_ (
    .A(_5762__bF$buf1),
    .B(_6513_),
    .Y(_6514_)
);

MUX2X1 _17167_ (
    .A(\datapath.registers.838[23] [14]),
    .B(\datapath.registers.838[21] [14]),
    .S(\datapath.idinstr_16_bF$buf37 ),
    .Y(_6515_)
);

NAND2X1 _17168_ (
    .A(\datapath.idinstr_15_bF$buf31 ),
    .B(_6515_),
    .Y(_6516_)
);

NAND3X1 _17169_ (
    .A(\datapath.idinstr_17_bF$buf4 ),
    .B(_6514_),
    .C(_6516_),
    .Y(_6517_)
);

AOI21X1 _17170_ (
    .A(_6512_),
    .B(_6517_),
    .C(\datapath.idinstr_18_bF$buf5 ),
    .Y(_6518_)
);

OAI21X1 _17171_ (
    .A(_6518_),
    .B(_6507_),
    .C(\datapath.idinstr_19_bF$buf4 ),
    .Y(_6519_)
);

MUX2X1 _17172_ (
    .A(\datapath.registers.838[9] [14]),
    .B(\datapath.registers.838[8] [14]),
    .S(\datapath.idinstr_15_bF$buf30 ),
    .Y(_6520_)
);

NOR2X1 _17173_ (
    .A(\datapath.registers.838[11] [14]),
    .B(_5762__bF$buf0),
    .Y(_6521_)
);

OAI21X1 _17174_ (
    .A(\datapath.registers.838[10] [14]),
    .B(\datapath.idinstr_15_bF$buf29 ),
    .C(\datapath.idinstr_16_bF$buf36 ),
    .Y(_6522_)
);

OAI22X1 _17175_ (
    .A(_6522_),
    .B(_6521_),
    .C(\datapath.idinstr_16_bF$buf35 ),
    .D(_6520_),
    .Y(_6523_)
);

INVX1 _17176_ (
    .A(\datapath.registers.838[15] [14]),
    .Y(_6524_)
);

AOI21X1 _17177_ (
    .A(_5762__bF$buf47),
    .B(\datapath.registers.838[14] [14]),
    .C(_5756__bF$buf7),
    .Y(_6525_)
);

OAI21X1 _17178_ (
    .A(_6524_),
    .B(_5762__bF$buf46),
    .C(_6525_),
    .Y(_6526_)
);

NAND2X1 _17179_ (
    .A(\datapath.registers.838[12] [14]),
    .B(_5762__bF$buf45),
    .Y(_6527_)
);

AOI21X1 _17180_ (
    .A(\datapath.registers.838[13] [14]),
    .B(\datapath.idinstr_15_bF$buf28 ),
    .C(\datapath.idinstr_16_bF$buf34 ),
    .Y(_6528_)
);

AOI21X1 _17181_ (
    .A(_6527_),
    .B(_6528_),
    .C(_5757__bF$buf6),
    .Y(_6529_)
);

AOI22X1 _17182_ (
    .A(_6526_),
    .B(_6529_),
    .C(_5757__bF$buf5),
    .D(_6523_),
    .Y(_6530_)
);

NOR2X1 _17183_ (
    .A(\datapath.registers.838[0] [14]),
    .B(\datapath.idinstr_15_bF$buf27 ),
    .Y(_6531_)
);

OAI21X1 _17184_ (
    .A(\datapath.registers.838[1] [14]),
    .B(_5762__bF$buf44),
    .C(_5756__bF$buf6),
    .Y(_6532_)
);

NOR2X1 _17185_ (
    .A(\datapath.registers.838[3] [14]),
    .B(_5762__bF$buf43),
    .Y(_6533_)
);

OAI21X1 _17186_ (
    .A(\datapath.registers.838[2] [14]),
    .B(\datapath.idinstr_15_bF$buf26 ),
    .C(\datapath.idinstr_16_bF$buf33 ),
    .Y(_6534_)
);

OAI22X1 _17187_ (
    .A(_6533_),
    .B(_6534_),
    .C(_6531_),
    .D(_6532_),
    .Y(_6535_)
);

NOR2X1 _17188_ (
    .A(\datapath.idinstr_17_bF$buf3 ),
    .B(_6535_),
    .Y(_6536_)
);

MUX2X1 _17189_ (
    .A(\datapath.registers.838[5] [14]),
    .B(\datapath.registers.838[4] [14]),
    .S(\datapath.idinstr_15_bF$buf25 ),
    .Y(_6537_)
);

NOR2X1 _17190_ (
    .A(\datapath.registers.838[7] [14]),
    .B(_5762__bF$buf42),
    .Y(_6538_)
);

OAI21X1 _17191_ (
    .A(\datapath.registers.838[6] [14]),
    .B(\datapath.idinstr_15_bF$buf24 ),
    .C(\datapath.idinstr_16_bF$buf32 ),
    .Y(_6539_)
);

OAI22X1 _17192_ (
    .A(_6539_),
    .B(_6538_),
    .C(\datapath.idinstr_16_bF$buf31 ),
    .D(_6537_),
    .Y(_6540_)
);

OAI21X1 _17193_ (
    .A(_5757__bF$buf4),
    .B(_6540_),
    .C(_5760__bF$buf6),
    .Y(_6541_)
);

OAI22X1 _17194_ (
    .A(_5760__bF$buf5),
    .B(_6530_),
    .C(_6536_),
    .D(_6541_),
    .Y(_6542_)
);

NAND2X1 _17195_ (
    .A(_5789__bF$buf0),
    .B(_6542_),
    .Y(_6543_)
);

AOI22X1 _17196_ (
    .A(_5755__bF$buf0),
    .B(_5759__bF$buf0),
    .C(_6519_),
    .D(_6543_),
    .Y(\datapath.registers.rega_data [14])
);

MUX2X1 _17197_ (
    .A(\datapath.registers.838[9] [15]),
    .B(\datapath.registers.838[8] [15]),
    .S(\datapath.idinstr_15_bF$buf23 ),
    .Y(_6544_)
);

NOR2X1 _17198_ (
    .A(\datapath.registers.838[11] [15]),
    .B(_5762__bF$buf41),
    .Y(_6545_)
);

OAI21X1 _17199_ (
    .A(\datapath.registers.838[10] [15]),
    .B(\datapath.idinstr_15_bF$buf22 ),
    .C(\datapath.idinstr_16_bF$buf30 ),
    .Y(_6546_)
);

OAI22X1 _17200_ (
    .A(_6546_),
    .B(_6545_),
    .C(\datapath.idinstr_16_bF$buf29 ),
    .D(_6544_),
    .Y(_6547_)
);

INVX1 _17201_ (
    .A(\datapath.registers.838[15] [15]),
    .Y(_6548_)
);

AOI21X1 _17202_ (
    .A(_5762__bF$buf40),
    .B(\datapath.registers.838[14] [15]),
    .C(_5756__bF$buf5),
    .Y(_6549_)
);

OAI21X1 _17203_ (
    .A(_6548_),
    .B(_5762__bF$buf39),
    .C(_6549_),
    .Y(_6550_)
);

NAND2X1 _17204_ (
    .A(\datapath.registers.838[12] [15]),
    .B(_5762__bF$buf38),
    .Y(_6551_)
);

AOI21X1 _17205_ (
    .A(\datapath.registers.838[13] [15]),
    .B(\datapath.idinstr_15_bF$buf21 ),
    .C(\datapath.idinstr_16_bF$buf28 ),
    .Y(_6552_)
);

AOI21X1 _17206_ (
    .A(_6551_),
    .B(_6552_),
    .C(_5757__bF$buf3),
    .Y(_6553_)
);

AOI22X1 _17207_ (
    .A(_6550_),
    .B(_6553_),
    .C(_5757__bF$buf2),
    .D(_6547_),
    .Y(_6554_)
);

NOR2X1 _17208_ (
    .A(\datapath.registers.838[0] [15]),
    .B(\datapath.idinstr_15_bF$buf20 ),
    .Y(_6555_)
);

OAI21X1 _17209_ (
    .A(\datapath.registers.838[1] [15]),
    .B(_5762__bF$buf37),
    .C(_5756__bF$buf4),
    .Y(_6556_)
);

NOR2X1 _17210_ (
    .A(\datapath.registers.838[3] [15]),
    .B(_5762__bF$buf36),
    .Y(_6557_)
);

OAI21X1 _17211_ (
    .A(\datapath.registers.838[2] [15]),
    .B(\datapath.idinstr_15_bF$buf19 ),
    .C(\datapath.idinstr_16_bF$buf27 ),
    .Y(_6558_)
);

OAI22X1 _17212_ (
    .A(_6557_),
    .B(_6558_),
    .C(_6555_),
    .D(_6556_),
    .Y(_6559_)
);

NOR2X1 _17213_ (
    .A(\datapath.idinstr_17_bF$buf2 ),
    .B(_6559_),
    .Y(_6560_)
);

MUX2X1 _17214_ (
    .A(\datapath.registers.838[5] [15]),
    .B(\datapath.registers.838[4] [15]),
    .S(\datapath.idinstr_15_bF$buf18 ),
    .Y(_6561_)
);

NOR2X1 _17215_ (
    .A(\datapath.registers.838[7] [15]),
    .B(_5762__bF$buf35),
    .Y(_6562_)
);

OAI21X1 _17216_ (
    .A(\datapath.registers.838[6] [15]),
    .B(\datapath.idinstr_15_bF$buf17 ),
    .C(\datapath.idinstr_16_bF$buf26 ),
    .Y(_6563_)
);

OAI22X1 _17217_ (
    .A(_6563_),
    .B(_6562_),
    .C(\datapath.idinstr_16_bF$buf25 ),
    .D(_6561_),
    .Y(_6564_)
);

OAI21X1 _17218_ (
    .A(_5757__bF$buf1),
    .B(_6564_),
    .C(_5760__bF$buf4),
    .Y(_6565_)
);

OAI22X1 _17219_ (
    .A(_5760__bF$buf3),
    .B(_6554_),
    .C(_6560_),
    .D(_6565_),
    .Y(_6566_)
);

NAND2X1 _17220_ (
    .A(_5789__bF$buf4),
    .B(_6566_),
    .Y(_6567_)
);

INVX1 _17221_ (
    .A(\datapath.registers.838[27] [15]),
    .Y(_6568_)
);

AOI21X1 _17222_ (
    .A(\datapath.registers.838[31] [15]),
    .B(\datapath.idinstr_17_bF$buf1 ),
    .C(_5762__bF$buf34),
    .Y(_6569_)
);

OAI21X1 _17223_ (
    .A(\datapath.idinstr_17_bF$buf0 ),
    .B(_6568_),
    .C(_6569_),
    .Y(_6570_)
);

INVX1 _17224_ (
    .A(\datapath.registers.838[26] [15]),
    .Y(_6571_)
);

AOI21X1 _17225_ (
    .A(\datapath.registers.838[30] [15]),
    .B(\datapath.idinstr_17_bF$buf15 ),
    .C(\datapath.idinstr_15_bF$buf16 ),
    .Y(_6572_)
);

OAI21X1 _17226_ (
    .A(\datapath.idinstr_17_bF$buf14 ),
    .B(_6571_),
    .C(_6572_),
    .Y(_6573_)
);

NAND3X1 _17227_ (
    .A(\datapath.idinstr_16_bF$buf24 ),
    .B(_6573_),
    .C(_6570_),
    .Y(_6574_)
);

INVX1 _17228_ (
    .A(\datapath.registers.838[25] [15]),
    .Y(_6575_)
);

AOI21X1 _17229_ (
    .A(\datapath.idinstr_17_bF$buf13 ),
    .B(\datapath.registers.838[29] [15]),
    .C(_5762__bF$buf33),
    .Y(_6576_)
);

OAI21X1 _17230_ (
    .A(\datapath.idinstr_17_bF$buf12 ),
    .B(_6575_),
    .C(_6576_),
    .Y(_6577_)
);

INVX1 _17231_ (
    .A(\datapath.registers.838[24] [15]),
    .Y(_6578_)
);

AOI21X1 _17232_ (
    .A(\datapath.idinstr_17_bF$buf11 ),
    .B(\datapath.registers.838[28] [15]),
    .C(\datapath.idinstr_15_bF$buf15 ),
    .Y(_6579_)
);

OAI21X1 _17233_ (
    .A(_6578_),
    .B(\datapath.idinstr_17_bF$buf10 ),
    .C(_6579_),
    .Y(_6580_)
);

NAND3X1 _17234_ (
    .A(_5756__bF$buf3),
    .B(_6580_),
    .C(_6577_),
    .Y(_6581_)
);

AOI21X1 _17235_ (
    .A(_6574_),
    .B(_6581_),
    .C(_5760__bF$buf2),
    .Y(_6582_)
);

MUX2X1 _17236_ (
    .A(\datapath.registers.838[18] [15]),
    .B(\datapath.registers.838[16] [15]),
    .S(\datapath.idinstr_16_bF$buf23 ),
    .Y(_6583_)
);

NAND2X1 _17237_ (
    .A(_5762__bF$buf32),
    .B(_6583_),
    .Y(_6584_)
);

MUX2X1 _17238_ (
    .A(\datapath.registers.838[19] [15]),
    .B(\datapath.registers.838[17] [15]),
    .S(\datapath.idinstr_16_bF$buf22 ),
    .Y(_6585_)
);

NAND2X1 _17239_ (
    .A(\datapath.idinstr_15_bF$buf14 ),
    .B(_6585_),
    .Y(_6586_)
);

NAND3X1 _17240_ (
    .A(_5757__bF$buf0),
    .B(_6584_),
    .C(_6586_),
    .Y(_6587_)
);

MUX2X1 _17241_ (
    .A(\datapath.registers.838[22] [15]),
    .B(\datapath.registers.838[20] [15]),
    .S(\datapath.idinstr_16_bF$buf21 ),
    .Y(_6588_)
);

NAND2X1 _17242_ (
    .A(_5762__bF$buf31),
    .B(_6588_),
    .Y(_6589_)
);

MUX2X1 _17243_ (
    .A(\datapath.registers.838[23] [15]),
    .B(\datapath.registers.838[21] [15]),
    .S(\datapath.idinstr_16_bF$buf20 ),
    .Y(_6590_)
);

NAND2X1 _17244_ (
    .A(\datapath.idinstr_15_bF$buf13 ),
    .B(_6590_),
    .Y(_6591_)
);

NAND3X1 _17245_ (
    .A(\datapath.idinstr_17_bF$buf9 ),
    .B(_6589_),
    .C(_6591_),
    .Y(_6592_)
);

AOI21X1 _17246_ (
    .A(_6587_),
    .B(_6592_),
    .C(\datapath.idinstr_18_bF$buf4 ),
    .Y(_6593_)
);

OAI21X1 _17247_ (
    .A(_6582_),
    .B(_6593_),
    .C(\datapath.idinstr_19_bF$buf3 ),
    .Y(_6594_)
);

AOI22X1 _17248_ (
    .A(_5755__bF$buf4),
    .B(_5759__bF$buf4),
    .C(_6594_),
    .D(_6567_),
    .Y(\datapath.registers.rega_data [15])
);

MUX2X1 _17249_ (
    .A(\datapath.registers.838[9] [16]),
    .B(\datapath.registers.838[8] [16]),
    .S(\datapath.idinstr_15_bF$buf12 ),
    .Y(_6595_)
);

NOR2X1 _17250_ (
    .A(\datapath.registers.838[11] [16]),
    .B(_5762__bF$buf30),
    .Y(_6596_)
);

OAI21X1 _17251_ (
    .A(\datapath.registers.838[10] [16]),
    .B(\datapath.idinstr_15_bF$buf11 ),
    .C(\datapath.idinstr_16_bF$buf19 ),
    .Y(_6597_)
);

OAI22X1 _17252_ (
    .A(_6597_),
    .B(_6596_),
    .C(\datapath.idinstr_16_bF$buf18 ),
    .D(_6595_),
    .Y(_6598_)
);

INVX1 _17253_ (
    .A(\datapath.registers.838[15] [16]),
    .Y(_6599_)
);

AOI21X1 _17254_ (
    .A(_5762__bF$buf29),
    .B(\datapath.registers.838[14] [16]),
    .C(_5756__bF$buf2),
    .Y(_6600_)
);

OAI21X1 _17255_ (
    .A(_6599_),
    .B(_5762__bF$buf28),
    .C(_6600_),
    .Y(_6601_)
);

NAND2X1 _17256_ (
    .A(\datapath.registers.838[12] [16]),
    .B(_5762__bF$buf27),
    .Y(_6602_)
);

AOI21X1 _17257_ (
    .A(\datapath.registers.838[13] [16]),
    .B(\datapath.idinstr_15_bF$buf10 ),
    .C(\datapath.idinstr_16_bF$buf17 ),
    .Y(_6603_)
);

AOI21X1 _17258_ (
    .A(_6602_),
    .B(_6603_),
    .C(_5757__bF$buf10),
    .Y(_6604_)
);

AOI22X1 _17259_ (
    .A(_6601_),
    .B(_6604_),
    .C(_5757__bF$buf9),
    .D(_6598_),
    .Y(_6605_)
);

NOR2X1 _17260_ (
    .A(\datapath.registers.838[0] [16]),
    .B(\datapath.idinstr_15_bF$buf9 ),
    .Y(_6606_)
);

OAI21X1 _17261_ (
    .A(\datapath.registers.838[1] [16]),
    .B(_5762__bF$buf26),
    .C(_5756__bF$buf1),
    .Y(_6607_)
);

NOR2X1 _17262_ (
    .A(\datapath.registers.838[3] [16]),
    .B(_5762__bF$buf25),
    .Y(_6608_)
);

OAI21X1 _17263_ (
    .A(\datapath.registers.838[2] [16]),
    .B(\datapath.idinstr_15_bF$buf8 ),
    .C(\datapath.idinstr_16_bF$buf16 ),
    .Y(_6609_)
);

OAI22X1 _17264_ (
    .A(_6608_),
    .B(_6609_),
    .C(_6606_),
    .D(_6607_),
    .Y(_6610_)
);

NOR2X1 _17265_ (
    .A(\datapath.idinstr_17_bF$buf8 ),
    .B(_6610_),
    .Y(_6611_)
);

MUX2X1 _17266_ (
    .A(\datapath.registers.838[5] [16]),
    .B(\datapath.registers.838[4] [16]),
    .S(\datapath.idinstr_15_bF$buf7 ),
    .Y(_6612_)
);

NOR2X1 _17267_ (
    .A(\datapath.registers.838[7] [16]),
    .B(_5762__bF$buf24),
    .Y(_6613_)
);

OAI21X1 _17268_ (
    .A(\datapath.registers.838[6] [16]),
    .B(\datapath.idinstr_15_bF$buf6 ),
    .C(\datapath.idinstr_16_bF$buf15 ),
    .Y(_6614_)
);

OAI22X1 _17269_ (
    .A(_6614_),
    .B(_6613_),
    .C(\datapath.idinstr_16_bF$buf14 ),
    .D(_6612_),
    .Y(_6615_)
);

OAI21X1 _17270_ (
    .A(_5757__bF$buf8),
    .B(_6615_),
    .C(_5760__bF$buf1),
    .Y(_6616_)
);

OAI22X1 _17271_ (
    .A(_5760__bF$buf0),
    .B(_6605_),
    .C(_6611_),
    .D(_6616_),
    .Y(_6617_)
);

NAND2X1 _17272_ (
    .A(_5789__bF$buf3),
    .B(_6617_),
    .Y(_6618_)
);

INVX1 _17273_ (
    .A(\datapath.registers.838[27] [16]),
    .Y(_6619_)
);

AOI21X1 _17274_ (
    .A(\datapath.registers.838[31] [16]),
    .B(\datapath.idinstr_17_bF$buf7 ),
    .C(_5762__bF$buf23),
    .Y(_6620_)
);

OAI21X1 _17275_ (
    .A(\datapath.idinstr_17_bF$buf6 ),
    .B(_6619_),
    .C(_6620_),
    .Y(_6621_)
);

INVX1 _17276_ (
    .A(\datapath.registers.838[26] [16]),
    .Y(_6622_)
);

AOI21X1 _17277_ (
    .A(\datapath.registers.838[30] [16]),
    .B(\datapath.idinstr_17_bF$buf5 ),
    .C(\datapath.idinstr_15_bF$buf5 ),
    .Y(_6623_)
);

OAI21X1 _17278_ (
    .A(\datapath.idinstr_17_bF$buf4 ),
    .B(_6622_),
    .C(_6623_),
    .Y(_6624_)
);

NAND3X1 _17279_ (
    .A(\datapath.idinstr_16_bF$buf13 ),
    .B(_6624_),
    .C(_6621_),
    .Y(_6625_)
);

INVX1 _17280_ (
    .A(\datapath.registers.838[25] [16]),
    .Y(_6626_)
);

AOI21X1 _17281_ (
    .A(\datapath.idinstr_17_bF$buf3 ),
    .B(\datapath.registers.838[29] [16]),
    .C(_5762__bF$buf22),
    .Y(_6627_)
);

OAI21X1 _17282_ (
    .A(\datapath.idinstr_17_bF$buf2 ),
    .B(_6626_),
    .C(_6627_),
    .Y(_6628_)
);

INVX1 _17283_ (
    .A(\datapath.registers.838[24] [16]),
    .Y(_6629_)
);

AOI21X1 _17284_ (
    .A(\datapath.idinstr_17_bF$buf1 ),
    .B(\datapath.registers.838[28] [16]),
    .C(\datapath.idinstr_15_bF$buf4 ),
    .Y(_6630_)
);

OAI21X1 _17285_ (
    .A(_6629_),
    .B(\datapath.idinstr_17_bF$buf0 ),
    .C(_6630_),
    .Y(_6631_)
);

NAND3X1 _17286_ (
    .A(_5756__bF$buf0),
    .B(_6631_),
    .C(_6628_),
    .Y(_6632_)
);

AOI21X1 _17287_ (
    .A(_6625_),
    .B(_6632_),
    .C(_5760__bF$buf7),
    .Y(_6633_)
);

MUX2X1 _17288_ (
    .A(\datapath.registers.838[18] [16]),
    .B(\datapath.registers.838[16] [16]),
    .S(\datapath.idinstr_16_bF$buf12 ),
    .Y(_6634_)
);

NAND2X1 _17289_ (
    .A(_5762__bF$buf21),
    .B(_6634_),
    .Y(_6635_)
);

MUX2X1 _17290_ (
    .A(\datapath.registers.838[19] [16]),
    .B(\datapath.registers.838[17] [16]),
    .S(\datapath.idinstr_16_bF$buf11 ),
    .Y(_6636_)
);

NAND2X1 _17291_ (
    .A(\datapath.idinstr_15_bF$buf3 ),
    .B(_6636_),
    .Y(_6637_)
);

NAND3X1 _17292_ (
    .A(_5757__bF$buf7),
    .B(_6635_),
    .C(_6637_),
    .Y(_6638_)
);

MUX2X1 _17293_ (
    .A(\datapath.registers.838[22] [16]),
    .B(\datapath.registers.838[20] [16]),
    .S(\datapath.idinstr_16_bF$buf10 ),
    .Y(_6639_)
);

NAND2X1 _17294_ (
    .A(_5762__bF$buf20),
    .B(_6639_),
    .Y(_6640_)
);

MUX2X1 _17295_ (
    .A(\datapath.registers.838[23] [16]),
    .B(\datapath.registers.838[21] [16]),
    .S(\datapath.idinstr_16_bF$buf9 ),
    .Y(_6641_)
);

NAND2X1 _17296_ (
    .A(\datapath.idinstr_15_bF$buf2 ),
    .B(_6641_),
    .Y(_6642_)
);

NAND3X1 _17297_ (
    .A(\datapath.idinstr_17_bF$buf15 ),
    .B(_6640_),
    .C(_6642_),
    .Y(_6643_)
);

AOI21X1 _17298_ (
    .A(_6638_),
    .B(_6643_),
    .C(\datapath.idinstr_18_bF$buf3 ),
    .Y(_6644_)
);

OAI21X1 _17299_ (
    .A(_6633_),
    .B(_6644_),
    .C(\datapath.idinstr_19_bF$buf2 ),
    .Y(_6645_)
);

AOI22X1 _17300_ (
    .A(_5755__bF$buf3),
    .B(_5759__bF$buf3),
    .C(_6645_),
    .D(_6618_),
    .Y(\datapath.registers.rega_data [16])
);

NAND2X1 _17301_ (
    .A(\datapath.idinstr_15_bF$buf1 ),
    .B(\datapath.registers.838[27] [17]),
    .Y(_6646_)
);

NAND2X1 _17302_ (
    .A(\datapath.registers.838[26] [17]),
    .B(_5762__bF$buf19),
    .Y(_6647_)
);

NAND3X1 _17303_ (
    .A(\datapath.idinstr_16_bF$buf8 ),
    .B(_6646_),
    .C(_6647_),
    .Y(_6648_)
);

NAND2X1 _17304_ (
    .A(\datapath.idinstr_15_bF$buf0 ),
    .B(\datapath.registers.838[25] [17]),
    .Y(_6649_)
);

AOI21X1 _17305_ (
    .A(_5762__bF$buf18),
    .B(\datapath.registers.838[24] [17]),
    .C(\datapath.idinstr_16_bF$buf7 ),
    .Y(_6650_)
);

NAND2X1 _17306_ (
    .A(_6649_),
    .B(_6650_),
    .Y(_6651_)
);

NAND3X1 _17307_ (
    .A(_5757__bF$buf6),
    .B(_6648_),
    .C(_6651_),
    .Y(_6652_)
);

NAND2X1 _17308_ (
    .A(\datapath.registers.838[31] [17]),
    .B(\datapath.idinstr_15_bF$buf54 ),
    .Y(_6653_)
);

AOI21X1 _17309_ (
    .A(_5762__bF$buf17),
    .B(\datapath.registers.838[30] [17]),
    .C(_5756__bF$buf9),
    .Y(_6654_)
);

NAND2X1 _17310_ (
    .A(_6653_),
    .B(_6654_),
    .Y(_6655_)
);

INVX1 _17311_ (
    .A(\datapath.registers.838[28] [17]),
    .Y(_6656_)
);

AOI21X1 _17312_ (
    .A(\datapath.idinstr_15_bF$buf53 ),
    .B(\datapath.registers.838[29] [17]),
    .C(\datapath.idinstr_16_bF$buf6 ),
    .Y(_6657_)
);

OAI21X1 _17313_ (
    .A(\datapath.idinstr_15_bF$buf52 ),
    .B(_6656_),
    .C(_6657_),
    .Y(_6658_)
);

NAND3X1 _17314_ (
    .A(\datapath.idinstr_17_bF$buf14 ),
    .B(_6658_),
    .C(_6655_),
    .Y(_6659_)
);

AOI21X1 _17315_ (
    .A(_6652_),
    .B(_6659_),
    .C(_5760__bF$buf6),
    .Y(_6660_)
);

MUX2X1 _17316_ (
    .A(\datapath.registers.838[18] [17]),
    .B(\datapath.registers.838[16] [17]),
    .S(\datapath.idinstr_16_bF$buf5 ),
    .Y(_6661_)
);

NAND2X1 _17317_ (
    .A(_5762__bF$buf16),
    .B(_6661_),
    .Y(_6662_)
);

MUX2X1 _17318_ (
    .A(\datapath.registers.838[19] [17]),
    .B(\datapath.registers.838[17] [17]),
    .S(\datapath.idinstr_16_bF$buf4 ),
    .Y(_6663_)
);

NAND2X1 _17319_ (
    .A(\datapath.idinstr_15_bF$buf51 ),
    .B(_6663_),
    .Y(_6664_)
);

NAND3X1 _17320_ (
    .A(_5757__bF$buf5),
    .B(_6662_),
    .C(_6664_),
    .Y(_6665_)
);

MUX2X1 _17321_ (
    .A(\datapath.registers.838[22] [17]),
    .B(\datapath.registers.838[20] [17]),
    .S(\datapath.idinstr_16_bF$buf3 ),
    .Y(_6666_)
);

NAND2X1 _17322_ (
    .A(_5762__bF$buf15),
    .B(_6666_),
    .Y(_6667_)
);

MUX2X1 _17323_ (
    .A(\datapath.registers.838[23] [17]),
    .B(\datapath.registers.838[21] [17]),
    .S(\datapath.idinstr_16_bF$buf2 ),
    .Y(_6668_)
);

NAND2X1 _17324_ (
    .A(\datapath.idinstr_15_bF$buf50 ),
    .B(_6668_),
    .Y(_6669_)
);

NAND3X1 _17325_ (
    .A(\datapath.idinstr_17_bF$buf13 ),
    .B(_6667_),
    .C(_6669_),
    .Y(_6670_)
);

AOI21X1 _17326_ (
    .A(_6665_),
    .B(_6670_),
    .C(\datapath.idinstr_18_bF$buf2 ),
    .Y(_6671_)
);

OAI21X1 _17327_ (
    .A(_6671_),
    .B(_6660_),
    .C(\datapath.idinstr_19_bF$buf1 ),
    .Y(_6672_)
);

MUX2X1 _17328_ (
    .A(\datapath.registers.838[9] [17]),
    .B(\datapath.registers.838[8] [17]),
    .S(\datapath.idinstr_15_bF$buf49 ),
    .Y(_6673_)
);

NOR2X1 _17329_ (
    .A(\datapath.registers.838[11] [17]),
    .B(_5762__bF$buf14),
    .Y(_6674_)
);

OAI21X1 _17330_ (
    .A(\datapath.registers.838[10] [17]),
    .B(\datapath.idinstr_15_bF$buf48 ),
    .C(\datapath.idinstr_16_bF$buf1 ),
    .Y(_6675_)
);

OAI22X1 _17331_ (
    .A(_6675_),
    .B(_6674_),
    .C(\datapath.idinstr_16_bF$buf0 ),
    .D(_6673_),
    .Y(_6676_)
);

INVX1 _17332_ (
    .A(\datapath.registers.838[15] [17]),
    .Y(_6677_)
);

AOI21X1 _17333_ (
    .A(_5762__bF$buf13),
    .B(\datapath.registers.838[14] [17]),
    .C(_5756__bF$buf8),
    .Y(_6678_)
);

OAI21X1 _17334_ (
    .A(_6677_),
    .B(_5762__bF$buf12),
    .C(_6678_),
    .Y(_6679_)
);

NAND2X1 _17335_ (
    .A(\datapath.registers.838[12] [17]),
    .B(_5762__bF$buf11),
    .Y(_6680_)
);

AOI21X1 _17336_ (
    .A(\datapath.registers.838[13] [17]),
    .B(\datapath.idinstr_15_bF$buf47 ),
    .C(\datapath.idinstr_16_bF$buf51 ),
    .Y(_6681_)
);

AOI21X1 _17337_ (
    .A(_6680_),
    .B(_6681_),
    .C(_5757__bF$buf4),
    .Y(_6682_)
);

AOI22X1 _17338_ (
    .A(_6679_),
    .B(_6682_),
    .C(_5757__bF$buf3),
    .D(_6676_),
    .Y(_6683_)
);

NOR2X1 _17339_ (
    .A(\datapath.registers.838[0] [17]),
    .B(\datapath.idinstr_15_bF$buf46 ),
    .Y(_6684_)
);

OAI21X1 _17340_ (
    .A(\datapath.registers.838[1] [17]),
    .B(_5762__bF$buf10),
    .C(_5756__bF$buf7),
    .Y(_6685_)
);

NOR2X1 _17341_ (
    .A(\datapath.registers.838[3] [17]),
    .B(_5762__bF$buf9),
    .Y(_6686_)
);

OAI21X1 _17342_ (
    .A(\datapath.registers.838[2] [17]),
    .B(\datapath.idinstr_15_bF$buf45 ),
    .C(\datapath.idinstr_16_bF$buf50 ),
    .Y(_6687_)
);

OAI22X1 _17343_ (
    .A(_6686_),
    .B(_6687_),
    .C(_6684_),
    .D(_6685_),
    .Y(_6688_)
);

NOR2X1 _17344_ (
    .A(\datapath.idinstr_17_bF$buf12 ),
    .B(_6688_),
    .Y(_6689_)
);

MUX2X1 _17345_ (
    .A(\datapath.registers.838[5] [17]),
    .B(\datapath.registers.838[4] [17]),
    .S(\datapath.idinstr_15_bF$buf44 ),
    .Y(_6690_)
);

NOR2X1 _17346_ (
    .A(\datapath.registers.838[7] [17]),
    .B(_5762__bF$buf8),
    .Y(_6691_)
);

OAI21X1 _17347_ (
    .A(\datapath.registers.838[6] [17]),
    .B(\datapath.idinstr_15_bF$buf43 ),
    .C(\datapath.idinstr_16_bF$buf49 ),
    .Y(_6692_)
);

OAI22X1 _17348_ (
    .A(_6692_),
    .B(_6691_),
    .C(\datapath.idinstr_16_bF$buf48 ),
    .D(_6690_),
    .Y(_6693_)
);

OAI21X1 _17349_ (
    .A(_5757__bF$buf2),
    .B(_6693_),
    .C(_5760__bF$buf5),
    .Y(_6694_)
);

OAI22X1 _17350_ (
    .A(_5760__bF$buf4),
    .B(_6683_),
    .C(_6689_),
    .D(_6694_),
    .Y(_6695_)
);

NAND2X1 _17351_ (
    .A(_5789__bF$buf2),
    .B(_6695_),
    .Y(_6696_)
);

AOI22X1 _17352_ (
    .A(_5755__bF$buf2),
    .B(_5759__bF$buf2),
    .C(_6672_),
    .D(_6696_),
    .Y(\datapath.registers.rega_data [17])
);

NAND2X1 _17353_ (
    .A(\datapath.idinstr_15_bF$buf42 ),
    .B(\datapath.registers.838[27] [18]),
    .Y(_6697_)
);

NAND2X1 _17354_ (
    .A(\datapath.registers.838[26] [18]),
    .B(_5762__bF$buf7),
    .Y(_6698_)
);

NAND3X1 _17355_ (
    .A(\datapath.idinstr_16_bF$buf47 ),
    .B(_6697_),
    .C(_6698_),
    .Y(_6699_)
);

NAND2X1 _17356_ (
    .A(\datapath.idinstr_15_bF$buf41 ),
    .B(\datapath.registers.838[25] [18]),
    .Y(_6700_)
);

AOI21X1 _17357_ (
    .A(_5762__bF$buf6),
    .B(\datapath.registers.838[24] [18]),
    .C(\datapath.idinstr_16_bF$buf46 ),
    .Y(_6701_)
);

NAND2X1 _17358_ (
    .A(_6700_),
    .B(_6701_),
    .Y(_6702_)
);

NAND3X1 _17359_ (
    .A(_5757__bF$buf1),
    .B(_6699_),
    .C(_6702_),
    .Y(_6703_)
);

NAND2X1 _17360_ (
    .A(\datapath.registers.838[31] [18]),
    .B(\datapath.idinstr_15_bF$buf40 ),
    .Y(_6704_)
);

AOI21X1 _17361_ (
    .A(_5762__bF$buf5),
    .B(\datapath.registers.838[30] [18]),
    .C(_5756__bF$buf6),
    .Y(_6705_)
);

NAND2X1 _17362_ (
    .A(_6704_),
    .B(_6705_),
    .Y(_6706_)
);

INVX1 _17363_ (
    .A(\datapath.registers.838[28] [18]),
    .Y(_6707_)
);

AOI21X1 _17364_ (
    .A(\datapath.idinstr_15_bF$buf39 ),
    .B(\datapath.registers.838[29] [18]),
    .C(\datapath.idinstr_16_bF$buf45 ),
    .Y(_6708_)
);

OAI21X1 _17365_ (
    .A(\datapath.idinstr_15_bF$buf38 ),
    .B(_6707_),
    .C(_6708_),
    .Y(_6709_)
);

NAND3X1 _17366_ (
    .A(\datapath.idinstr_17_bF$buf11 ),
    .B(_6709_),
    .C(_6706_),
    .Y(_6710_)
);

AOI21X1 _17367_ (
    .A(_6703_),
    .B(_6710_),
    .C(_5760__bF$buf3),
    .Y(_6711_)
);

MUX2X1 _17368_ (
    .A(\datapath.registers.838[18] [18]),
    .B(\datapath.registers.838[16] [18]),
    .S(\datapath.idinstr_16_bF$buf44 ),
    .Y(_6712_)
);

NAND2X1 _17369_ (
    .A(_5762__bF$buf4),
    .B(_6712_),
    .Y(_6713_)
);

MUX2X1 _17370_ (
    .A(\datapath.registers.838[19] [18]),
    .B(\datapath.registers.838[17] [18]),
    .S(\datapath.idinstr_16_bF$buf43 ),
    .Y(_6714_)
);

NAND2X1 _17371_ (
    .A(\datapath.idinstr_15_bF$buf37 ),
    .B(_6714_),
    .Y(_6715_)
);

NAND3X1 _17372_ (
    .A(_5757__bF$buf0),
    .B(_6713_),
    .C(_6715_),
    .Y(_6716_)
);

MUX2X1 _17373_ (
    .A(\datapath.registers.838[22] [18]),
    .B(\datapath.registers.838[20] [18]),
    .S(\datapath.idinstr_16_bF$buf42 ),
    .Y(_6717_)
);

NAND2X1 _17374_ (
    .A(_5762__bF$buf3),
    .B(_6717_),
    .Y(_6718_)
);

MUX2X1 _17375_ (
    .A(\datapath.registers.838[23] [18]),
    .B(\datapath.registers.838[21] [18]),
    .S(\datapath.idinstr_16_bF$buf41 ),
    .Y(_6719_)
);

NAND2X1 _17376_ (
    .A(\datapath.idinstr_15_bF$buf36 ),
    .B(_6719_),
    .Y(_6720_)
);

NAND3X1 _17377_ (
    .A(\datapath.idinstr_17_bF$buf10 ),
    .B(_6718_),
    .C(_6720_),
    .Y(_6721_)
);

AOI21X1 _17378_ (
    .A(_6716_),
    .B(_6721_),
    .C(\datapath.idinstr_18_bF$buf1 ),
    .Y(_6722_)
);

OAI21X1 _17379_ (
    .A(_6722_),
    .B(_6711_),
    .C(\datapath.idinstr_19_bF$buf0 ),
    .Y(_6723_)
);

MUX2X1 _17380_ (
    .A(\datapath.registers.838[9] [18]),
    .B(\datapath.registers.838[8] [18]),
    .S(\datapath.idinstr_15_bF$buf35 ),
    .Y(_6724_)
);

NOR2X1 _17381_ (
    .A(\datapath.registers.838[11] [18]),
    .B(_5762__bF$buf2),
    .Y(_6725_)
);

OAI21X1 _17382_ (
    .A(\datapath.registers.838[10] [18]),
    .B(\datapath.idinstr_15_bF$buf34 ),
    .C(\datapath.idinstr_16_bF$buf40 ),
    .Y(_6726_)
);

OAI22X1 _17383_ (
    .A(_6726_),
    .B(_6725_),
    .C(\datapath.idinstr_16_bF$buf39 ),
    .D(_6724_),
    .Y(_6727_)
);

INVX1 _17384_ (
    .A(\datapath.registers.838[15] [18]),
    .Y(_6728_)
);

AOI21X1 _17385_ (
    .A(_5762__bF$buf1),
    .B(\datapath.registers.838[14] [18]),
    .C(_5756__bF$buf5),
    .Y(_6729_)
);

OAI21X1 _17386_ (
    .A(_6728_),
    .B(_5762__bF$buf0),
    .C(_6729_),
    .Y(_6730_)
);

NAND2X1 _17387_ (
    .A(\datapath.registers.838[12] [18]),
    .B(_5762__bF$buf47),
    .Y(_6731_)
);

AOI21X1 _17388_ (
    .A(\datapath.registers.838[13] [18]),
    .B(\datapath.idinstr_15_bF$buf33 ),
    .C(\datapath.idinstr_16_bF$buf38 ),
    .Y(_6732_)
);

AOI21X1 _17389_ (
    .A(_6731_),
    .B(_6732_),
    .C(_5757__bF$buf10),
    .Y(_6733_)
);

AOI22X1 _17390_ (
    .A(_6730_),
    .B(_6733_),
    .C(_5757__bF$buf9),
    .D(_6727_),
    .Y(_6734_)
);

NOR2X1 _17391_ (
    .A(\datapath.registers.838[0] [18]),
    .B(\datapath.idinstr_15_bF$buf32 ),
    .Y(_6735_)
);

OAI21X1 _17392_ (
    .A(\datapath.registers.838[1] [18]),
    .B(_5762__bF$buf46),
    .C(_5756__bF$buf4),
    .Y(_6736_)
);

NOR2X1 _17393_ (
    .A(\datapath.registers.838[3] [18]),
    .B(_5762__bF$buf45),
    .Y(_6737_)
);

OAI21X1 _17394_ (
    .A(\datapath.registers.838[2] [18]),
    .B(\datapath.idinstr_15_bF$buf31 ),
    .C(\datapath.idinstr_16_bF$buf37 ),
    .Y(_6738_)
);

OAI22X1 _17395_ (
    .A(_6737_),
    .B(_6738_),
    .C(_6735_),
    .D(_6736_),
    .Y(_6739_)
);

NOR2X1 _17396_ (
    .A(\datapath.idinstr_17_bF$buf9 ),
    .B(_6739_),
    .Y(_6740_)
);

MUX2X1 _17397_ (
    .A(\datapath.registers.838[5] [18]),
    .B(\datapath.registers.838[4] [18]),
    .S(\datapath.idinstr_15_bF$buf30 ),
    .Y(_6741_)
);

NOR2X1 _17398_ (
    .A(\datapath.registers.838[7] [18]),
    .B(_5762__bF$buf44),
    .Y(_6742_)
);

OAI21X1 _17399_ (
    .A(\datapath.registers.838[6] [18]),
    .B(\datapath.idinstr_15_bF$buf29 ),
    .C(\datapath.idinstr_16_bF$buf36 ),
    .Y(_6743_)
);

OAI22X1 _17400_ (
    .A(_6743_),
    .B(_6742_),
    .C(\datapath.idinstr_16_bF$buf35 ),
    .D(_6741_),
    .Y(_6744_)
);

OAI21X1 _17401_ (
    .A(_5757__bF$buf8),
    .B(_6744_),
    .C(_5760__bF$buf2),
    .Y(_6745_)
);

OAI22X1 _17402_ (
    .A(_5760__bF$buf1),
    .B(_6734_),
    .C(_6740_),
    .D(_6745_),
    .Y(_6746_)
);

NAND2X1 _17403_ (
    .A(_5789__bF$buf1),
    .B(_6746_),
    .Y(_6747_)
);

AOI22X1 _17404_ (
    .A(_5755__bF$buf1),
    .B(_5759__bF$buf1),
    .C(_6723_),
    .D(_6747_),
    .Y(\datapath.registers.rega_data [18])
);

NAND2X1 _17405_ (
    .A(\datapath.idinstr_15_bF$buf28 ),
    .B(\datapath.registers.838[27] [19]),
    .Y(_6748_)
);

NAND2X1 _17406_ (
    .A(\datapath.registers.838[26] [19]),
    .B(_5762__bF$buf43),
    .Y(_6749_)
);

NAND3X1 _17407_ (
    .A(\datapath.idinstr_16_bF$buf34 ),
    .B(_6748_),
    .C(_6749_),
    .Y(_6750_)
);

NAND2X1 _17408_ (
    .A(\datapath.idinstr_15_bF$buf27 ),
    .B(\datapath.registers.838[25] [19]),
    .Y(_6751_)
);

AOI21X1 _17409_ (
    .A(_5762__bF$buf42),
    .B(\datapath.registers.838[24] [19]),
    .C(\datapath.idinstr_16_bF$buf33 ),
    .Y(_6752_)
);

NAND2X1 _17410_ (
    .A(_6751_),
    .B(_6752_),
    .Y(_6753_)
);

NAND3X1 _17411_ (
    .A(_5757__bF$buf7),
    .B(_6750_),
    .C(_6753_),
    .Y(_6754_)
);

NAND2X1 _17412_ (
    .A(\datapath.registers.838[31] [19]),
    .B(\datapath.idinstr_15_bF$buf26 ),
    .Y(_6755_)
);

AOI21X1 _17413_ (
    .A(_5762__bF$buf41),
    .B(\datapath.registers.838[30] [19]),
    .C(_5756__bF$buf3),
    .Y(_6756_)
);

NAND2X1 _17414_ (
    .A(_6755_),
    .B(_6756_),
    .Y(_6757_)
);

INVX1 _17415_ (
    .A(\datapath.registers.838[28] [19]),
    .Y(_6758_)
);

AOI21X1 _17416_ (
    .A(\datapath.idinstr_15_bF$buf25 ),
    .B(\datapath.registers.838[29] [19]),
    .C(\datapath.idinstr_16_bF$buf32 ),
    .Y(_6759_)
);

OAI21X1 _17417_ (
    .A(\datapath.idinstr_15_bF$buf24 ),
    .B(_6758_),
    .C(_6759_),
    .Y(_6760_)
);

NAND3X1 _17418_ (
    .A(\datapath.idinstr_17_bF$buf8 ),
    .B(_6760_),
    .C(_6757_),
    .Y(_6761_)
);

AOI21X1 _17419_ (
    .A(_6754_),
    .B(_6761_),
    .C(_5760__bF$buf0),
    .Y(_6762_)
);

MUX2X1 _17420_ (
    .A(\datapath.registers.838[18] [19]),
    .B(\datapath.registers.838[16] [19]),
    .S(\datapath.idinstr_16_bF$buf31 ),
    .Y(_6763_)
);

NAND2X1 _17421_ (
    .A(_5762__bF$buf40),
    .B(_6763_),
    .Y(_6764_)
);

MUX2X1 _17422_ (
    .A(\datapath.registers.838[19] [19]),
    .B(\datapath.registers.838[17] [19]),
    .S(\datapath.idinstr_16_bF$buf30 ),
    .Y(_6765_)
);

NAND2X1 _17423_ (
    .A(\datapath.idinstr_15_bF$buf23 ),
    .B(_6765_),
    .Y(_6766_)
);

NAND3X1 _17424_ (
    .A(_5757__bF$buf6),
    .B(_6764_),
    .C(_6766_),
    .Y(_6767_)
);

MUX2X1 _17425_ (
    .A(\datapath.registers.838[22] [19]),
    .B(\datapath.registers.838[20] [19]),
    .S(\datapath.idinstr_16_bF$buf29 ),
    .Y(_6768_)
);

NAND2X1 _17426_ (
    .A(_5762__bF$buf39),
    .B(_6768_),
    .Y(_6769_)
);

MUX2X1 _17427_ (
    .A(\datapath.registers.838[23] [19]),
    .B(\datapath.registers.838[21] [19]),
    .S(\datapath.idinstr_16_bF$buf28 ),
    .Y(_6770_)
);

NAND2X1 _17428_ (
    .A(\datapath.idinstr_15_bF$buf22 ),
    .B(_6770_),
    .Y(_6771_)
);

NAND3X1 _17429_ (
    .A(\datapath.idinstr_17_bF$buf7 ),
    .B(_6769_),
    .C(_6771_),
    .Y(_6772_)
);

AOI21X1 _17430_ (
    .A(_6767_),
    .B(_6772_),
    .C(\datapath.idinstr_18_bF$buf0 ),
    .Y(_6773_)
);

OAI21X1 _17431_ (
    .A(_6773_),
    .B(_6762_),
    .C(\datapath.idinstr_19_bF$buf5 ),
    .Y(_6774_)
);

MUX2X1 _17432_ (
    .A(\datapath.registers.838[9] [19]),
    .B(\datapath.registers.838[8] [19]),
    .S(\datapath.idinstr_15_bF$buf21 ),
    .Y(_6775_)
);

NOR2X1 _17433_ (
    .A(\datapath.registers.838[11] [19]),
    .B(_5762__bF$buf38),
    .Y(_6776_)
);

OAI21X1 _17434_ (
    .A(\datapath.registers.838[10] [19]),
    .B(\datapath.idinstr_15_bF$buf20 ),
    .C(\datapath.idinstr_16_bF$buf27 ),
    .Y(_6777_)
);

OAI22X1 _17435_ (
    .A(_6777_),
    .B(_6776_),
    .C(\datapath.idinstr_16_bF$buf26 ),
    .D(_6775_),
    .Y(_6778_)
);

INVX1 _17436_ (
    .A(\datapath.registers.838[15] [19]),
    .Y(_6779_)
);

AOI21X1 _17437_ (
    .A(_5762__bF$buf37),
    .B(\datapath.registers.838[14] [19]),
    .C(_5756__bF$buf2),
    .Y(_6780_)
);

OAI21X1 _17438_ (
    .A(_6779_),
    .B(_5762__bF$buf36),
    .C(_6780_),
    .Y(_6781_)
);

NAND2X1 _17439_ (
    .A(\datapath.registers.838[12] [19]),
    .B(_5762__bF$buf35),
    .Y(_6782_)
);

AOI21X1 _17440_ (
    .A(\datapath.registers.838[13] [19]),
    .B(\datapath.idinstr_15_bF$buf19 ),
    .C(\datapath.idinstr_16_bF$buf25 ),
    .Y(_6783_)
);

AOI21X1 _17441_ (
    .A(_6782_),
    .B(_6783_),
    .C(_5757__bF$buf5),
    .Y(_6784_)
);

AOI22X1 _17442_ (
    .A(_6781_),
    .B(_6784_),
    .C(_5757__bF$buf4),
    .D(_6778_),
    .Y(_6785_)
);

NOR2X1 _17443_ (
    .A(\datapath.registers.838[0] [19]),
    .B(\datapath.idinstr_15_bF$buf18 ),
    .Y(_6786_)
);

OAI21X1 _17444_ (
    .A(\datapath.registers.838[1] [19]),
    .B(_5762__bF$buf34),
    .C(_5756__bF$buf1),
    .Y(_6787_)
);

NOR2X1 _17445_ (
    .A(\datapath.registers.838[3] [19]),
    .B(_5762__bF$buf33),
    .Y(_6788_)
);

OAI21X1 _17446_ (
    .A(\datapath.registers.838[2] [19]),
    .B(\datapath.idinstr_15_bF$buf17 ),
    .C(\datapath.idinstr_16_bF$buf24 ),
    .Y(_6789_)
);

OAI22X1 _17447_ (
    .A(_6788_),
    .B(_6789_),
    .C(_6786_),
    .D(_6787_),
    .Y(_6790_)
);

NOR2X1 _17448_ (
    .A(\datapath.idinstr_17_bF$buf6 ),
    .B(_6790_),
    .Y(_6791_)
);

MUX2X1 _17449_ (
    .A(\datapath.registers.838[5] [19]),
    .B(\datapath.registers.838[4] [19]),
    .S(\datapath.idinstr_15_bF$buf16 ),
    .Y(_6792_)
);

NOR2X1 _17450_ (
    .A(\datapath.registers.838[7] [19]),
    .B(_5762__bF$buf32),
    .Y(_6793_)
);

OAI21X1 _17451_ (
    .A(\datapath.registers.838[6] [19]),
    .B(\datapath.idinstr_15_bF$buf15 ),
    .C(\datapath.idinstr_16_bF$buf23 ),
    .Y(_6794_)
);

OAI22X1 _17452_ (
    .A(_6794_),
    .B(_6793_),
    .C(\datapath.idinstr_16_bF$buf22 ),
    .D(_6792_),
    .Y(_6795_)
);

OAI21X1 _17453_ (
    .A(_5757__bF$buf3),
    .B(_6795_),
    .C(_5760__bF$buf7),
    .Y(_6796_)
);

OAI22X1 _17454_ (
    .A(_5760__bF$buf6),
    .B(_6785_),
    .C(_6791_),
    .D(_6796_),
    .Y(_6797_)
);

NAND2X1 _17455_ (
    .A(_5789__bF$buf0),
    .B(_6797_),
    .Y(_6798_)
);

AOI22X1 _17456_ (
    .A(_5755__bF$buf0),
    .B(_5759__bF$buf0),
    .C(_6774_),
    .D(_6798_),
    .Y(\datapath.registers.rega_data [19])
);

MUX2X1 _17457_ (
    .A(\datapath.registers.838[9] [20]),
    .B(\datapath.registers.838[8] [20]),
    .S(\datapath.idinstr_15_bF$buf14 ),
    .Y(_6799_)
);

NOR2X1 _17458_ (
    .A(\datapath.registers.838[11] [20]),
    .B(_5762__bF$buf31),
    .Y(_6800_)
);

OAI21X1 _17459_ (
    .A(\datapath.registers.838[10] [20]),
    .B(\datapath.idinstr_15_bF$buf13 ),
    .C(\datapath.idinstr_16_bF$buf21 ),
    .Y(_6801_)
);

OAI22X1 _17460_ (
    .A(_6801_),
    .B(_6800_),
    .C(\datapath.idinstr_16_bF$buf20 ),
    .D(_6799_),
    .Y(_6802_)
);

INVX1 _17461_ (
    .A(\datapath.registers.838[15] [20]),
    .Y(_6803_)
);

AOI21X1 _17462_ (
    .A(_5762__bF$buf30),
    .B(\datapath.registers.838[14] [20]),
    .C(_5756__bF$buf0),
    .Y(_6804_)
);

OAI21X1 _17463_ (
    .A(_6803_),
    .B(_5762__bF$buf29),
    .C(_6804_),
    .Y(_6805_)
);

NAND2X1 _17464_ (
    .A(\datapath.registers.838[12] [20]),
    .B(_5762__bF$buf28),
    .Y(_6806_)
);

AOI21X1 _17465_ (
    .A(\datapath.registers.838[13] [20]),
    .B(\datapath.idinstr_15_bF$buf12 ),
    .C(\datapath.idinstr_16_bF$buf19 ),
    .Y(_6807_)
);

AOI21X1 _17466_ (
    .A(_6806_),
    .B(_6807_),
    .C(_5757__bF$buf2),
    .Y(_6808_)
);

AOI22X1 _17467_ (
    .A(_6805_),
    .B(_6808_),
    .C(_5757__bF$buf1),
    .D(_6802_),
    .Y(_6809_)
);

NOR2X1 _17468_ (
    .A(\datapath.registers.838[0] [20]),
    .B(\datapath.idinstr_15_bF$buf11 ),
    .Y(_6810_)
);

OAI21X1 _17469_ (
    .A(\datapath.registers.838[1] [20]),
    .B(_5762__bF$buf27),
    .C(_5756__bF$buf9),
    .Y(_6811_)
);

NOR2X1 _17470_ (
    .A(\datapath.registers.838[3] [20]),
    .B(_5762__bF$buf26),
    .Y(_6812_)
);

OAI21X1 _17471_ (
    .A(\datapath.registers.838[2] [20]),
    .B(\datapath.idinstr_15_bF$buf10 ),
    .C(\datapath.idinstr_16_bF$buf18 ),
    .Y(_6813_)
);

OAI22X1 _17472_ (
    .A(_6812_),
    .B(_6813_),
    .C(_6810_),
    .D(_6811_),
    .Y(_6814_)
);

NOR2X1 _17473_ (
    .A(\datapath.idinstr_17_bF$buf5 ),
    .B(_6814_),
    .Y(_6815_)
);

MUX2X1 _17474_ (
    .A(\datapath.registers.838[5] [20]),
    .B(\datapath.registers.838[4] [20]),
    .S(\datapath.idinstr_15_bF$buf9 ),
    .Y(_6816_)
);

NOR2X1 _17475_ (
    .A(\datapath.registers.838[7] [20]),
    .B(_5762__bF$buf25),
    .Y(_6817_)
);

OAI21X1 _17476_ (
    .A(\datapath.registers.838[6] [20]),
    .B(\datapath.idinstr_15_bF$buf8 ),
    .C(\datapath.idinstr_16_bF$buf17 ),
    .Y(_6818_)
);

OAI22X1 _17477_ (
    .A(_6818_),
    .B(_6817_),
    .C(\datapath.idinstr_16_bF$buf16 ),
    .D(_6816_),
    .Y(_6819_)
);

OAI21X1 _17478_ (
    .A(_5757__bF$buf0),
    .B(_6819_),
    .C(_5760__bF$buf5),
    .Y(_6820_)
);

OAI22X1 _17479_ (
    .A(_5760__bF$buf4),
    .B(_6809_),
    .C(_6815_),
    .D(_6820_),
    .Y(_6821_)
);

NAND2X1 _17480_ (
    .A(_5789__bF$buf4),
    .B(_6821_),
    .Y(_6822_)
);

INVX1 _17481_ (
    .A(\datapath.registers.838[27] [20]),
    .Y(_6823_)
);

AOI21X1 _17482_ (
    .A(\datapath.registers.838[31] [20]),
    .B(\datapath.idinstr_17_bF$buf4 ),
    .C(_5762__bF$buf24),
    .Y(_6824_)
);

OAI21X1 _17483_ (
    .A(\datapath.idinstr_17_bF$buf3 ),
    .B(_6823_),
    .C(_6824_),
    .Y(_6825_)
);

INVX1 _17484_ (
    .A(\datapath.registers.838[26] [20]),
    .Y(_6826_)
);

AOI21X1 _17485_ (
    .A(\datapath.registers.838[30] [20]),
    .B(\datapath.idinstr_17_bF$buf2 ),
    .C(\datapath.idinstr_15_bF$buf7 ),
    .Y(_6827_)
);

OAI21X1 _17486_ (
    .A(\datapath.idinstr_17_bF$buf1 ),
    .B(_6826_),
    .C(_6827_),
    .Y(_6828_)
);

NAND3X1 _17487_ (
    .A(\datapath.idinstr_16_bF$buf15 ),
    .B(_6828_),
    .C(_6825_),
    .Y(_6829_)
);

INVX1 _17488_ (
    .A(\datapath.registers.838[25] [20]),
    .Y(_6830_)
);

AOI21X1 _17489_ (
    .A(\datapath.idinstr_17_bF$buf0 ),
    .B(\datapath.registers.838[29] [20]),
    .C(_5762__bF$buf23),
    .Y(_6831_)
);

OAI21X1 _17490_ (
    .A(\datapath.idinstr_17_bF$buf15 ),
    .B(_6830_),
    .C(_6831_),
    .Y(_6832_)
);

INVX1 _17491_ (
    .A(\datapath.registers.838[24] [20]),
    .Y(_6833_)
);

AOI21X1 _17492_ (
    .A(\datapath.idinstr_17_bF$buf14 ),
    .B(\datapath.registers.838[28] [20]),
    .C(\datapath.idinstr_15_bF$buf6 ),
    .Y(_6834_)
);

OAI21X1 _17493_ (
    .A(_6833_),
    .B(\datapath.idinstr_17_bF$buf13 ),
    .C(_6834_),
    .Y(_6835_)
);

NAND3X1 _17494_ (
    .A(_5756__bF$buf8),
    .B(_6835_),
    .C(_6832_),
    .Y(_6836_)
);

AOI21X1 _17495_ (
    .A(_6829_),
    .B(_6836_),
    .C(_5760__bF$buf3),
    .Y(_6837_)
);

MUX2X1 _17496_ (
    .A(\datapath.registers.838[18] [20]),
    .B(\datapath.registers.838[16] [20]),
    .S(\datapath.idinstr_16_bF$buf14 ),
    .Y(_6838_)
);

NAND2X1 _17497_ (
    .A(_5762__bF$buf22),
    .B(_6838_),
    .Y(_6839_)
);

MUX2X1 _17498_ (
    .A(\datapath.registers.838[19] [20]),
    .B(\datapath.registers.838[17] [20]),
    .S(\datapath.idinstr_16_bF$buf13 ),
    .Y(_6840_)
);

NAND2X1 _17499_ (
    .A(\datapath.idinstr_15_bF$buf5 ),
    .B(_6840_),
    .Y(_6841_)
);

NAND3X1 _17500_ (
    .A(_5757__bF$buf10),
    .B(_6839_),
    .C(_6841_),
    .Y(_6842_)
);

MUX2X1 _17501_ (
    .A(\datapath.registers.838[22] [20]),
    .B(\datapath.registers.838[20] [20]),
    .S(\datapath.idinstr_16_bF$buf12 ),
    .Y(_6843_)
);

NAND2X1 _17502_ (
    .A(_5762__bF$buf21),
    .B(_6843_),
    .Y(_6844_)
);

MUX2X1 _17503_ (
    .A(\datapath.registers.838[23] [20]),
    .B(\datapath.registers.838[21] [20]),
    .S(\datapath.idinstr_16_bF$buf11 ),
    .Y(_6845_)
);

NAND2X1 _17504_ (
    .A(\datapath.idinstr_15_bF$buf4 ),
    .B(_6845_),
    .Y(_6846_)
);

NAND3X1 _17505_ (
    .A(\datapath.idinstr_17_bF$buf12 ),
    .B(_6844_),
    .C(_6846_),
    .Y(_6847_)
);

AOI21X1 _17506_ (
    .A(_6842_),
    .B(_6847_),
    .C(\datapath.idinstr_18_bF$buf6 ),
    .Y(_6848_)
);

OAI21X1 _17507_ (
    .A(_6837_),
    .B(_6848_),
    .C(\datapath.idinstr_19_bF$buf4 ),
    .Y(_6849_)
);

AOI22X1 _17508_ (
    .A(_5755__bF$buf4),
    .B(_5759__bF$buf4),
    .C(_6849_),
    .D(_6822_),
    .Y(\datapath.registers.rega_data [20])
);

NAND2X1 _17509_ (
    .A(\datapath.idinstr_15_bF$buf3 ),
    .B(\datapath.registers.838[27] [21]),
    .Y(_6850_)
);

NAND2X1 _17510_ (
    .A(\datapath.registers.838[26] [21]),
    .B(_5762__bF$buf20),
    .Y(_6851_)
);

NAND3X1 _17511_ (
    .A(\datapath.idinstr_16_bF$buf10 ),
    .B(_6850_),
    .C(_6851_),
    .Y(_6852_)
);

NAND2X1 _17512_ (
    .A(\datapath.idinstr_15_bF$buf2 ),
    .B(\datapath.registers.838[25] [21]),
    .Y(_6853_)
);

AOI21X1 _17513_ (
    .A(_5762__bF$buf19),
    .B(\datapath.registers.838[24] [21]),
    .C(\datapath.idinstr_16_bF$buf9 ),
    .Y(_6854_)
);

NAND2X1 _17514_ (
    .A(_6853_),
    .B(_6854_),
    .Y(_6855_)
);

NAND3X1 _17515_ (
    .A(_5757__bF$buf9),
    .B(_6852_),
    .C(_6855_),
    .Y(_6856_)
);

NAND2X1 _17516_ (
    .A(\datapath.registers.838[31] [21]),
    .B(\datapath.idinstr_15_bF$buf1 ),
    .Y(_6857_)
);

AOI21X1 _17517_ (
    .A(_5762__bF$buf18),
    .B(\datapath.registers.838[30] [21]),
    .C(_5756__bF$buf7),
    .Y(_6858_)
);

NAND2X1 _17518_ (
    .A(_6857_),
    .B(_6858_),
    .Y(_6859_)
);

INVX1 _17519_ (
    .A(\datapath.registers.838[28] [21]),
    .Y(_6860_)
);

AOI21X1 _17520_ (
    .A(\datapath.idinstr_15_bF$buf0 ),
    .B(\datapath.registers.838[29] [21]),
    .C(\datapath.idinstr_16_bF$buf8 ),
    .Y(_6861_)
);

OAI21X1 _17521_ (
    .A(\datapath.idinstr_15_bF$buf54 ),
    .B(_6860_),
    .C(_6861_),
    .Y(_6862_)
);

NAND3X1 _17522_ (
    .A(\datapath.idinstr_17_bF$buf11 ),
    .B(_6862_),
    .C(_6859_),
    .Y(_6863_)
);

AOI21X1 _17523_ (
    .A(_6856_),
    .B(_6863_),
    .C(_5760__bF$buf2),
    .Y(_6864_)
);

MUX2X1 _17524_ (
    .A(\datapath.registers.838[17] [21]),
    .B(\datapath.registers.838[16] [21]),
    .S(\datapath.idinstr_15_bF$buf53 ),
    .Y(_6865_)
);

NOR2X1 _17525_ (
    .A(\datapath.registers.838[19] [21]),
    .B(_5762__bF$buf17),
    .Y(_6866_)
);

OAI21X1 _17526_ (
    .A(\datapath.registers.838[18] [21]),
    .B(\datapath.idinstr_15_bF$buf52 ),
    .C(\datapath.idinstr_16_bF$buf7 ),
    .Y(_6867_)
);

OAI22X1 _17527_ (
    .A(_6867_),
    .B(_6866_),
    .C(\datapath.idinstr_16_bF$buf6 ),
    .D(_6865_),
    .Y(_6868_)
);

NAND2X1 _17528_ (
    .A(_5757__bF$buf8),
    .B(_6868_),
    .Y(_6869_)
);

MUX2X1 _17529_ (
    .A(\datapath.registers.838[21] [21]),
    .B(\datapath.registers.838[20] [21]),
    .S(\datapath.idinstr_15_bF$buf51 ),
    .Y(_6870_)
);

NOR2X1 _17530_ (
    .A(\datapath.registers.838[23] [21]),
    .B(_5762__bF$buf16),
    .Y(_6871_)
);

OAI21X1 _17531_ (
    .A(\datapath.registers.838[22] [21]),
    .B(\datapath.idinstr_15_bF$buf50 ),
    .C(\datapath.idinstr_16_bF$buf5 ),
    .Y(_6872_)
);

OAI22X1 _17532_ (
    .A(_6872_),
    .B(_6871_),
    .C(\datapath.idinstr_16_bF$buf4 ),
    .D(_6870_),
    .Y(_6873_)
);

NAND2X1 _17533_ (
    .A(\datapath.idinstr_17_bF$buf10 ),
    .B(_6873_),
    .Y(_6874_)
);

AOI21X1 _17534_ (
    .A(_6869_),
    .B(_6874_),
    .C(\datapath.idinstr_18_bF$buf5 ),
    .Y(_6875_)
);

OAI21X1 _17535_ (
    .A(_6864_),
    .B(_6875_),
    .C(\datapath.idinstr_19_bF$buf3 ),
    .Y(_6876_)
);

NAND2X1 _17536_ (
    .A(\datapath.registers.838[11] [21]),
    .B(\datapath.idinstr_16_bF$buf3 ),
    .Y(_6877_)
);

NAND2X1 _17537_ (
    .A(\datapath.registers.838[9] [21]),
    .B(_5756__bF$buf6),
    .Y(_6878_)
);

NAND3X1 _17538_ (
    .A(\datapath.idinstr_15_bF$buf49 ),
    .B(_6877_),
    .C(_6878_),
    .Y(_6879_)
);

NAND2X1 _17539_ (
    .A(\datapath.registers.838[10] [21]),
    .B(\datapath.idinstr_16_bF$buf2 ),
    .Y(_6880_)
);

AOI21X1 _17540_ (
    .A(_5756__bF$buf5),
    .B(\datapath.registers.838[8] [21]),
    .C(\datapath.idinstr_15_bF$buf48 ),
    .Y(_6881_)
);

NAND2X1 _17541_ (
    .A(_6880_),
    .B(_6881_),
    .Y(_6882_)
);

NAND3X1 _17542_ (
    .A(_5757__bF$buf7),
    .B(_6879_),
    .C(_6882_),
    .Y(_6883_)
);

NAND2X1 _17543_ (
    .A(\datapath.registers.838[15] [21]),
    .B(\datapath.idinstr_16_bF$buf1 ),
    .Y(_6884_)
);

NAND2X1 _17544_ (
    .A(\datapath.registers.838[13] [21]),
    .B(_5756__bF$buf4),
    .Y(_6885_)
);

NAND3X1 _17545_ (
    .A(\datapath.idinstr_15_bF$buf47 ),
    .B(_6884_),
    .C(_6885_),
    .Y(_6886_)
);

NAND2X1 _17546_ (
    .A(\datapath.registers.838[14] [21]),
    .B(\datapath.idinstr_16_bF$buf0 ),
    .Y(_6887_)
);

AOI21X1 _17547_ (
    .A(_5756__bF$buf3),
    .B(\datapath.registers.838[12] [21]),
    .C(\datapath.idinstr_15_bF$buf46 ),
    .Y(_6888_)
);

NAND2X1 _17548_ (
    .A(_6887_),
    .B(_6888_),
    .Y(_6889_)
);

NAND3X1 _17549_ (
    .A(\datapath.idinstr_17_bF$buf9 ),
    .B(_6886_),
    .C(_6889_),
    .Y(_6890_)
);

AOI21X1 _17550_ (
    .A(_6883_),
    .B(_6890_),
    .C(_5760__bF$buf1),
    .Y(_6891_)
);

INVX1 _17551_ (
    .A(\datapath.registers.838[1] [21]),
    .Y(_6892_)
);

AOI21X1 _17552_ (
    .A(\datapath.registers.838[5] [21]),
    .B(\datapath.idinstr_17_bF$buf8 ),
    .C(_5762__bF$buf15),
    .Y(_6893_)
);

OAI21X1 _17553_ (
    .A(_6892_),
    .B(\datapath.idinstr_17_bF$buf7 ),
    .C(_6893_),
    .Y(_6894_)
);

INVX1 _17554_ (
    .A(\datapath.registers.838[0] [21]),
    .Y(_6895_)
);

AOI21X1 _17555_ (
    .A(\datapath.registers.838[4] [21]),
    .B(\datapath.idinstr_17_bF$buf6 ),
    .C(\datapath.idinstr_15_bF$buf45 ),
    .Y(_6896_)
);

OAI21X1 _17556_ (
    .A(_6895_),
    .B(\datapath.idinstr_17_bF$buf5 ),
    .C(_6896_),
    .Y(_6897_)
);

NAND3X1 _17557_ (
    .A(_5756__bF$buf2),
    .B(_6897_),
    .C(_6894_),
    .Y(_6898_)
);

AOI21X1 _17558_ (
    .A(\datapath.registers.838[7] [21]),
    .B(\datapath.idinstr_17_bF$buf4 ),
    .C(_5762__bF$buf14),
    .Y(_6899_)
);

OAI21X1 _17559_ (
    .A(_5536_),
    .B(\datapath.idinstr_17_bF$buf3 ),
    .C(_6899_),
    .Y(_6900_)
);

INVX1 _17560_ (
    .A(\datapath.registers.838[2] [21]),
    .Y(_6901_)
);

AOI21X1 _17561_ (
    .A(\datapath.registers.838[6] [21]),
    .B(\datapath.idinstr_17_bF$buf2 ),
    .C(\datapath.idinstr_15_bF$buf44 ),
    .Y(_6902_)
);

OAI21X1 _17562_ (
    .A(_6901_),
    .B(\datapath.idinstr_17_bF$buf1 ),
    .C(_6902_),
    .Y(_6903_)
);

NAND3X1 _17563_ (
    .A(\datapath.idinstr_16_bF$buf51 ),
    .B(_6903_),
    .C(_6900_),
    .Y(_6904_)
);

AOI21X1 _17564_ (
    .A(_6898_),
    .B(_6904_),
    .C(\datapath.idinstr_18_bF$buf4 ),
    .Y(_6905_)
);

OAI21X1 _17565_ (
    .A(_6905_),
    .B(_6891_),
    .C(_5789__bF$buf3),
    .Y(_6906_)
);

AOI22X1 _17566_ (
    .A(_5755__bF$buf3),
    .B(_5759__bF$buf3),
    .C(_6906_),
    .D(_6876_),
    .Y(\datapath.registers.rega_data [21])
);

MUX2X1 _17567_ (
    .A(\datapath.registers.838[9] [22]),
    .B(\datapath.registers.838[8] [22]),
    .S(\datapath.idinstr_15_bF$buf43 ),
    .Y(_6907_)
);

NOR2X1 _17568_ (
    .A(\datapath.registers.838[11] [22]),
    .B(_5762__bF$buf13),
    .Y(_6908_)
);

OAI21X1 _17569_ (
    .A(\datapath.registers.838[10] [22]),
    .B(\datapath.idinstr_15_bF$buf42 ),
    .C(\datapath.idinstr_16_bF$buf50 ),
    .Y(_6909_)
);

OAI22X1 _17570_ (
    .A(_6909_),
    .B(_6908_),
    .C(\datapath.idinstr_16_bF$buf49 ),
    .D(_6907_),
    .Y(_6910_)
);

INVX1 _17571_ (
    .A(\datapath.registers.838[15] [22]),
    .Y(_6911_)
);

AOI21X1 _17572_ (
    .A(_5762__bF$buf12),
    .B(\datapath.registers.838[14] [22]),
    .C(_5756__bF$buf1),
    .Y(_6912_)
);

OAI21X1 _17573_ (
    .A(_6911_),
    .B(_5762__bF$buf11),
    .C(_6912_),
    .Y(_6913_)
);

NAND2X1 _17574_ (
    .A(\datapath.registers.838[12] [22]),
    .B(_5762__bF$buf10),
    .Y(_6914_)
);

AOI21X1 _17575_ (
    .A(\datapath.registers.838[13] [22]),
    .B(\datapath.idinstr_15_bF$buf41 ),
    .C(\datapath.idinstr_16_bF$buf48 ),
    .Y(_6915_)
);

AOI21X1 _17576_ (
    .A(_6914_),
    .B(_6915_),
    .C(_5757__bF$buf6),
    .Y(_6916_)
);

AOI22X1 _17577_ (
    .A(_6913_),
    .B(_6916_),
    .C(_5757__bF$buf5),
    .D(_6910_),
    .Y(_6917_)
);

NOR2X1 _17578_ (
    .A(\datapath.registers.838[0] [22]),
    .B(\datapath.idinstr_15_bF$buf40 ),
    .Y(_6918_)
);

OAI21X1 _17579_ (
    .A(\datapath.registers.838[1] [22]),
    .B(_5762__bF$buf9),
    .C(_5756__bF$buf0),
    .Y(_6919_)
);

NOR2X1 _17580_ (
    .A(\datapath.registers.838[3] [22]),
    .B(_5762__bF$buf8),
    .Y(_6920_)
);

OAI21X1 _17581_ (
    .A(\datapath.registers.838[2] [22]),
    .B(\datapath.idinstr_15_bF$buf39 ),
    .C(\datapath.idinstr_16_bF$buf47 ),
    .Y(_6921_)
);

OAI22X1 _17582_ (
    .A(_6920_),
    .B(_6921_),
    .C(_6918_),
    .D(_6919_),
    .Y(_6922_)
);

NOR2X1 _17583_ (
    .A(\datapath.idinstr_17_bF$buf0 ),
    .B(_6922_),
    .Y(_6923_)
);

MUX2X1 _17584_ (
    .A(\datapath.registers.838[5] [22]),
    .B(\datapath.registers.838[4] [22]),
    .S(\datapath.idinstr_15_bF$buf38 ),
    .Y(_6924_)
);

NOR2X1 _17585_ (
    .A(\datapath.registers.838[7] [22]),
    .B(_5762__bF$buf7),
    .Y(_6925_)
);

OAI21X1 _17586_ (
    .A(\datapath.registers.838[6] [22]),
    .B(\datapath.idinstr_15_bF$buf37 ),
    .C(\datapath.idinstr_16_bF$buf46 ),
    .Y(_6926_)
);

OAI22X1 _17587_ (
    .A(_6926_),
    .B(_6925_),
    .C(\datapath.idinstr_16_bF$buf45 ),
    .D(_6924_),
    .Y(_6927_)
);

OAI21X1 _17588_ (
    .A(_5757__bF$buf4),
    .B(_6927_),
    .C(_5760__bF$buf0),
    .Y(_6928_)
);

OAI22X1 _17589_ (
    .A(_5760__bF$buf7),
    .B(_6917_),
    .C(_6923_),
    .D(_6928_),
    .Y(_6929_)
);

NAND2X1 _17590_ (
    .A(_5789__bF$buf2),
    .B(_6929_),
    .Y(_6930_)
);

INVX1 _17591_ (
    .A(\datapath.registers.838[19] [22]),
    .Y(_6931_)
);

AOI21X1 _17592_ (
    .A(\datapath.registers.838[23] [22]),
    .B(\datapath.idinstr_17_bF$buf15 ),
    .C(_5762__bF$buf6),
    .Y(_6932_)
);

OAI21X1 _17593_ (
    .A(_6931_),
    .B(\datapath.idinstr_17_bF$buf14 ),
    .C(_6932_),
    .Y(_6933_)
);

NAND2X1 _17594_ (
    .A(\datapath.registers.838[18] [22]),
    .B(_5757__bF$buf3),
    .Y(_6934_)
);

AOI21X1 _17595_ (
    .A(\datapath.registers.838[22] [22]),
    .B(\datapath.idinstr_17_bF$buf13 ),
    .C(\datapath.idinstr_15_bF$buf36 ),
    .Y(_6935_)
);

AOI21X1 _17596_ (
    .A(_6934_),
    .B(_6935_),
    .C(_5756__bF$buf9),
    .Y(_6936_)
);

AOI21X1 _17597_ (
    .A(\datapath.registers.838[21] [22]),
    .B(\datapath.idinstr_17_bF$buf12 ),
    .C(_5762__bF$buf5),
    .Y(_6937_)
);

OAI21X1 _17598_ (
    .A(_5000_),
    .B(\datapath.idinstr_17_bF$buf11 ),
    .C(_6937_),
    .Y(_6938_)
);

NAND2X1 _17599_ (
    .A(\datapath.registers.838[16] [22]),
    .B(_5757__bF$buf2),
    .Y(_6939_)
);

AOI21X1 _17600_ (
    .A(\datapath.registers.838[20] [22]),
    .B(\datapath.idinstr_17_bF$buf10 ),
    .C(\datapath.idinstr_15_bF$buf35 ),
    .Y(_6940_)
);

AOI21X1 _17601_ (
    .A(_6939_),
    .B(_6940_),
    .C(\datapath.idinstr_16_bF$buf44 ),
    .Y(_6941_)
);

AOI22X1 _17602_ (
    .A(_6936_),
    .B(_6933_),
    .C(_6938_),
    .D(_6941_),
    .Y(_6942_)
);

NOR2X1 _17603_ (
    .A(\datapath.registers.838[24] [22]),
    .B(\datapath.idinstr_15_bF$buf34 ),
    .Y(_6943_)
);

OAI21X1 _17604_ (
    .A(\datapath.registers.838[25] [22]),
    .B(_5762__bF$buf4),
    .C(_5756__bF$buf8),
    .Y(_6944_)
);

NOR2X1 _17605_ (
    .A(\datapath.registers.838[27] [22]),
    .B(_5762__bF$buf3),
    .Y(_6945_)
);

OAI21X1 _17606_ (
    .A(\datapath.idinstr_15_bF$buf33 ),
    .B(\datapath.registers.838[26] [22]),
    .C(\datapath.idinstr_16_bF$buf43 ),
    .Y(_6946_)
);

OAI22X1 _17607_ (
    .A(_6945_),
    .B(_6946_),
    .C(_6943_),
    .D(_6944_),
    .Y(_6947_)
);

NOR2X1 _17608_ (
    .A(\datapath.idinstr_17_bF$buf9 ),
    .B(_6947_),
    .Y(_6948_)
);

MUX2X1 _17609_ (
    .A(\datapath.registers.838[29] [22]),
    .B(\datapath.registers.838[28] [22]),
    .S(\datapath.idinstr_15_bF$buf32 ),
    .Y(_6949_)
);

NOR2X1 _17610_ (
    .A(\datapath.registers.838[31] [22]),
    .B(_5762__bF$buf2),
    .Y(_6950_)
);

OAI21X1 _17611_ (
    .A(\datapath.registers.838[30] [22]),
    .B(\datapath.idinstr_15_bF$buf31 ),
    .C(\datapath.idinstr_16_bF$buf42 ),
    .Y(_6951_)
);

OAI22X1 _17612_ (
    .A(_6951_),
    .B(_6950_),
    .C(\datapath.idinstr_16_bF$buf41 ),
    .D(_6949_),
    .Y(_6952_)
);

OAI21X1 _17613_ (
    .A(_5757__bF$buf1),
    .B(_6952_),
    .C(\datapath.idinstr_18_bF$buf3 ),
    .Y(_6953_)
);

OAI22X1 _17614_ (
    .A(\datapath.idinstr_18_bF$buf2 ),
    .B(_6942_),
    .C(_6948_),
    .D(_6953_),
    .Y(_6954_)
);

NAND2X1 _17615_ (
    .A(\datapath.idinstr_19_bF$buf2 ),
    .B(_6954_),
    .Y(_6955_)
);

AOI22X1 _17616_ (
    .A(_5755__bF$buf2),
    .B(_5759__bF$buf2),
    .C(_6955_),
    .D(_6930_),
    .Y(\datapath.registers.rega_data [22])
);

MUX2X1 _17617_ (
    .A(\datapath.registers.838[9] [23]),
    .B(\datapath.registers.838[8] [23]),
    .S(\datapath.idinstr_15_bF$buf30 ),
    .Y(_6956_)
);

NOR2X1 _17618_ (
    .A(\datapath.registers.838[11] [23]),
    .B(_5762__bF$buf1),
    .Y(_6957_)
);

OAI21X1 _17619_ (
    .A(\datapath.registers.838[10] [23]),
    .B(\datapath.idinstr_15_bF$buf29 ),
    .C(\datapath.idinstr_16_bF$buf40 ),
    .Y(_6958_)
);

OAI22X1 _17620_ (
    .A(_6958_),
    .B(_6957_),
    .C(\datapath.idinstr_16_bF$buf39 ),
    .D(_6956_),
    .Y(_6959_)
);

INVX1 _17621_ (
    .A(\datapath.registers.838[15] [23]),
    .Y(_6960_)
);

AOI21X1 _17622_ (
    .A(_5762__bF$buf0),
    .B(\datapath.registers.838[14] [23]),
    .C(_5756__bF$buf7),
    .Y(_6961_)
);

OAI21X1 _17623_ (
    .A(_6960_),
    .B(_5762__bF$buf47),
    .C(_6961_),
    .Y(_6962_)
);

NAND2X1 _17624_ (
    .A(\datapath.registers.838[12] [23]),
    .B(_5762__bF$buf46),
    .Y(_6963_)
);

AOI21X1 _17625_ (
    .A(\datapath.registers.838[13] [23]),
    .B(\datapath.idinstr_15_bF$buf28 ),
    .C(\datapath.idinstr_16_bF$buf38 ),
    .Y(_6964_)
);

AOI21X1 _17626_ (
    .A(_6963_),
    .B(_6964_),
    .C(_5757__bF$buf0),
    .Y(_6965_)
);

AOI22X1 _17627_ (
    .A(_6962_),
    .B(_6965_),
    .C(_5757__bF$buf10),
    .D(_6959_),
    .Y(_6966_)
);

NOR2X1 _17628_ (
    .A(\datapath.registers.838[0] [23]),
    .B(\datapath.idinstr_15_bF$buf27 ),
    .Y(_6967_)
);

OAI21X1 _17629_ (
    .A(\datapath.registers.838[1] [23]),
    .B(_5762__bF$buf45),
    .C(_5756__bF$buf6),
    .Y(_6968_)
);

NOR2X1 _17630_ (
    .A(\datapath.registers.838[3] [23]),
    .B(_5762__bF$buf44),
    .Y(_6969_)
);

OAI21X1 _17631_ (
    .A(\datapath.registers.838[2] [23]),
    .B(\datapath.idinstr_15_bF$buf26 ),
    .C(\datapath.idinstr_16_bF$buf37 ),
    .Y(_6970_)
);

OAI22X1 _17632_ (
    .A(_6969_),
    .B(_6970_),
    .C(_6967_),
    .D(_6968_),
    .Y(_6971_)
);

NOR2X1 _17633_ (
    .A(\datapath.idinstr_17_bF$buf8 ),
    .B(_6971_),
    .Y(_6972_)
);

MUX2X1 _17634_ (
    .A(\datapath.registers.838[5] [23]),
    .B(\datapath.registers.838[4] [23]),
    .S(\datapath.idinstr_15_bF$buf25 ),
    .Y(_6973_)
);

NOR2X1 _17635_ (
    .A(\datapath.registers.838[7] [23]),
    .B(_5762__bF$buf43),
    .Y(_6974_)
);

OAI21X1 _17636_ (
    .A(\datapath.registers.838[6] [23]),
    .B(\datapath.idinstr_15_bF$buf24 ),
    .C(\datapath.idinstr_16_bF$buf36 ),
    .Y(_6975_)
);

OAI22X1 _17637_ (
    .A(_6975_),
    .B(_6974_),
    .C(\datapath.idinstr_16_bF$buf35 ),
    .D(_6973_),
    .Y(_6976_)
);

OAI21X1 _17638_ (
    .A(_5757__bF$buf9),
    .B(_6976_),
    .C(_5760__bF$buf6),
    .Y(_6977_)
);

OAI22X1 _17639_ (
    .A(_5760__bF$buf5),
    .B(_6966_),
    .C(_6972_),
    .D(_6977_),
    .Y(_6978_)
);

NAND2X1 _17640_ (
    .A(_5789__bF$buf1),
    .B(_6978_),
    .Y(_6979_)
);

INVX1 _17641_ (
    .A(\datapath.registers.838[27] [23]),
    .Y(_6980_)
);

AOI21X1 _17642_ (
    .A(\datapath.registers.838[31] [23]),
    .B(\datapath.idinstr_17_bF$buf7 ),
    .C(_5762__bF$buf42),
    .Y(_6981_)
);

OAI21X1 _17643_ (
    .A(\datapath.idinstr_17_bF$buf6 ),
    .B(_6980_),
    .C(_6981_),
    .Y(_6982_)
);

INVX1 _17644_ (
    .A(\datapath.registers.838[26] [23]),
    .Y(_6983_)
);

AOI21X1 _17645_ (
    .A(\datapath.registers.838[30] [23]),
    .B(\datapath.idinstr_17_bF$buf5 ),
    .C(\datapath.idinstr_15_bF$buf23 ),
    .Y(_6984_)
);

OAI21X1 _17646_ (
    .A(\datapath.idinstr_17_bF$buf4 ),
    .B(_6983_),
    .C(_6984_),
    .Y(_6985_)
);

NAND3X1 _17647_ (
    .A(\datapath.idinstr_16_bF$buf34 ),
    .B(_6985_),
    .C(_6982_),
    .Y(_6986_)
);

INVX1 _17648_ (
    .A(\datapath.registers.838[25] [23]),
    .Y(_6987_)
);

AOI21X1 _17649_ (
    .A(\datapath.idinstr_17_bF$buf3 ),
    .B(\datapath.registers.838[29] [23]),
    .C(_5762__bF$buf41),
    .Y(_6988_)
);

OAI21X1 _17650_ (
    .A(\datapath.idinstr_17_bF$buf2 ),
    .B(_6987_),
    .C(_6988_),
    .Y(_6989_)
);

INVX1 _17651_ (
    .A(\datapath.registers.838[24] [23]),
    .Y(_6990_)
);

AOI21X1 _17652_ (
    .A(\datapath.idinstr_17_bF$buf1 ),
    .B(\datapath.registers.838[28] [23]),
    .C(\datapath.idinstr_15_bF$buf22 ),
    .Y(_6991_)
);

OAI21X1 _17653_ (
    .A(_6990_),
    .B(\datapath.idinstr_17_bF$buf0 ),
    .C(_6991_),
    .Y(_6992_)
);

NAND3X1 _17654_ (
    .A(_5756__bF$buf5),
    .B(_6992_),
    .C(_6989_),
    .Y(_6993_)
);

AOI21X1 _17655_ (
    .A(_6986_),
    .B(_6993_),
    .C(_5760__bF$buf4),
    .Y(_6994_)
);

MUX2X1 _17656_ (
    .A(\datapath.registers.838[18] [23]),
    .B(\datapath.registers.838[16] [23]),
    .S(\datapath.idinstr_16_bF$buf33 ),
    .Y(_6995_)
);

NAND2X1 _17657_ (
    .A(_5762__bF$buf40),
    .B(_6995_),
    .Y(_6996_)
);

MUX2X1 _17658_ (
    .A(\datapath.registers.838[19] [23]),
    .B(\datapath.registers.838[17] [23]),
    .S(\datapath.idinstr_16_bF$buf32 ),
    .Y(_6997_)
);

NAND2X1 _17659_ (
    .A(\datapath.idinstr_15_bF$buf21 ),
    .B(_6997_),
    .Y(_6998_)
);

NAND3X1 _17660_ (
    .A(_5757__bF$buf8),
    .B(_6996_),
    .C(_6998_),
    .Y(_6999_)
);

MUX2X1 _17661_ (
    .A(\datapath.registers.838[22] [23]),
    .B(\datapath.registers.838[20] [23]),
    .S(\datapath.idinstr_16_bF$buf31 ),
    .Y(_7000_)
);

NAND2X1 _17662_ (
    .A(_5762__bF$buf39),
    .B(_7000_),
    .Y(_7001_)
);

MUX2X1 _17663_ (
    .A(\datapath.registers.838[23] [23]),
    .B(\datapath.registers.838[21] [23]),
    .S(\datapath.idinstr_16_bF$buf30 ),
    .Y(_7002_)
);

NAND2X1 _17664_ (
    .A(\datapath.idinstr_15_bF$buf20 ),
    .B(_7002_),
    .Y(_7003_)
);

NAND3X1 _17665_ (
    .A(\datapath.idinstr_17_bF$buf15 ),
    .B(_7001_),
    .C(_7003_),
    .Y(_7004_)
);

AOI21X1 _17666_ (
    .A(_6999_),
    .B(_7004_),
    .C(\datapath.idinstr_18_bF$buf1 ),
    .Y(_7005_)
);

OAI21X1 _17667_ (
    .A(_6994_),
    .B(_7005_),
    .C(\datapath.idinstr_19_bF$buf1 ),
    .Y(_7006_)
);

AOI22X1 _17668_ (
    .A(_5755__bF$buf1),
    .B(_5759__bF$buf1),
    .C(_7006_),
    .D(_6979_),
    .Y(\datapath.registers.rega_data [23])
);

MUX2X1 _17669_ (
    .A(\datapath.registers.838[2] [24]),
    .B(\datapath.registers.838[0] [24]),
    .S(\datapath.idinstr_16_bF$buf29 ),
    .Y(_7007_)
);

NAND2X1 _17670_ (
    .A(_5762__bF$buf38),
    .B(_7007_),
    .Y(_7008_)
);

MUX2X1 _17671_ (
    .A(\datapath.registers.838[3] [24]),
    .B(\datapath.registers.838[1] [24]),
    .S(\datapath.idinstr_16_bF$buf28 ),
    .Y(_7009_)
);

NAND2X1 _17672_ (
    .A(\datapath.idinstr_15_bF$buf19 ),
    .B(_7009_),
    .Y(_7010_)
);

NAND3X1 _17673_ (
    .A(_5757__bF$buf7),
    .B(_7008_),
    .C(_7010_),
    .Y(_7011_)
);

MUX2X1 _17674_ (
    .A(\datapath.registers.838[6] [24]),
    .B(\datapath.registers.838[4] [24]),
    .S(\datapath.idinstr_16_bF$buf27 ),
    .Y(_7012_)
);

NAND2X1 _17675_ (
    .A(_5762__bF$buf37),
    .B(_7012_),
    .Y(_7013_)
);

MUX2X1 _17676_ (
    .A(\datapath.registers.838[7] [24]),
    .B(\datapath.registers.838[5] [24]),
    .S(\datapath.idinstr_16_bF$buf26 ),
    .Y(_7014_)
);

NAND2X1 _17677_ (
    .A(\datapath.idinstr_15_bF$buf18 ),
    .B(_7014_),
    .Y(_7015_)
);

NAND3X1 _17678_ (
    .A(\datapath.idinstr_17_bF$buf14 ),
    .B(_7013_),
    .C(_7015_),
    .Y(_7016_)
);

AOI21X1 _17679_ (
    .A(_7011_),
    .B(_7016_),
    .C(\datapath.idinstr_18_bF$buf0 ),
    .Y(_7017_)
);

AOI21X1 _17680_ (
    .A(\datapath.registers.838[13] [24]),
    .B(\datapath.idinstr_17_bF$buf13 ),
    .C(_5762__bF$buf36),
    .Y(_7018_)
);

OAI21X1 _17681_ (
    .A(_5297_),
    .B(\datapath.idinstr_17_bF$buf12 ),
    .C(_7018_),
    .Y(_7019_)
);

INVX1 _17682_ (
    .A(\datapath.registers.838[8] [24]),
    .Y(_7020_)
);

AOI21X1 _17683_ (
    .A(\datapath.registers.838[12] [24]),
    .B(\datapath.idinstr_17_bF$buf11 ),
    .C(\datapath.idinstr_15_bF$buf17 ),
    .Y(_7021_)
);

OAI21X1 _17684_ (
    .A(_7020_),
    .B(\datapath.idinstr_17_bF$buf10 ),
    .C(_7021_),
    .Y(_7022_)
);

NAND3X1 _17685_ (
    .A(_5756__bF$buf4),
    .B(_7022_),
    .C(_7019_),
    .Y(_7023_)
);

INVX1 _17686_ (
    .A(\datapath.registers.838[11] [24]),
    .Y(_7024_)
);

AOI21X1 _17687_ (
    .A(\datapath.registers.838[15] [24]),
    .B(\datapath.idinstr_17_bF$buf9 ),
    .C(_5762__bF$buf35),
    .Y(_7025_)
);

OAI21X1 _17688_ (
    .A(_7024_),
    .B(\datapath.idinstr_17_bF$buf8 ),
    .C(_7025_),
    .Y(_7026_)
);

AOI21X1 _17689_ (
    .A(\datapath.registers.838[14] [24]),
    .B(\datapath.idinstr_17_bF$buf7 ),
    .C(\datapath.idinstr_15_bF$buf16 ),
    .Y(_7027_)
);

OAI21X1 _17690_ (
    .A(_5253_),
    .B(\datapath.idinstr_17_bF$buf6 ),
    .C(_7027_),
    .Y(_7028_)
);

NAND3X1 _17691_ (
    .A(\datapath.idinstr_16_bF$buf25 ),
    .B(_7028_),
    .C(_7026_),
    .Y(_7029_)
);

AOI21X1 _17692_ (
    .A(_7023_),
    .B(_7029_),
    .C(_5760__bF$buf3),
    .Y(_7030_)
);

OAI21X1 _17693_ (
    .A(_7030_),
    .B(_7017_),
    .C(_5789__bF$buf0),
    .Y(_7031_)
);

NOR2X1 _17694_ (
    .A(\datapath.registers.838[24] [24]),
    .B(\datapath.idinstr_15_bF$buf15 ),
    .Y(_7032_)
);

OAI21X1 _17695_ (
    .A(\datapath.registers.838[25] [24]),
    .B(_5762__bF$buf34),
    .C(_5756__bF$buf3),
    .Y(_7033_)
);

NOR2X1 _17696_ (
    .A(\datapath.registers.838[27] [24]),
    .B(_5762__bF$buf33),
    .Y(_7034_)
);

OAI21X1 _17697_ (
    .A(\datapath.idinstr_15_bF$buf14 ),
    .B(\datapath.registers.838[26] [24]),
    .C(\datapath.idinstr_16_bF$buf24 ),
    .Y(_7035_)
);

OAI22X1 _17698_ (
    .A(_7034_),
    .B(_7035_),
    .C(_7032_),
    .D(_7033_),
    .Y(_7036_)
);

NOR2X1 _17699_ (
    .A(\datapath.idinstr_17_bF$buf5 ),
    .B(_7036_),
    .Y(_7037_)
);

MUX2X1 _17700_ (
    .A(\datapath.registers.838[29] [24]),
    .B(\datapath.registers.838[28] [24]),
    .S(\datapath.idinstr_15_bF$buf13 ),
    .Y(_7038_)
);

NOR2X1 _17701_ (
    .A(\datapath.registers.838[31] [24]),
    .B(_5762__bF$buf32),
    .Y(_7039_)
);

OAI21X1 _17702_ (
    .A(\datapath.registers.838[30] [24]),
    .B(\datapath.idinstr_15_bF$buf12 ),
    .C(\datapath.idinstr_16_bF$buf23 ),
    .Y(_7040_)
);

OAI22X1 _17703_ (
    .A(_7040_),
    .B(_7039_),
    .C(\datapath.idinstr_16_bF$buf22 ),
    .D(_7038_),
    .Y(_7041_)
);

OAI21X1 _17704_ (
    .A(_5757__bF$buf6),
    .B(_7041_),
    .C(\datapath.idinstr_18_bF$buf6 ),
    .Y(_7042_)
);

INVX1 _17705_ (
    .A(\datapath.registers.838[19] [24]),
    .Y(_7043_)
);

AOI21X1 _17706_ (
    .A(\datapath.registers.838[23] [24]),
    .B(\datapath.idinstr_17_bF$buf4 ),
    .C(_5762__bF$buf31),
    .Y(_7044_)
);

OAI21X1 _17707_ (
    .A(_7043_),
    .B(\datapath.idinstr_17_bF$buf3 ),
    .C(_7044_),
    .Y(_7045_)
);

NAND2X1 _17708_ (
    .A(\datapath.registers.838[18] [24]),
    .B(_5757__bF$buf5),
    .Y(_7046_)
);

AOI21X1 _17709_ (
    .A(\datapath.registers.838[22] [24]),
    .B(\datapath.idinstr_17_bF$buf2 ),
    .C(\datapath.idinstr_15_bF$buf11 ),
    .Y(_7047_)
);

AOI21X1 _17710_ (
    .A(_7046_),
    .B(_7047_),
    .C(_5756__bF$buf2),
    .Y(_7048_)
);

AOI21X1 _17711_ (
    .A(\datapath.registers.838[21] [24]),
    .B(\datapath.idinstr_17_bF$buf1 ),
    .C(_5762__bF$buf30),
    .Y(_7049_)
);

OAI21X1 _17712_ (
    .A(_5004_),
    .B(\datapath.idinstr_17_bF$buf0 ),
    .C(_7049_),
    .Y(_7050_)
);

NAND2X1 _17713_ (
    .A(\datapath.registers.838[16] [24]),
    .B(_5757__bF$buf4),
    .Y(_7051_)
);

AOI21X1 _17714_ (
    .A(\datapath.registers.838[20] [24]),
    .B(\datapath.idinstr_17_bF$buf15 ),
    .C(\datapath.idinstr_15_bF$buf10 ),
    .Y(_7052_)
);

AOI21X1 _17715_ (
    .A(_7051_),
    .B(_7052_),
    .C(\datapath.idinstr_16_bF$buf21 ),
    .Y(_7053_)
);

AOI22X1 _17716_ (
    .A(_7048_),
    .B(_7045_),
    .C(_7050_),
    .D(_7053_),
    .Y(_7054_)
);

OAI22X1 _17717_ (
    .A(\datapath.idinstr_18_bF$buf5 ),
    .B(_7054_),
    .C(_7037_),
    .D(_7042_),
    .Y(_7055_)
);

NAND2X1 _17718_ (
    .A(\datapath.idinstr_19_bF$buf0 ),
    .B(_7055_),
    .Y(_7056_)
);

AOI22X1 _17719_ (
    .A(_5755__bF$buf0),
    .B(_5759__bF$buf0),
    .C(_7031_),
    .D(_7056_),
    .Y(\datapath.registers.rega_data [24])
);

NAND2X1 _17720_ (
    .A(\datapath.idinstr_15_bF$buf9 ),
    .B(\datapath.registers.838[27] [25]),
    .Y(_7057_)
);

NAND2X1 _17721_ (
    .A(\datapath.registers.838[26] [25]),
    .B(_5762__bF$buf29),
    .Y(_7058_)
);

NAND3X1 _17722_ (
    .A(\datapath.idinstr_16_bF$buf20 ),
    .B(_7057_),
    .C(_7058_),
    .Y(_7059_)
);

NAND2X1 _17723_ (
    .A(\datapath.idinstr_15_bF$buf8 ),
    .B(\datapath.registers.838[25] [25]),
    .Y(_7060_)
);

AOI21X1 _17724_ (
    .A(_5762__bF$buf28),
    .B(\datapath.registers.838[24] [25]),
    .C(\datapath.idinstr_16_bF$buf19 ),
    .Y(_7061_)
);

NAND2X1 _17725_ (
    .A(_7060_),
    .B(_7061_),
    .Y(_7062_)
);

NAND3X1 _17726_ (
    .A(_5757__bF$buf3),
    .B(_7059_),
    .C(_7062_),
    .Y(_7063_)
);

NAND2X1 _17727_ (
    .A(\datapath.registers.838[31] [25]),
    .B(\datapath.idinstr_15_bF$buf7 ),
    .Y(_7064_)
);

AOI21X1 _17728_ (
    .A(_5762__bF$buf27),
    .B(\datapath.registers.838[30] [25]),
    .C(_5756__bF$buf1),
    .Y(_7065_)
);

NAND2X1 _17729_ (
    .A(_7064_),
    .B(_7065_),
    .Y(_7066_)
);

INVX1 _17730_ (
    .A(\datapath.registers.838[28] [25]),
    .Y(_7067_)
);

AOI21X1 _17731_ (
    .A(\datapath.idinstr_15_bF$buf6 ),
    .B(\datapath.registers.838[29] [25]),
    .C(\datapath.idinstr_16_bF$buf18 ),
    .Y(_7068_)
);

OAI21X1 _17732_ (
    .A(\datapath.idinstr_15_bF$buf5 ),
    .B(_7067_),
    .C(_7068_),
    .Y(_7069_)
);

NAND3X1 _17733_ (
    .A(\datapath.idinstr_17_bF$buf14 ),
    .B(_7069_),
    .C(_7066_),
    .Y(_7070_)
);

AOI21X1 _17734_ (
    .A(_7063_),
    .B(_7070_),
    .C(_5760__bF$buf2),
    .Y(_7071_)
);

MUX2X1 _17735_ (
    .A(\datapath.registers.838[17] [25]),
    .B(\datapath.registers.838[16] [25]),
    .S(\datapath.idinstr_15_bF$buf4 ),
    .Y(_7072_)
);

NOR2X1 _17736_ (
    .A(\datapath.registers.838[19] [25]),
    .B(_5762__bF$buf26),
    .Y(_7073_)
);

OAI21X1 _17737_ (
    .A(\datapath.registers.838[18] [25]),
    .B(\datapath.idinstr_15_bF$buf3 ),
    .C(\datapath.idinstr_16_bF$buf17 ),
    .Y(_7074_)
);

OAI22X1 _17738_ (
    .A(_7074_),
    .B(_7073_),
    .C(\datapath.idinstr_16_bF$buf16 ),
    .D(_7072_),
    .Y(_7075_)
);

NAND2X1 _17739_ (
    .A(_5757__bF$buf2),
    .B(_7075_),
    .Y(_7076_)
);

MUX2X1 _17740_ (
    .A(\datapath.registers.838[21] [25]),
    .B(\datapath.registers.838[20] [25]),
    .S(\datapath.idinstr_15_bF$buf2 ),
    .Y(_7077_)
);

NOR2X1 _17741_ (
    .A(\datapath.registers.838[23] [25]),
    .B(_5762__bF$buf25),
    .Y(_7078_)
);

OAI21X1 _17742_ (
    .A(\datapath.registers.838[22] [25]),
    .B(\datapath.idinstr_15_bF$buf1 ),
    .C(\datapath.idinstr_16_bF$buf15 ),
    .Y(_7079_)
);

OAI22X1 _17743_ (
    .A(_7079_),
    .B(_7078_),
    .C(\datapath.idinstr_16_bF$buf14 ),
    .D(_7077_),
    .Y(_7080_)
);

NAND2X1 _17744_ (
    .A(\datapath.idinstr_17_bF$buf13 ),
    .B(_7080_),
    .Y(_7081_)
);

AOI21X1 _17745_ (
    .A(_7076_),
    .B(_7081_),
    .C(\datapath.idinstr_18_bF$buf4 ),
    .Y(_7082_)
);

OAI21X1 _17746_ (
    .A(_7071_),
    .B(_7082_),
    .C(\datapath.idinstr_19_bF$buf5 ),
    .Y(_7083_)
);

NAND2X1 _17747_ (
    .A(\datapath.registers.838[11] [25]),
    .B(\datapath.idinstr_16_bF$buf13 ),
    .Y(_7084_)
);

NAND2X1 _17748_ (
    .A(\datapath.registers.838[9] [25]),
    .B(_5756__bF$buf0),
    .Y(_7085_)
);

NAND3X1 _17749_ (
    .A(\datapath.idinstr_15_bF$buf0 ),
    .B(_7084_),
    .C(_7085_),
    .Y(_7086_)
);

NAND2X1 _17750_ (
    .A(\datapath.registers.838[10] [25]),
    .B(\datapath.idinstr_16_bF$buf12 ),
    .Y(_7087_)
);

AOI21X1 _17751_ (
    .A(_5756__bF$buf9),
    .B(\datapath.registers.838[8] [25]),
    .C(\datapath.idinstr_15_bF$buf54 ),
    .Y(_7088_)
);

NAND2X1 _17752_ (
    .A(_7087_),
    .B(_7088_),
    .Y(_7089_)
);

NAND3X1 _17753_ (
    .A(_5757__bF$buf1),
    .B(_7086_),
    .C(_7089_),
    .Y(_7090_)
);

NAND2X1 _17754_ (
    .A(\datapath.registers.838[15] [25]),
    .B(\datapath.idinstr_16_bF$buf11 ),
    .Y(_7091_)
);

NAND2X1 _17755_ (
    .A(\datapath.registers.838[13] [25]),
    .B(_5756__bF$buf8),
    .Y(_7092_)
);

NAND3X1 _17756_ (
    .A(\datapath.idinstr_15_bF$buf53 ),
    .B(_7091_),
    .C(_7092_),
    .Y(_7093_)
);

NAND2X1 _17757_ (
    .A(\datapath.registers.838[14] [25]),
    .B(\datapath.idinstr_16_bF$buf10 ),
    .Y(_7094_)
);

AOI21X1 _17758_ (
    .A(_5756__bF$buf7),
    .B(\datapath.registers.838[12] [25]),
    .C(\datapath.idinstr_15_bF$buf52 ),
    .Y(_7095_)
);

NAND2X1 _17759_ (
    .A(_7094_),
    .B(_7095_),
    .Y(_7096_)
);

NAND3X1 _17760_ (
    .A(\datapath.idinstr_17_bF$buf12 ),
    .B(_7093_),
    .C(_7096_),
    .Y(_7097_)
);

AOI21X1 _17761_ (
    .A(_7090_),
    .B(_7097_),
    .C(_5760__bF$buf1),
    .Y(_7098_)
);

INVX1 _17762_ (
    .A(\datapath.registers.838[1] [25]),
    .Y(_7099_)
);

AOI21X1 _17763_ (
    .A(\datapath.registers.838[5] [25]),
    .B(\datapath.idinstr_17_bF$buf11 ),
    .C(_5762__bF$buf24),
    .Y(_7100_)
);

OAI21X1 _17764_ (
    .A(_7099_),
    .B(\datapath.idinstr_17_bF$buf10 ),
    .C(_7100_),
    .Y(_7101_)
);

INVX1 _17765_ (
    .A(\datapath.registers.838[0] [25]),
    .Y(_7102_)
);

AOI21X1 _17766_ (
    .A(\datapath.registers.838[4] [25]),
    .B(\datapath.idinstr_17_bF$buf9 ),
    .C(\datapath.idinstr_15_bF$buf51 ),
    .Y(_7103_)
);

OAI21X1 _17767_ (
    .A(_7102_),
    .B(\datapath.idinstr_17_bF$buf8 ),
    .C(_7103_),
    .Y(_7104_)
);

NAND3X1 _17768_ (
    .A(_5756__bF$buf6),
    .B(_7104_),
    .C(_7101_),
    .Y(_7105_)
);

AOI21X1 _17769_ (
    .A(\datapath.registers.838[7] [25]),
    .B(\datapath.idinstr_17_bF$buf7 ),
    .C(_5762__bF$buf23),
    .Y(_7106_)
);

OAI21X1 _17770_ (
    .A(_5543_),
    .B(\datapath.idinstr_17_bF$buf6 ),
    .C(_7106_),
    .Y(_7107_)
);

INVX1 _17771_ (
    .A(\datapath.registers.838[2] [25]),
    .Y(_7108_)
);

AOI21X1 _17772_ (
    .A(\datapath.registers.838[6] [25]),
    .B(\datapath.idinstr_17_bF$buf5 ),
    .C(\datapath.idinstr_15_bF$buf50 ),
    .Y(_7109_)
);

OAI21X1 _17773_ (
    .A(_7108_),
    .B(\datapath.idinstr_17_bF$buf4 ),
    .C(_7109_),
    .Y(_7110_)
);

NAND3X1 _17774_ (
    .A(\datapath.idinstr_16_bF$buf9 ),
    .B(_7110_),
    .C(_7107_),
    .Y(_7111_)
);

AOI21X1 _17775_ (
    .A(_7105_),
    .B(_7111_),
    .C(\datapath.idinstr_18_bF$buf3 ),
    .Y(_7112_)
);

OAI21X1 _17776_ (
    .A(_7112_),
    .B(_7098_),
    .C(_5789__bF$buf4),
    .Y(_7113_)
);

AOI22X1 _17777_ (
    .A(_5755__bF$buf4),
    .B(_5759__bF$buf4),
    .C(_7113_),
    .D(_7083_),
    .Y(\datapath.registers.rega_data [25])
);

NAND2X1 _17778_ (
    .A(\datapath.idinstr_15_bF$buf49 ),
    .B(\datapath.registers.838[27] [26]),
    .Y(_7114_)
);

NAND2X1 _17779_ (
    .A(\datapath.registers.838[26] [26]),
    .B(_5762__bF$buf22),
    .Y(_7115_)
);

NAND3X1 _17780_ (
    .A(\datapath.idinstr_16_bF$buf8 ),
    .B(_7114_),
    .C(_7115_),
    .Y(_7116_)
);

NAND2X1 _17781_ (
    .A(\datapath.idinstr_15_bF$buf48 ),
    .B(\datapath.registers.838[25] [26]),
    .Y(_7117_)
);

AOI21X1 _17782_ (
    .A(_5762__bF$buf21),
    .B(\datapath.registers.838[24] [26]),
    .C(\datapath.idinstr_16_bF$buf7 ),
    .Y(_7118_)
);

NAND2X1 _17783_ (
    .A(_7117_),
    .B(_7118_),
    .Y(_7119_)
);

NAND3X1 _17784_ (
    .A(_5757__bF$buf0),
    .B(_7116_),
    .C(_7119_),
    .Y(_7120_)
);

NAND2X1 _17785_ (
    .A(\datapath.registers.838[31] [26]),
    .B(\datapath.idinstr_15_bF$buf47 ),
    .Y(_7121_)
);

AOI21X1 _17786_ (
    .A(_5762__bF$buf20),
    .B(\datapath.registers.838[30] [26]),
    .C(_5756__bF$buf5),
    .Y(_7122_)
);

NAND2X1 _17787_ (
    .A(_7121_),
    .B(_7122_),
    .Y(_7123_)
);

INVX1 _17788_ (
    .A(\datapath.registers.838[28] [26]),
    .Y(_7124_)
);

AOI21X1 _17789_ (
    .A(\datapath.idinstr_15_bF$buf46 ),
    .B(\datapath.registers.838[29] [26]),
    .C(\datapath.idinstr_16_bF$buf6 ),
    .Y(_7125_)
);

OAI21X1 _17790_ (
    .A(\datapath.idinstr_15_bF$buf45 ),
    .B(_7124_),
    .C(_7125_),
    .Y(_7126_)
);

NAND3X1 _17791_ (
    .A(\datapath.idinstr_17_bF$buf3 ),
    .B(_7126_),
    .C(_7123_),
    .Y(_7127_)
);

AOI21X1 _17792_ (
    .A(_7120_),
    .B(_7127_),
    .C(_5760__bF$buf0),
    .Y(_7128_)
);

MUX2X1 _17793_ (
    .A(\datapath.registers.838[18] [26]),
    .B(\datapath.registers.838[16] [26]),
    .S(\datapath.idinstr_16_bF$buf5 ),
    .Y(_7129_)
);

NAND2X1 _17794_ (
    .A(_5762__bF$buf19),
    .B(_7129_),
    .Y(_7130_)
);

MUX2X1 _17795_ (
    .A(\datapath.registers.838[19] [26]),
    .B(\datapath.registers.838[17] [26]),
    .S(\datapath.idinstr_16_bF$buf4 ),
    .Y(_7131_)
);

NAND2X1 _17796_ (
    .A(\datapath.idinstr_15_bF$buf44 ),
    .B(_7131_),
    .Y(_7132_)
);

NAND3X1 _17797_ (
    .A(_5757__bF$buf10),
    .B(_7130_),
    .C(_7132_),
    .Y(_7133_)
);

MUX2X1 _17798_ (
    .A(\datapath.registers.838[22] [26]),
    .B(\datapath.registers.838[20] [26]),
    .S(\datapath.idinstr_16_bF$buf3 ),
    .Y(_7134_)
);

NAND2X1 _17799_ (
    .A(_5762__bF$buf18),
    .B(_7134_),
    .Y(_7135_)
);

MUX2X1 _17800_ (
    .A(\datapath.registers.838[23] [26]),
    .B(\datapath.registers.838[21] [26]),
    .S(\datapath.idinstr_16_bF$buf2 ),
    .Y(_7136_)
);

NAND2X1 _17801_ (
    .A(\datapath.idinstr_15_bF$buf43 ),
    .B(_7136_),
    .Y(_7137_)
);

NAND3X1 _17802_ (
    .A(\datapath.idinstr_17_bF$buf2 ),
    .B(_7135_),
    .C(_7137_),
    .Y(_7138_)
);

AOI21X1 _17803_ (
    .A(_7133_),
    .B(_7138_),
    .C(\datapath.idinstr_18_bF$buf2 ),
    .Y(_7139_)
);

OAI21X1 _17804_ (
    .A(_7139_),
    .B(_7128_),
    .C(\datapath.idinstr_19_bF$buf4 ),
    .Y(_7140_)
);

MUX2X1 _17805_ (
    .A(\datapath.registers.838[9] [26]),
    .B(\datapath.registers.838[8] [26]),
    .S(\datapath.idinstr_15_bF$buf42 ),
    .Y(_7141_)
);

NOR2X1 _17806_ (
    .A(\datapath.registers.838[11] [26]),
    .B(_5762__bF$buf17),
    .Y(_7142_)
);

OAI21X1 _17807_ (
    .A(\datapath.registers.838[10] [26]),
    .B(\datapath.idinstr_15_bF$buf41 ),
    .C(\datapath.idinstr_16_bF$buf1 ),
    .Y(_7143_)
);

OAI22X1 _17808_ (
    .A(_7143_),
    .B(_7142_),
    .C(\datapath.idinstr_16_bF$buf0 ),
    .D(_7141_),
    .Y(_7144_)
);

INVX1 _17809_ (
    .A(\datapath.registers.838[15] [26]),
    .Y(_7145_)
);

AOI21X1 _17810_ (
    .A(_5762__bF$buf16),
    .B(\datapath.registers.838[14] [26]),
    .C(_5756__bF$buf4),
    .Y(_7146_)
);

OAI21X1 _17811_ (
    .A(_7145_),
    .B(_5762__bF$buf15),
    .C(_7146_),
    .Y(_7147_)
);

NAND2X1 _17812_ (
    .A(\datapath.registers.838[12] [26]),
    .B(_5762__bF$buf14),
    .Y(_7148_)
);

AOI21X1 _17813_ (
    .A(\datapath.registers.838[13] [26]),
    .B(\datapath.idinstr_15_bF$buf40 ),
    .C(\datapath.idinstr_16_bF$buf51 ),
    .Y(_7149_)
);

AOI21X1 _17814_ (
    .A(_7148_),
    .B(_7149_),
    .C(_5757__bF$buf9),
    .Y(_7150_)
);

AOI22X1 _17815_ (
    .A(_7147_),
    .B(_7150_),
    .C(_5757__bF$buf8),
    .D(_7144_),
    .Y(_7151_)
);

NOR2X1 _17816_ (
    .A(\datapath.registers.838[0] [26]),
    .B(\datapath.idinstr_15_bF$buf39 ),
    .Y(_7152_)
);

OAI21X1 _17817_ (
    .A(\datapath.registers.838[1] [26]),
    .B(_5762__bF$buf13),
    .C(_5756__bF$buf3),
    .Y(_7153_)
);

NOR2X1 _17818_ (
    .A(\datapath.registers.838[3] [26]),
    .B(_5762__bF$buf12),
    .Y(_7154_)
);

OAI21X1 _17819_ (
    .A(\datapath.registers.838[2] [26]),
    .B(\datapath.idinstr_15_bF$buf38 ),
    .C(\datapath.idinstr_16_bF$buf50 ),
    .Y(_7155_)
);

OAI22X1 _17820_ (
    .A(_7154_),
    .B(_7155_),
    .C(_7152_),
    .D(_7153_),
    .Y(_7156_)
);

NOR2X1 _17821_ (
    .A(\datapath.idinstr_17_bF$buf1 ),
    .B(_7156_),
    .Y(_7157_)
);

MUX2X1 _17822_ (
    .A(\datapath.registers.838[5] [26]),
    .B(\datapath.registers.838[4] [26]),
    .S(\datapath.idinstr_15_bF$buf37 ),
    .Y(_7158_)
);

NOR2X1 _17823_ (
    .A(\datapath.registers.838[7] [26]),
    .B(_5762__bF$buf11),
    .Y(_7159_)
);

OAI21X1 _17824_ (
    .A(\datapath.registers.838[6] [26]),
    .B(\datapath.idinstr_15_bF$buf36 ),
    .C(\datapath.idinstr_16_bF$buf49 ),
    .Y(_7160_)
);

OAI22X1 _17825_ (
    .A(_7160_),
    .B(_7159_),
    .C(\datapath.idinstr_16_bF$buf48 ),
    .D(_7158_),
    .Y(_7161_)
);

OAI21X1 _17826_ (
    .A(_5757__bF$buf7),
    .B(_7161_),
    .C(_5760__bF$buf7),
    .Y(_7162_)
);

OAI22X1 _17827_ (
    .A(_5760__bF$buf6),
    .B(_7151_),
    .C(_7157_),
    .D(_7162_),
    .Y(_7163_)
);

NAND2X1 _17828_ (
    .A(_5789__bF$buf3),
    .B(_7163_),
    .Y(_7164_)
);

AOI22X1 _17829_ (
    .A(_5755__bF$buf3),
    .B(_5759__bF$buf3),
    .C(_7140_),
    .D(_7164_),
    .Y(\datapath.registers.rega_data [26])
);

MUX2X1 _17830_ (
    .A(\datapath.registers.838[9] [27]),
    .B(\datapath.registers.838[8] [27]),
    .S(\datapath.idinstr_15_bF$buf35 ),
    .Y(_7165_)
);

NOR2X1 _17831_ (
    .A(\datapath.registers.838[11] [27]),
    .B(_5762__bF$buf10),
    .Y(_7166_)
);

OAI21X1 _17832_ (
    .A(\datapath.registers.838[10] [27]),
    .B(\datapath.idinstr_15_bF$buf34 ),
    .C(\datapath.idinstr_16_bF$buf47 ),
    .Y(_7167_)
);

OAI22X1 _17833_ (
    .A(_7167_),
    .B(_7166_),
    .C(\datapath.idinstr_16_bF$buf46 ),
    .D(_7165_),
    .Y(_7168_)
);

INVX1 _17834_ (
    .A(\datapath.registers.838[15] [27]),
    .Y(_7169_)
);

AOI21X1 _17835_ (
    .A(_5762__bF$buf9),
    .B(\datapath.registers.838[14] [27]),
    .C(_5756__bF$buf2),
    .Y(_7170_)
);

OAI21X1 _17836_ (
    .A(_7169_),
    .B(_5762__bF$buf8),
    .C(_7170_),
    .Y(_7171_)
);

NAND2X1 _17837_ (
    .A(\datapath.registers.838[12] [27]),
    .B(_5762__bF$buf7),
    .Y(_7172_)
);

AOI21X1 _17838_ (
    .A(\datapath.registers.838[13] [27]),
    .B(\datapath.idinstr_15_bF$buf33 ),
    .C(\datapath.idinstr_16_bF$buf45 ),
    .Y(_7173_)
);

AOI21X1 _17839_ (
    .A(_7172_),
    .B(_7173_),
    .C(_5757__bF$buf6),
    .Y(_7174_)
);

AOI22X1 _17840_ (
    .A(_7171_),
    .B(_7174_),
    .C(_5757__bF$buf5),
    .D(_7168_),
    .Y(_7175_)
);

NOR2X1 _17841_ (
    .A(\datapath.registers.838[0] [27]),
    .B(\datapath.idinstr_15_bF$buf32 ),
    .Y(_7176_)
);

OAI21X1 _17842_ (
    .A(\datapath.registers.838[1] [27]),
    .B(_5762__bF$buf6),
    .C(_5756__bF$buf1),
    .Y(_7177_)
);

NOR2X1 _17843_ (
    .A(\datapath.registers.838[3] [27]),
    .B(_5762__bF$buf5),
    .Y(_7178_)
);

OAI21X1 _17844_ (
    .A(\datapath.registers.838[2] [27]),
    .B(\datapath.idinstr_15_bF$buf31 ),
    .C(\datapath.idinstr_16_bF$buf44 ),
    .Y(_7179_)
);

OAI22X1 _17845_ (
    .A(_7178_),
    .B(_7179_),
    .C(_7176_),
    .D(_7177_),
    .Y(_7180_)
);

NOR2X1 _17846_ (
    .A(\datapath.idinstr_17_bF$buf0 ),
    .B(_7180_),
    .Y(_7181_)
);

MUX2X1 _17847_ (
    .A(\datapath.registers.838[5] [27]),
    .B(\datapath.registers.838[4] [27]),
    .S(\datapath.idinstr_15_bF$buf30 ),
    .Y(_7182_)
);

NOR2X1 _17848_ (
    .A(\datapath.registers.838[7] [27]),
    .B(_5762__bF$buf4),
    .Y(_7183_)
);

OAI21X1 _17849_ (
    .A(\datapath.registers.838[6] [27]),
    .B(\datapath.idinstr_15_bF$buf29 ),
    .C(\datapath.idinstr_16_bF$buf43 ),
    .Y(_7184_)
);

OAI22X1 _17850_ (
    .A(_7184_),
    .B(_7183_),
    .C(\datapath.idinstr_16_bF$buf42 ),
    .D(_7182_),
    .Y(_7185_)
);

OAI21X1 _17851_ (
    .A(_5757__bF$buf4),
    .B(_7185_),
    .C(_5760__bF$buf5),
    .Y(_7186_)
);

OAI22X1 _17852_ (
    .A(_5760__bF$buf4),
    .B(_7175_),
    .C(_7181_),
    .D(_7186_),
    .Y(_7187_)
);

NAND2X1 _17853_ (
    .A(_5789__bF$buf2),
    .B(_7187_),
    .Y(_7188_)
);

INVX1 _17854_ (
    .A(\datapath.registers.838[19] [27]),
    .Y(_7189_)
);

AOI21X1 _17855_ (
    .A(\datapath.registers.838[23] [27]),
    .B(\datapath.idinstr_17_bF$buf15 ),
    .C(_5762__bF$buf3),
    .Y(_7190_)
);

OAI21X1 _17856_ (
    .A(_7189_),
    .B(\datapath.idinstr_17_bF$buf14 ),
    .C(_7190_),
    .Y(_7191_)
);

NAND2X1 _17857_ (
    .A(\datapath.registers.838[18] [27]),
    .B(_5757__bF$buf3),
    .Y(_7192_)
);

AOI21X1 _17858_ (
    .A(\datapath.registers.838[22] [27]),
    .B(\datapath.idinstr_17_bF$buf13 ),
    .C(\datapath.idinstr_15_bF$buf28 ),
    .Y(_7193_)
);

AOI21X1 _17859_ (
    .A(_7192_),
    .B(_7193_),
    .C(_5756__bF$buf0),
    .Y(_7194_)
);

AOI21X1 _17860_ (
    .A(\datapath.registers.838[21] [27]),
    .B(\datapath.idinstr_17_bF$buf12 ),
    .C(_5762__bF$buf2),
    .Y(_7195_)
);

OAI21X1 _17861_ (
    .A(_5009_),
    .B(\datapath.idinstr_17_bF$buf11 ),
    .C(_7195_),
    .Y(_7196_)
);

NAND2X1 _17862_ (
    .A(\datapath.registers.838[16] [27]),
    .B(_5757__bF$buf2),
    .Y(_7197_)
);

AOI21X1 _17863_ (
    .A(\datapath.registers.838[20] [27]),
    .B(\datapath.idinstr_17_bF$buf10 ),
    .C(\datapath.idinstr_15_bF$buf27 ),
    .Y(_7198_)
);

AOI21X1 _17864_ (
    .A(_7197_),
    .B(_7198_),
    .C(\datapath.idinstr_16_bF$buf41 ),
    .Y(_7199_)
);

AOI22X1 _17865_ (
    .A(_7194_),
    .B(_7191_),
    .C(_7196_),
    .D(_7199_),
    .Y(_7200_)
);

NOR2X1 _17866_ (
    .A(\datapath.registers.838[24] [27]),
    .B(\datapath.idinstr_15_bF$buf26 ),
    .Y(_7201_)
);

OAI21X1 _17867_ (
    .A(\datapath.registers.838[25] [27]),
    .B(_5762__bF$buf1),
    .C(_5756__bF$buf9),
    .Y(_7202_)
);

NOR2X1 _17868_ (
    .A(\datapath.registers.838[27] [27]),
    .B(_5762__bF$buf0),
    .Y(_7203_)
);

OAI21X1 _17869_ (
    .A(\datapath.idinstr_15_bF$buf25 ),
    .B(\datapath.registers.838[26] [27]),
    .C(\datapath.idinstr_16_bF$buf40 ),
    .Y(_7204_)
);

OAI22X1 _17870_ (
    .A(_7203_),
    .B(_7204_),
    .C(_7201_),
    .D(_7202_),
    .Y(_7205_)
);

NOR2X1 _17871_ (
    .A(\datapath.idinstr_17_bF$buf9 ),
    .B(_7205_),
    .Y(_7206_)
);

MUX2X1 _17872_ (
    .A(\datapath.registers.838[29] [27]),
    .B(\datapath.registers.838[28] [27]),
    .S(\datapath.idinstr_15_bF$buf24 ),
    .Y(_7207_)
);

NOR2X1 _17873_ (
    .A(\datapath.registers.838[31] [27]),
    .B(_5762__bF$buf47),
    .Y(_7208_)
);

OAI21X1 _17874_ (
    .A(\datapath.registers.838[30] [27]),
    .B(\datapath.idinstr_15_bF$buf23 ),
    .C(\datapath.idinstr_16_bF$buf39 ),
    .Y(_7209_)
);

OAI22X1 _17875_ (
    .A(_7209_),
    .B(_7208_),
    .C(\datapath.idinstr_16_bF$buf38 ),
    .D(_7207_),
    .Y(_7210_)
);

OAI21X1 _17876_ (
    .A(_5757__bF$buf1),
    .B(_7210_),
    .C(\datapath.idinstr_18_bF$buf1 ),
    .Y(_7211_)
);

OAI22X1 _17877_ (
    .A(\datapath.idinstr_18_bF$buf0 ),
    .B(_7200_),
    .C(_7206_),
    .D(_7211_),
    .Y(_7212_)
);

NAND2X1 _17878_ (
    .A(\datapath.idinstr_19_bF$buf3 ),
    .B(_7212_),
    .Y(_7213_)
);

AOI22X1 _17879_ (
    .A(_5755__bF$buf2),
    .B(_5759__bF$buf2),
    .C(_7213_),
    .D(_7188_),
    .Y(\datapath.registers.rega_data [27])
);

MUX2X1 _17880_ (
    .A(\datapath.registers.838[9] [28]),
    .B(\datapath.registers.838[8] [28]),
    .S(\datapath.idinstr_15_bF$buf22 ),
    .Y(_7214_)
);

NOR2X1 _17881_ (
    .A(\datapath.registers.838[11] [28]),
    .B(_5762__bF$buf46),
    .Y(_7215_)
);

OAI21X1 _17882_ (
    .A(\datapath.registers.838[10] [28]),
    .B(\datapath.idinstr_15_bF$buf21 ),
    .C(\datapath.idinstr_16_bF$buf37 ),
    .Y(_7216_)
);

OAI22X1 _17883_ (
    .A(_7216_),
    .B(_7215_),
    .C(\datapath.idinstr_16_bF$buf36 ),
    .D(_7214_),
    .Y(_7217_)
);

INVX1 _17884_ (
    .A(\datapath.registers.838[15] [28]),
    .Y(_7218_)
);

AOI21X1 _17885_ (
    .A(_5762__bF$buf45),
    .B(\datapath.registers.838[14] [28]),
    .C(_5756__bF$buf8),
    .Y(_7219_)
);

OAI21X1 _17886_ (
    .A(_7218_),
    .B(_5762__bF$buf44),
    .C(_7219_),
    .Y(_7220_)
);

NAND2X1 _17887_ (
    .A(\datapath.registers.838[12] [28]),
    .B(_5762__bF$buf43),
    .Y(_7221_)
);

AOI21X1 _17888_ (
    .A(\datapath.registers.838[13] [28]),
    .B(\datapath.idinstr_15_bF$buf20 ),
    .C(\datapath.idinstr_16_bF$buf35 ),
    .Y(_7222_)
);

AOI21X1 _17889_ (
    .A(_7221_),
    .B(_7222_),
    .C(_5757__bF$buf0),
    .Y(_7223_)
);

AOI22X1 _17890_ (
    .A(_7220_),
    .B(_7223_),
    .C(_5757__bF$buf10),
    .D(_7217_),
    .Y(_7224_)
);

NOR2X1 _17891_ (
    .A(\datapath.registers.838[0] [28]),
    .B(\datapath.idinstr_15_bF$buf19 ),
    .Y(_7225_)
);

OAI21X1 _17892_ (
    .A(\datapath.registers.838[1] [28]),
    .B(_5762__bF$buf42),
    .C(_5756__bF$buf7),
    .Y(_7226_)
);

NOR2X1 _17893_ (
    .A(\datapath.registers.838[3] [28]),
    .B(_5762__bF$buf41),
    .Y(_7227_)
);

OAI21X1 _17894_ (
    .A(\datapath.registers.838[2] [28]),
    .B(\datapath.idinstr_15_bF$buf18 ),
    .C(\datapath.idinstr_16_bF$buf34 ),
    .Y(_7228_)
);

OAI22X1 _17895_ (
    .A(_7227_),
    .B(_7228_),
    .C(_7225_),
    .D(_7226_),
    .Y(_7229_)
);

NOR2X1 _17896_ (
    .A(\datapath.idinstr_17_bF$buf8 ),
    .B(_7229_),
    .Y(_7230_)
);

MUX2X1 _17897_ (
    .A(\datapath.registers.838[5] [28]),
    .B(\datapath.registers.838[4] [28]),
    .S(\datapath.idinstr_15_bF$buf17 ),
    .Y(_7231_)
);

NOR2X1 _17898_ (
    .A(\datapath.registers.838[7] [28]),
    .B(_5762__bF$buf40),
    .Y(_7232_)
);

OAI21X1 _17899_ (
    .A(\datapath.registers.838[6] [28]),
    .B(\datapath.idinstr_15_bF$buf16 ),
    .C(\datapath.idinstr_16_bF$buf33 ),
    .Y(_7233_)
);

OAI22X1 _17900_ (
    .A(_7233_),
    .B(_7232_),
    .C(\datapath.idinstr_16_bF$buf32 ),
    .D(_7231_),
    .Y(_7234_)
);

OAI21X1 _17901_ (
    .A(_5757__bF$buf9),
    .B(_7234_),
    .C(_5760__bF$buf3),
    .Y(_7235_)
);

OAI22X1 _17902_ (
    .A(_5760__bF$buf2),
    .B(_7224_),
    .C(_7230_),
    .D(_7235_),
    .Y(_7236_)
);

NAND2X1 _17903_ (
    .A(_5789__bF$buf1),
    .B(_7236_),
    .Y(_7237_)
);

INVX1 _17904_ (
    .A(\datapath.registers.838[27] [28]),
    .Y(_7238_)
);

AOI21X1 _17905_ (
    .A(\datapath.registers.838[31] [28]),
    .B(\datapath.idinstr_17_bF$buf7 ),
    .C(_5762__bF$buf39),
    .Y(_7239_)
);

OAI21X1 _17906_ (
    .A(\datapath.idinstr_17_bF$buf6 ),
    .B(_7238_),
    .C(_7239_),
    .Y(_7240_)
);

INVX1 _17907_ (
    .A(\datapath.registers.838[26] [28]),
    .Y(_7241_)
);

AOI21X1 _17908_ (
    .A(\datapath.registers.838[30] [28]),
    .B(\datapath.idinstr_17_bF$buf5 ),
    .C(\datapath.idinstr_15_bF$buf15 ),
    .Y(_7242_)
);

OAI21X1 _17909_ (
    .A(\datapath.idinstr_17_bF$buf4 ),
    .B(_7241_),
    .C(_7242_),
    .Y(_7243_)
);

NAND3X1 _17910_ (
    .A(\datapath.idinstr_16_bF$buf31 ),
    .B(_7243_),
    .C(_7240_),
    .Y(_7244_)
);

INVX1 _17911_ (
    .A(\datapath.registers.838[25] [28]),
    .Y(_7245_)
);

AOI21X1 _17912_ (
    .A(\datapath.idinstr_17_bF$buf3 ),
    .B(\datapath.registers.838[29] [28]),
    .C(_5762__bF$buf38),
    .Y(_7246_)
);

OAI21X1 _17913_ (
    .A(\datapath.idinstr_17_bF$buf2 ),
    .B(_7245_),
    .C(_7246_),
    .Y(_7247_)
);

INVX1 _17914_ (
    .A(\datapath.registers.838[24] [28]),
    .Y(_7248_)
);

AOI21X1 _17915_ (
    .A(\datapath.idinstr_17_bF$buf1 ),
    .B(\datapath.registers.838[28] [28]),
    .C(\datapath.idinstr_15_bF$buf14 ),
    .Y(_7249_)
);

OAI21X1 _17916_ (
    .A(_7248_),
    .B(\datapath.idinstr_17_bF$buf0 ),
    .C(_7249_),
    .Y(_7250_)
);

NAND3X1 _17917_ (
    .A(_5756__bF$buf6),
    .B(_7250_),
    .C(_7247_),
    .Y(_7251_)
);

AOI21X1 _17918_ (
    .A(_7244_),
    .B(_7251_),
    .C(_5760__bF$buf1),
    .Y(_7252_)
);

MUX2X1 _17919_ (
    .A(\datapath.registers.838[18] [28]),
    .B(\datapath.registers.838[16] [28]),
    .S(\datapath.idinstr_16_bF$buf30 ),
    .Y(_7253_)
);

NAND2X1 _17920_ (
    .A(_5762__bF$buf37),
    .B(_7253_),
    .Y(_7254_)
);

MUX2X1 _17921_ (
    .A(\datapath.registers.838[19] [28]),
    .B(\datapath.registers.838[17] [28]),
    .S(\datapath.idinstr_16_bF$buf29 ),
    .Y(_7255_)
);

NAND2X1 _17922_ (
    .A(\datapath.idinstr_15_bF$buf13 ),
    .B(_7255_),
    .Y(_7256_)
);

NAND3X1 _17923_ (
    .A(_5757__bF$buf8),
    .B(_7254_),
    .C(_7256_),
    .Y(_7257_)
);

MUX2X1 _17924_ (
    .A(\datapath.registers.838[22] [28]),
    .B(\datapath.registers.838[20] [28]),
    .S(\datapath.idinstr_16_bF$buf28 ),
    .Y(_7258_)
);

NAND2X1 _17925_ (
    .A(_5762__bF$buf36),
    .B(_7258_),
    .Y(_7259_)
);

MUX2X1 _17926_ (
    .A(\datapath.registers.838[23] [28]),
    .B(\datapath.registers.838[21] [28]),
    .S(\datapath.idinstr_16_bF$buf27 ),
    .Y(_7260_)
);

NAND2X1 _17927_ (
    .A(\datapath.idinstr_15_bF$buf12 ),
    .B(_7260_),
    .Y(_7261_)
);

NAND3X1 _17928_ (
    .A(\datapath.idinstr_17_bF$buf15 ),
    .B(_7259_),
    .C(_7261_),
    .Y(_7262_)
);

AOI21X1 _17929_ (
    .A(_7257_),
    .B(_7262_),
    .C(\datapath.idinstr_18_bF$buf6 ),
    .Y(_7263_)
);

OAI21X1 _17930_ (
    .A(_7252_),
    .B(_7263_),
    .C(\datapath.idinstr_19_bF$buf2 ),
    .Y(_7264_)
);

AOI22X1 _17931_ (
    .A(_5755__bF$buf1),
    .B(_5759__bF$buf1),
    .C(_7264_),
    .D(_7237_),
    .Y(\datapath.registers.rega_data [28])
);

NAND2X1 _17932_ (
    .A(\datapath.idinstr_15_bF$buf11 ),
    .B(\datapath.registers.838[27] [29]),
    .Y(_7265_)
);

NAND2X1 _17933_ (
    .A(\datapath.registers.838[26] [29]),
    .B(_5762__bF$buf35),
    .Y(_7266_)
);

NAND3X1 _17934_ (
    .A(\datapath.idinstr_16_bF$buf26 ),
    .B(_7265_),
    .C(_7266_),
    .Y(_7267_)
);

NAND2X1 _17935_ (
    .A(\datapath.idinstr_15_bF$buf10 ),
    .B(\datapath.registers.838[25] [29]),
    .Y(_7268_)
);

AOI21X1 _17936_ (
    .A(_5762__bF$buf34),
    .B(\datapath.registers.838[24] [29]),
    .C(\datapath.idinstr_16_bF$buf25 ),
    .Y(_7269_)
);

NAND2X1 _17937_ (
    .A(_7268_),
    .B(_7269_),
    .Y(_7270_)
);

NAND3X1 _17938_ (
    .A(_5757__bF$buf7),
    .B(_7267_),
    .C(_7270_),
    .Y(_7271_)
);

NAND2X1 _17939_ (
    .A(\datapath.registers.838[31] [29]),
    .B(\datapath.idinstr_15_bF$buf9 ),
    .Y(_7272_)
);

AOI21X1 _17940_ (
    .A(_5762__bF$buf33),
    .B(\datapath.registers.838[30] [29]),
    .C(_5756__bF$buf5),
    .Y(_7273_)
);

NAND2X1 _17941_ (
    .A(_7272_),
    .B(_7273_),
    .Y(_7274_)
);

INVX1 _17942_ (
    .A(\datapath.registers.838[28] [29]),
    .Y(_7275_)
);

AOI21X1 _17943_ (
    .A(\datapath.idinstr_15_bF$buf8 ),
    .B(\datapath.registers.838[29] [29]),
    .C(\datapath.idinstr_16_bF$buf24 ),
    .Y(_7276_)
);

OAI21X1 _17944_ (
    .A(\datapath.idinstr_15_bF$buf7 ),
    .B(_7275_),
    .C(_7276_),
    .Y(_7277_)
);

NAND3X1 _17945_ (
    .A(\datapath.idinstr_17_bF$buf14 ),
    .B(_7277_),
    .C(_7274_),
    .Y(_7278_)
);

AOI21X1 _17946_ (
    .A(_7271_),
    .B(_7278_),
    .C(_5760__bF$buf0),
    .Y(_7279_)
);

MUX2X1 _17947_ (
    .A(\datapath.registers.838[18] [29]),
    .B(\datapath.registers.838[16] [29]),
    .S(\datapath.idinstr_16_bF$buf23 ),
    .Y(_7280_)
);

NAND2X1 _17948_ (
    .A(_5762__bF$buf32),
    .B(_7280_),
    .Y(_7281_)
);

MUX2X1 _17949_ (
    .A(\datapath.registers.838[19] [29]),
    .B(\datapath.registers.838[17] [29]),
    .S(\datapath.idinstr_16_bF$buf22 ),
    .Y(_7282_)
);

NAND2X1 _17950_ (
    .A(\datapath.idinstr_15_bF$buf6 ),
    .B(_7282_),
    .Y(_7283_)
);

NAND3X1 _17951_ (
    .A(_5757__bF$buf6),
    .B(_7281_),
    .C(_7283_),
    .Y(_7284_)
);

MUX2X1 _17952_ (
    .A(\datapath.registers.838[22] [29]),
    .B(\datapath.registers.838[20] [29]),
    .S(\datapath.idinstr_16_bF$buf21 ),
    .Y(_7285_)
);

NAND2X1 _17953_ (
    .A(_5762__bF$buf31),
    .B(_7285_),
    .Y(_7286_)
);

MUX2X1 _17954_ (
    .A(\datapath.registers.838[23] [29]),
    .B(\datapath.registers.838[21] [29]),
    .S(\datapath.idinstr_16_bF$buf20 ),
    .Y(_7287_)
);

NAND2X1 _17955_ (
    .A(\datapath.idinstr_15_bF$buf5 ),
    .B(_7287_),
    .Y(_7288_)
);

NAND3X1 _17956_ (
    .A(\datapath.idinstr_17_bF$buf13 ),
    .B(_7286_),
    .C(_7288_),
    .Y(_7289_)
);

AOI21X1 _17957_ (
    .A(_7284_),
    .B(_7289_),
    .C(\datapath.idinstr_18_bF$buf5 ),
    .Y(_7290_)
);

OAI21X1 _17958_ (
    .A(_7290_),
    .B(_7279_),
    .C(\datapath.idinstr_19_bF$buf1 ),
    .Y(_7291_)
);

MUX2X1 _17959_ (
    .A(\datapath.registers.838[9] [29]),
    .B(\datapath.registers.838[8] [29]),
    .S(\datapath.idinstr_15_bF$buf4 ),
    .Y(_7292_)
);

NOR2X1 _17960_ (
    .A(\datapath.registers.838[11] [29]),
    .B(_5762__bF$buf30),
    .Y(_7293_)
);

OAI21X1 _17961_ (
    .A(\datapath.registers.838[10] [29]),
    .B(\datapath.idinstr_15_bF$buf3 ),
    .C(\datapath.idinstr_16_bF$buf19 ),
    .Y(_7294_)
);

OAI22X1 _17962_ (
    .A(_7294_),
    .B(_7293_),
    .C(\datapath.idinstr_16_bF$buf18 ),
    .D(_7292_),
    .Y(_7295_)
);

INVX1 _17963_ (
    .A(\datapath.registers.838[15] [29]),
    .Y(_7296_)
);

AOI21X1 _17964_ (
    .A(_5762__bF$buf29),
    .B(\datapath.registers.838[14] [29]),
    .C(_5756__bF$buf4),
    .Y(_7297_)
);

OAI21X1 _17965_ (
    .A(_7296_),
    .B(_5762__bF$buf28),
    .C(_7297_),
    .Y(_7298_)
);

NAND2X1 _17966_ (
    .A(\datapath.registers.838[12] [29]),
    .B(_5762__bF$buf27),
    .Y(_7299_)
);

AOI21X1 _17967_ (
    .A(\datapath.registers.838[13] [29]),
    .B(\datapath.idinstr_15_bF$buf2 ),
    .C(\datapath.idinstr_16_bF$buf17 ),
    .Y(_7300_)
);

AOI21X1 _17968_ (
    .A(_7299_),
    .B(_7300_),
    .C(_5757__bF$buf5),
    .Y(_7301_)
);

AOI22X1 _17969_ (
    .A(_7298_),
    .B(_7301_),
    .C(_5757__bF$buf4),
    .D(_7295_),
    .Y(_7302_)
);

NOR2X1 _17970_ (
    .A(\datapath.registers.838[0] [29]),
    .B(\datapath.idinstr_15_bF$buf1 ),
    .Y(_7303_)
);

OAI21X1 _17971_ (
    .A(\datapath.registers.838[1] [29]),
    .B(_5762__bF$buf26),
    .C(_5756__bF$buf3),
    .Y(_7304_)
);

NOR2X1 _17972_ (
    .A(\datapath.registers.838[3] [29]),
    .B(_5762__bF$buf25),
    .Y(_7305_)
);

OAI21X1 _17973_ (
    .A(\datapath.registers.838[2] [29]),
    .B(\datapath.idinstr_15_bF$buf0 ),
    .C(\datapath.idinstr_16_bF$buf16 ),
    .Y(_7306_)
);

OAI22X1 _17974_ (
    .A(_7305_),
    .B(_7306_),
    .C(_7303_),
    .D(_7304_),
    .Y(_7307_)
);

NOR2X1 _17975_ (
    .A(\datapath.idinstr_17_bF$buf12 ),
    .B(_7307_),
    .Y(_7308_)
);

MUX2X1 _17976_ (
    .A(\datapath.registers.838[5] [29]),
    .B(\datapath.registers.838[4] [29]),
    .S(\datapath.idinstr_15_bF$buf54 ),
    .Y(_7309_)
);

NOR2X1 _17977_ (
    .A(\datapath.registers.838[7] [29]),
    .B(_5762__bF$buf24),
    .Y(_7310_)
);

OAI21X1 _17978_ (
    .A(\datapath.registers.838[6] [29]),
    .B(\datapath.idinstr_15_bF$buf53 ),
    .C(\datapath.idinstr_16_bF$buf15 ),
    .Y(_7311_)
);

OAI22X1 _17979_ (
    .A(_7311_),
    .B(_7310_),
    .C(\datapath.idinstr_16_bF$buf14 ),
    .D(_7309_),
    .Y(_7312_)
);

OAI21X1 _17980_ (
    .A(_5757__bF$buf3),
    .B(_7312_),
    .C(_5760__bF$buf7),
    .Y(_7313_)
);

OAI22X1 _17981_ (
    .A(_5760__bF$buf6),
    .B(_7302_),
    .C(_7308_),
    .D(_7313_),
    .Y(_7314_)
);

NAND2X1 _17982_ (
    .A(_5789__bF$buf0),
    .B(_7314_),
    .Y(_7315_)
);

AOI22X1 _17983_ (
    .A(_5755__bF$buf0),
    .B(_5759__bF$buf0),
    .C(_7291_),
    .D(_7315_),
    .Y(\datapath.registers.rega_data [29])
);

NAND2X1 _17984_ (
    .A(\datapath.idinstr_15_bF$buf52 ),
    .B(\datapath.registers.838[27] [30]),
    .Y(_7316_)
);

NAND2X1 _17985_ (
    .A(\datapath.registers.838[26] [30]),
    .B(_5762__bF$buf23),
    .Y(_7317_)
);

NAND3X1 _17986_ (
    .A(\datapath.idinstr_16_bF$buf13 ),
    .B(_7316_),
    .C(_7317_),
    .Y(_7318_)
);

NAND2X1 _17987_ (
    .A(\datapath.idinstr_15_bF$buf51 ),
    .B(\datapath.registers.838[25] [30]),
    .Y(_7319_)
);

AOI21X1 _17988_ (
    .A(_5762__bF$buf22),
    .B(\datapath.registers.838[24] [30]),
    .C(\datapath.idinstr_16_bF$buf12 ),
    .Y(_7320_)
);

NAND2X1 _17989_ (
    .A(_7319_),
    .B(_7320_),
    .Y(_7321_)
);

NAND3X1 _17990_ (
    .A(_5757__bF$buf2),
    .B(_7318_),
    .C(_7321_),
    .Y(_7322_)
);

NAND2X1 _17991_ (
    .A(\datapath.registers.838[31] [30]),
    .B(\datapath.idinstr_15_bF$buf50 ),
    .Y(_7323_)
);

AOI21X1 _17992_ (
    .A(_5762__bF$buf21),
    .B(\datapath.registers.838[30] [30]),
    .C(_5756__bF$buf2),
    .Y(_7324_)
);

NAND2X1 _17993_ (
    .A(_7323_),
    .B(_7324_),
    .Y(_7325_)
);

INVX1 _17994_ (
    .A(\datapath.registers.838[28] [30]),
    .Y(_7326_)
);

AOI21X1 _17995_ (
    .A(\datapath.idinstr_15_bF$buf49 ),
    .B(\datapath.registers.838[29] [30]),
    .C(\datapath.idinstr_16_bF$buf11 ),
    .Y(_7327_)
);

OAI21X1 _17996_ (
    .A(\datapath.idinstr_15_bF$buf48 ),
    .B(_7326_),
    .C(_7327_),
    .Y(_7328_)
);

NAND3X1 _17997_ (
    .A(\datapath.idinstr_17_bF$buf11 ),
    .B(_7328_),
    .C(_7325_),
    .Y(_7329_)
);

AOI21X1 _17998_ (
    .A(_7322_),
    .B(_7329_),
    .C(_5760__bF$buf5),
    .Y(_7330_)
);

MUX2X1 _17999_ (
    .A(\datapath.registers.838[18] [30]),
    .B(\datapath.registers.838[16] [30]),
    .S(\datapath.idinstr_16_bF$buf10 ),
    .Y(_7331_)
);

NAND2X1 _18000_ (
    .A(_5762__bF$buf20),
    .B(_7331_),
    .Y(_7332_)
);

MUX2X1 _18001_ (
    .A(\datapath.registers.838[19] [30]),
    .B(\datapath.registers.838[17] [30]),
    .S(\datapath.idinstr_16_bF$buf9 ),
    .Y(_7333_)
);

NAND2X1 _18002_ (
    .A(\datapath.idinstr_15_bF$buf47 ),
    .B(_7333_),
    .Y(_7334_)
);

NAND3X1 _18003_ (
    .A(_5757__bF$buf1),
    .B(_7332_),
    .C(_7334_),
    .Y(_7335_)
);

MUX2X1 _18004_ (
    .A(\datapath.registers.838[22] [30]),
    .B(\datapath.registers.838[20] [30]),
    .S(\datapath.idinstr_16_bF$buf8 ),
    .Y(_7336_)
);

NAND2X1 _18005_ (
    .A(_5762__bF$buf19),
    .B(_7336_),
    .Y(_7337_)
);

MUX2X1 _18006_ (
    .A(\datapath.registers.838[23] [30]),
    .B(\datapath.registers.838[21] [30]),
    .S(\datapath.idinstr_16_bF$buf7 ),
    .Y(_7338_)
);

NAND2X1 _18007_ (
    .A(\datapath.idinstr_15_bF$buf46 ),
    .B(_7338_),
    .Y(_7339_)
);

NAND3X1 _18008_ (
    .A(\datapath.idinstr_17_bF$buf10 ),
    .B(_7337_),
    .C(_7339_),
    .Y(_7340_)
);

AOI21X1 _18009_ (
    .A(_7335_),
    .B(_7340_),
    .C(\datapath.idinstr_18_bF$buf4 ),
    .Y(_7341_)
);

OAI21X1 _18010_ (
    .A(_7341_),
    .B(_7330_),
    .C(\datapath.idinstr_19_bF$buf0 ),
    .Y(_7342_)
);

MUX2X1 _18011_ (
    .A(\datapath.registers.838[9] [30]),
    .B(\datapath.registers.838[8] [30]),
    .S(\datapath.idinstr_15_bF$buf45 ),
    .Y(_7343_)
);

NOR2X1 _18012_ (
    .A(\datapath.registers.838[11] [30]),
    .B(_5762__bF$buf18),
    .Y(_7344_)
);

OAI21X1 _18013_ (
    .A(\datapath.registers.838[10] [30]),
    .B(\datapath.idinstr_15_bF$buf44 ),
    .C(\datapath.idinstr_16_bF$buf6 ),
    .Y(_7345_)
);

OAI22X1 _18014_ (
    .A(_7345_),
    .B(_7344_),
    .C(\datapath.idinstr_16_bF$buf5 ),
    .D(_7343_),
    .Y(_7346_)
);

INVX1 _18015_ (
    .A(\datapath.registers.838[15] [30]),
    .Y(_7347_)
);

AOI21X1 _18016_ (
    .A(_5762__bF$buf17),
    .B(\datapath.registers.838[14] [30]),
    .C(_5756__bF$buf1),
    .Y(_7348_)
);

OAI21X1 _18017_ (
    .A(_7347_),
    .B(_5762__bF$buf16),
    .C(_7348_),
    .Y(_7349_)
);

NAND2X1 _18018_ (
    .A(\datapath.registers.838[12] [30]),
    .B(_5762__bF$buf15),
    .Y(_7350_)
);

AOI21X1 _18019_ (
    .A(\datapath.registers.838[13] [30]),
    .B(\datapath.idinstr_15_bF$buf43 ),
    .C(\datapath.idinstr_16_bF$buf4 ),
    .Y(_7351_)
);

AOI21X1 _18020_ (
    .A(_7350_),
    .B(_7351_),
    .C(_5757__bF$buf0),
    .Y(_7352_)
);

AOI22X1 _18021_ (
    .A(_7349_),
    .B(_7352_),
    .C(_5757__bF$buf10),
    .D(_7346_),
    .Y(_7353_)
);

NOR2X1 _18022_ (
    .A(\datapath.registers.838[0] [30]),
    .B(\datapath.idinstr_15_bF$buf42 ),
    .Y(_7354_)
);

OAI21X1 _18023_ (
    .A(\datapath.registers.838[1] [30]),
    .B(_5762__bF$buf14),
    .C(_5756__bF$buf0),
    .Y(_7355_)
);

NOR2X1 _18024_ (
    .A(\datapath.registers.838[3] [30]),
    .B(_5762__bF$buf13),
    .Y(_7356_)
);

OAI21X1 _18025_ (
    .A(\datapath.registers.838[2] [30]),
    .B(\datapath.idinstr_15_bF$buf41 ),
    .C(\datapath.idinstr_16_bF$buf3 ),
    .Y(_7357_)
);

OAI22X1 _18026_ (
    .A(_7356_),
    .B(_7357_),
    .C(_7354_),
    .D(_7355_),
    .Y(_7358_)
);

NOR2X1 _18027_ (
    .A(\datapath.idinstr_17_bF$buf9 ),
    .B(_7358_),
    .Y(_7359_)
);

MUX2X1 _18028_ (
    .A(\datapath.registers.838[5] [30]),
    .B(\datapath.registers.838[4] [30]),
    .S(\datapath.idinstr_15_bF$buf40 ),
    .Y(_7360_)
);

NOR2X1 _18029_ (
    .A(\datapath.registers.838[7] [30]),
    .B(_5762__bF$buf12),
    .Y(_7361_)
);

OAI21X1 _18030_ (
    .A(\datapath.registers.838[6] [30]),
    .B(\datapath.idinstr_15_bF$buf39 ),
    .C(\datapath.idinstr_16_bF$buf2 ),
    .Y(_7362_)
);

OAI22X1 _18031_ (
    .A(_7362_),
    .B(_7361_),
    .C(\datapath.idinstr_16_bF$buf1 ),
    .D(_7360_),
    .Y(_7363_)
);

OAI21X1 _18032_ (
    .A(_5757__bF$buf9),
    .B(_7363_),
    .C(_5760__bF$buf4),
    .Y(_7364_)
);

OAI22X1 _18033_ (
    .A(_5760__bF$buf3),
    .B(_7353_),
    .C(_7359_),
    .D(_7364_),
    .Y(_7365_)
);

NAND2X1 _18034_ (
    .A(_5789__bF$buf4),
    .B(_7365_),
    .Y(_7366_)
);

AOI22X1 _18035_ (
    .A(_5755__bF$buf4),
    .B(_5759__bF$buf4),
    .C(_7342_),
    .D(_7366_),
    .Y(\datapath.registers.rega_data [30])
);

NAND2X1 _18036_ (
    .A(\datapath.idinstr_15_bF$buf38 ),
    .B(\datapath.registers.838[27] [31]),
    .Y(_7367_)
);

NAND2X1 _18037_ (
    .A(\datapath.registers.838[26] [31]),
    .B(_5762__bF$buf11),
    .Y(_7368_)
);

NAND3X1 _18038_ (
    .A(\datapath.idinstr_16_bF$buf0 ),
    .B(_7367_),
    .C(_7368_),
    .Y(_7369_)
);

NAND2X1 _18039_ (
    .A(\datapath.idinstr_15_bF$buf37 ),
    .B(\datapath.registers.838[25] [31]),
    .Y(_7370_)
);

AOI21X1 _18040_ (
    .A(_5762__bF$buf10),
    .B(\datapath.registers.838[24] [31]),
    .C(\datapath.idinstr_16_bF$buf51 ),
    .Y(_7371_)
);

NAND2X1 _18041_ (
    .A(_7370_),
    .B(_7371_),
    .Y(_7372_)
);

NAND3X1 _18042_ (
    .A(_5757__bF$buf8),
    .B(_7369_),
    .C(_7372_),
    .Y(_7373_)
);

NAND2X1 _18043_ (
    .A(\datapath.registers.838[31] [31]),
    .B(\datapath.idinstr_15_bF$buf36 ),
    .Y(_7374_)
);

AOI21X1 _18044_ (
    .A(_5762__bF$buf9),
    .B(\datapath.registers.838[30] [31]),
    .C(_5756__bF$buf9),
    .Y(_7375_)
);

NAND2X1 _18045_ (
    .A(_7374_),
    .B(_7375_),
    .Y(_7376_)
);

INVX1 _18046_ (
    .A(\datapath.registers.838[28] [31]),
    .Y(_7377_)
);

AOI21X1 _18047_ (
    .A(\datapath.idinstr_15_bF$buf35 ),
    .B(\datapath.registers.838[29] [31]),
    .C(\datapath.idinstr_16_bF$buf50 ),
    .Y(_7378_)
);

OAI21X1 _18048_ (
    .A(\datapath.idinstr_15_bF$buf34 ),
    .B(_7377_),
    .C(_7378_),
    .Y(_7379_)
);

NAND3X1 _18049_ (
    .A(\datapath.idinstr_17_bF$buf8 ),
    .B(_7379_),
    .C(_7376_),
    .Y(_7380_)
);

AOI21X1 _18050_ (
    .A(_7373_),
    .B(_7380_),
    .C(_5760__bF$buf2),
    .Y(_7381_)
);

MUX2X1 _18051_ (
    .A(\datapath.registers.838[18] [31]),
    .B(\datapath.registers.838[16] [31]),
    .S(\datapath.idinstr_16_bF$buf49 ),
    .Y(_7382_)
);

NAND2X1 _18052_ (
    .A(_5762__bF$buf8),
    .B(_7382_),
    .Y(_7383_)
);

MUX2X1 _18053_ (
    .A(\datapath.registers.838[19] [31]),
    .B(\datapath.registers.838[17] [31]),
    .S(\datapath.idinstr_16_bF$buf48 ),
    .Y(_7384_)
);

NAND2X1 _18054_ (
    .A(\datapath.idinstr_15_bF$buf33 ),
    .B(_7384_),
    .Y(_7385_)
);

NAND3X1 _18055_ (
    .A(_5757__bF$buf7),
    .B(_7383_),
    .C(_7385_),
    .Y(_7386_)
);

MUX2X1 _18056_ (
    .A(\datapath.registers.838[22] [31]),
    .B(\datapath.registers.838[20] [31]),
    .S(\datapath.idinstr_16_bF$buf47 ),
    .Y(_7387_)
);

NAND2X1 _18057_ (
    .A(_5762__bF$buf7),
    .B(_7387_),
    .Y(_7388_)
);

MUX2X1 _18058_ (
    .A(\datapath.registers.838[23] [31]),
    .B(\datapath.registers.838[21] [31]),
    .S(\datapath.idinstr_16_bF$buf46 ),
    .Y(_7389_)
);

NAND2X1 _18059_ (
    .A(\datapath.idinstr_15_bF$buf32 ),
    .B(_7389_),
    .Y(_7390_)
);

NAND3X1 _18060_ (
    .A(\datapath.idinstr_17_bF$buf7 ),
    .B(_7388_),
    .C(_7390_),
    .Y(_7391_)
);

AOI21X1 _18061_ (
    .A(_7386_),
    .B(_7391_),
    .C(\datapath.idinstr_18_bF$buf3 ),
    .Y(_7392_)
);

OAI21X1 _18062_ (
    .A(_7392_),
    .B(_7381_),
    .C(\datapath.idinstr_19_bF$buf5 ),
    .Y(_7393_)
);

MUX2X1 _18063_ (
    .A(\datapath.registers.838[9] [31]),
    .B(\datapath.registers.838[8] [31]),
    .S(\datapath.idinstr_15_bF$buf31 ),
    .Y(_7394_)
);

NOR2X1 _18064_ (
    .A(\datapath.registers.838[11] [31]),
    .B(_5762__bF$buf6),
    .Y(_7395_)
);

OAI21X1 _18065_ (
    .A(\datapath.registers.838[10] [31]),
    .B(\datapath.idinstr_15_bF$buf30 ),
    .C(\datapath.idinstr_16_bF$buf45 ),
    .Y(_7396_)
);

OAI22X1 _18066_ (
    .A(_7396_),
    .B(_7395_),
    .C(\datapath.idinstr_16_bF$buf44 ),
    .D(_7394_),
    .Y(_7397_)
);

INVX1 _18067_ (
    .A(\datapath.registers.838[15] [31]),
    .Y(_7398_)
);

AOI21X1 _18068_ (
    .A(_5762__bF$buf5),
    .B(\datapath.registers.838[14] [31]),
    .C(_5756__bF$buf8),
    .Y(_7399_)
);

OAI21X1 _18069_ (
    .A(_7398_),
    .B(_5762__bF$buf4),
    .C(_7399_),
    .Y(_7400_)
);

NAND2X1 _18070_ (
    .A(\datapath.registers.838[12] [31]),
    .B(_5762__bF$buf3),
    .Y(_7401_)
);

AOI21X1 _18071_ (
    .A(\datapath.registers.838[13] [31]),
    .B(\datapath.idinstr_15_bF$buf29 ),
    .C(\datapath.idinstr_16_bF$buf43 ),
    .Y(_7402_)
);

AOI21X1 _18072_ (
    .A(_7401_),
    .B(_7402_),
    .C(_5757__bF$buf6),
    .Y(_7403_)
);

AOI22X1 _18073_ (
    .A(_7400_),
    .B(_7403_),
    .C(_5757__bF$buf5),
    .D(_7397_),
    .Y(_7404_)
);

NOR2X1 _18074_ (
    .A(\datapath.registers.838[0] [31]),
    .B(\datapath.idinstr_15_bF$buf28 ),
    .Y(_7405_)
);

OAI21X1 _18075_ (
    .A(\datapath.registers.838[1] [31]),
    .B(_5762__bF$buf2),
    .C(_5756__bF$buf7),
    .Y(_7406_)
);

NOR2X1 _18076_ (
    .A(\datapath.registers.838[3] [31]),
    .B(_5762__bF$buf1),
    .Y(_7407_)
);

OAI21X1 _18077_ (
    .A(\datapath.registers.838[2] [31]),
    .B(\datapath.idinstr_15_bF$buf27 ),
    .C(\datapath.idinstr_16_bF$buf42 ),
    .Y(_7408_)
);

OAI22X1 _18078_ (
    .A(_7407_),
    .B(_7408_),
    .C(_7405_),
    .D(_7406_),
    .Y(_7409_)
);

NOR2X1 _18079_ (
    .A(\datapath.idinstr_17_bF$buf6 ),
    .B(_7409_),
    .Y(_7410_)
);

MUX2X1 _18080_ (
    .A(\datapath.registers.838[5] [31]),
    .B(\datapath.registers.838[4] [31]),
    .S(\datapath.idinstr_15_bF$buf26 ),
    .Y(_7411_)
);

NOR2X1 _18081_ (
    .A(\datapath.registers.838[7] [31]),
    .B(_5762__bF$buf0),
    .Y(_7412_)
);

OAI21X1 _18082_ (
    .A(\datapath.registers.838[6] [31]),
    .B(\datapath.idinstr_15_bF$buf25 ),
    .C(\datapath.idinstr_16_bF$buf41 ),
    .Y(_7413_)
);

OAI22X1 _18083_ (
    .A(_7413_),
    .B(_7412_),
    .C(\datapath.idinstr_16_bF$buf40 ),
    .D(_7411_),
    .Y(_7414_)
);

OAI21X1 _18084_ (
    .A(_5757__bF$buf4),
    .B(_7414_),
    .C(_5760__bF$buf1),
    .Y(_7415_)
);

OAI22X1 _18085_ (
    .A(_5760__bF$buf0),
    .B(_7404_),
    .C(_7410_),
    .D(_7415_),
    .Y(_7416_)
);

NAND2X1 _18086_ (
    .A(_5789__bF$buf3),
    .B(_7416_),
    .Y(_7417_)
);

AOI22X1 _18087_ (
    .A(_5755__bF$buf3),
    .B(_5759__bF$buf3),
    .C(_7393_),
    .D(_7417_),
    .Y(\datapath.registers.rega_data [31])
);

NOR2X1 _18088_ (
    .A(\datapath.idinstr_24_bF$buf1 ),
    .B(\datapath.idinstr_20_bF$buf49 ),
    .Y(_7418_)
);

INVX8 _18089_ (
    .A(\datapath.idinstr_21_bF$buf45 ),
    .Y(_7419_)
);

INVX8 _18090_ (
    .A(\datapath.idinstr_22_bF$buf35 ),
    .Y(_7420_)
);

NAND2X1 _18091_ (
    .A(_7419__bF$buf9),
    .B(_7420__bF$buf10),
    .Y(_7421_)
);

NOR2X1 _18092_ (
    .A(\datapath.idinstr_23_bF$buf1 ),
    .B(_7421_),
    .Y(_7422_)
);

INVX8 _18093_ (
    .A(\datapath.idinstr_23_bF$buf0 ),
    .Y(_7423_)
);

NAND2X1 _18094_ (
    .A(\datapath.registers.838[27] [0]),
    .B(\datapath.idinstr_20_bF$buf48 ),
    .Y(_7424_)
);

INVX8 _18095_ (
    .A(\datapath.idinstr_20_bF$buf47 ),
    .Y(_7425_)
);

NAND2X1 _18096_ (
    .A(\datapath.registers.838[26] [0]),
    .B(_7425__bF$buf47),
    .Y(_7426_)
);

NAND3X1 _18097_ (
    .A(\datapath.idinstr_21_bF$buf44 ),
    .B(_7424_),
    .C(_7426_),
    .Y(_7427_)
);

NAND2X1 _18098_ (
    .A(\datapath.registers.838[25] [0]),
    .B(\datapath.idinstr_20_bF$buf46 ),
    .Y(_7428_)
);

AOI21X1 _18099_ (
    .A(_7425__bF$buf46),
    .B(\datapath.registers.838[24] [0]),
    .C(\datapath.idinstr_21_bF$buf43 ),
    .Y(_7429_)
);

NAND2X1 _18100_ (
    .A(_7428_),
    .B(_7429_),
    .Y(_7430_)
);

NAND3X1 _18101_ (
    .A(_7420__bF$buf9),
    .B(_7427_),
    .C(_7430_),
    .Y(_7431_)
);

NAND2X1 _18102_ (
    .A(\datapath.registers.838[31] [0]),
    .B(\datapath.idinstr_20_bF$buf45 ),
    .Y(_7432_)
);

AOI21X1 _18103_ (
    .A(_7425__bF$buf45),
    .B(\datapath.registers.838[30] [0]),
    .C(_7419__bF$buf8),
    .Y(_7433_)
);

NAND2X1 _18104_ (
    .A(_7432_),
    .B(_7433_),
    .Y(_7434_)
);

AOI21X1 _18105_ (
    .A(\datapath.registers.838[29] [0]),
    .B(\datapath.idinstr_20_bF$buf44 ),
    .C(\datapath.idinstr_21_bF$buf42 ),
    .Y(_7435_)
);

OAI21X1 _18106_ (
    .A(_5772_),
    .B(\datapath.idinstr_20_bF$buf43 ),
    .C(_7435_),
    .Y(_7436_)
);

NAND3X1 _18107_ (
    .A(\datapath.idinstr_22_bF$buf34 ),
    .B(_7436_),
    .C(_7434_),
    .Y(_7437_)
);

AOI21X1 _18108_ (
    .A(_7431_),
    .B(_7437_),
    .C(_7423__bF$buf7),
    .Y(_7438_)
);

MUX2X1 _18109_ (
    .A(\datapath.registers.838[18] [0]),
    .B(\datapath.registers.838[16] [0]),
    .S(\datapath.idinstr_21_bF$buf41 ),
    .Y(_7439_)
);

NAND2X1 _18110_ (
    .A(_7425__bF$buf44),
    .B(_7439_),
    .Y(_7440_)
);

MUX2X1 _18111_ (
    .A(\datapath.registers.838[19] [0]),
    .B(\datapath.registers.838[17] [0]),
    .S(\datapath.idinstr_21_bF$buf40 ),
    .Y(_7441_)
);

NAND2X1 _18112_ (
    .A(\datapath.idinstr_20_bF$buf42 ),
    .B(_7441_),
    .Y(_7442_)
);

NAND3X1 _18113_ (
    .A(_7420__bF$buf8),
    .B(_7440_),
    .C(_7442_),
    .Y(_7443_)
);

MUX2X1 _18114_ (
    .A(\datapath.registers.838[22] [0]),
    .B(\datapath.registers.838[20] [0]),
    .S(\datapath.idinstr_21_bF$buf39 ),
    .Y(_7444_)
);

NAND2X1 _18115_ (
    .A(_7425__bF$buf43),
    .B(_7444_),
    .Y(_7445_)
);

MUX2X1 _18116_ (
    .A(\datapath.registers.838[23] [0]),
    .B(\datapath.registers.838[21] [0]),
    .S(\datapath.idinstr_21_bF$buf38 ),
    .Y(_7446_)
);

NAND2X1 _18117_ (
    .A(\datapath.idinstr_20_bF$buf41 ),
    .B(_7446_),
    .Y(_7447_)
);

NAND3X1 _18118_ (
    .A(\datapath.idinstr_22_bF$buf33 ),
    .B(_7445_),
    .C(_7447_),
    .Y(_7448_)
);

AOI21X1 _18119_ (
    .A(_7443_),
    .B(_7448_),
    .C(\datapath.idinstr_23_bF$buf6 ),
    .Y(_7449_)
);

OAI21X1 _18120_ (
    .A(_7449_),
    .B(_7438_),
    .C(\datapath.idinstr_24_bF$buf0 ),
    .Y(_7450_)
);

INVX8 _18121_ (
    .A(\datapath.idinstr_24_bF$buf5 ),
    .Y(_7451_)
);

MUX2X1 _18122_ (
    .A(\datapath.registers.838[9] [0]),
    .B(\datapath.registers.838[8] [0]),
    .S(\datapath.idinstr_20_bF$buf40 ),
    .Y(_7452_)
);

NOR2X1 _18123_ (
    .A(\datapath.registers.838[11] [0]),
    .B(_7425__bF$buf42),
    .Y(_7453_)
);

OAI21X1 _18124_ (
    .A(\datapath.registers.838[10] [0]),
    .B(\datapath.idinstr_20_bF$buf39 ),
    .C(\datapath.idinstr_21_bF$buf37 ),
    .Y(_7454_)
);

OAI22X1 _18125_ (
    .A(_7454_),
    .B(_7453_),
    .C(\datapath.idinstr_21_bF$buf36 ),
    .D(_7452_),
    .Y(_7455_)
);

INVX1 _18126_ (
    .A(\datapath.registers.838[15] [0]),
    .Y(_7456_)
);

AOI21X1 _18127_ (
    .A(_7425__bF$buf41),
    .B(\datapath.registers.838[14] [0]),
    .C(_7419__bF$buf7),
    .Y(_7457_)
);

OAI21X1 _18128_ (
    .A(_7456_),
    .B(_7425__bF$buf40),
    .C(_7457_),
    .Y(_7458_)
);

NAND2X1 _18129_ (
    .A(\datapath.registers.838[12] [0]),
    .B(_7425__bF$buf39),
    .Y(_7459_)
);

AOI21X1 _18130_ (
    .A(\datapath.registers.838[13] [0]),
    .B(\datapath.idinstr_20_bF$buf38 ),
    .C(\datapath.idinstr_21_bF$buf35 ),
    .Y(_7460_)
);

AOI21X1 _18131_ (
    .A(_7459_),
    .B(_7460_),
    .C(_7420__bF$buf7),
    .Y(_7461_)
);

AOI22X1 _18132_ (
    .A(_7458_),
    .B(_7461_),
    .C(_7420__bF$buf6),
    .D(_7455_),
    .Y(_7462_)
);

NOR2X1 _18133_ (
    .A(\datapath.registers.838[0] [0]),
    .B(\datapath.idinstr_20_bF$buf37 ),
    .Y(_7463_)
);

OAI21X1 _18134_ (
    .A(\datapath.registers.838[1] [0]),
    .B(_7425__bF$buf38),
    .C(_7419__bF$buf6),
    .Y(_7464_)
);

NOR2X1 _18135_ (
    .A(\datapath.registers.838[3] [0]),
    .B(_7425__bF$buf37),
    .Y(_7465_)
);

OAI21X1 _18136_ (
    .A(\datapath.registers.838[2] [0]),
    .B(\datapath.idinstr_20_bF$buf36 ),
    .C(\datapath.idinstr_21_bF$buf34 ),
    .Y(_7466_)
);

OAI22X1 _18137_ (
    .A(_7465_),
    .B(_7466_),
    .C(_7463_),
    .D(_7464_),
    .Y(_7467_)
);

NOR2X1 _18138_ (
    .A(\datapath.idinstr_22_bF$buf32 ),
    .B(_7467_),
    .Y(_7468_)
);

MUX2X1 _18139_ (
    .A(\datapath.registers.838[5] [0]),
    .B(\datapath.registers.838[4] [0]),
    .S(\datapath.idinstr_20_bF$buf35 ),
    .Y(_7469_)
);

NOR2X1 _18140_ (
    .A(\datapath.registers.838[7] [0]),
    .B(_7425__bF$buf36),
    .Y(_7470_)
);

OAI21X1 _18141_ (
    .A(\datapath.registers.838[6] [0]),
    .B(\datapath.idinstr_20_bF$buf34 ),
    .C(\datapath.idinstr_21_bF$buf33 ),
    .Y(_7471_)
);

OAI22X1 _18142_ (
    .A(_7471_),
    .B(_7470_),
    .C(\datapath.idinstr_21_bF$buf32 ),
    .D(_7469_),
    .Y(_7472_)
);

OAI21X1 _18143_ (
    .A(_7420__bF$buf5),
    .B(_7472_),
    .C(_7423__bF$buf6),
    .Y(_7473_)
);

OAI22X1 _18144_ (
    .A(_7423__bF$buf5),
    .B(_7462_),
    .C(_7468_),
    .D(_7473_),
    .Y(_7474_)
);

NAND2X1 _18145_ (
    .A(_7451__bF$buf4),
    .B(_7474_),
    .Y(_7475_)
);

AOI22X1 _18146_ (
    .A(_7418__bF$buf4),
    .B(_7422__bF$buf4),
    .C(_7450_),
    .D(_7475_),
    .Y(\datapath.registers.regb_data [0])
);

MUX2X1 _18147_ (
    .A(\datapath.registers.838[9] [1]),
    .B(\datapath.registers.838[8] [1]),
    .S(\datapath.idinstr_20_bF$buf33 ),
    .Y(_7476_)
);

NOR2X1 _18148_ (
    .A(\datapath.registers.838[11] [1]),
    .B(_7425__bF$buf35),
    .Y(_7477_)
);

OAI21X1 _18149_ (
    .A(\datapath.registers.838[10] [1]),
    .B(\datapath.idinstr_20_bF$buf32 ),
    .C(\datapath.idinstr_21_bF$buf31 ),
    .Y(_7478_)
);

OAI22X1 _18150_ (
    .A(_7478_),
    .B(_7477_),
    .C(\datapath.idinstr_21_bF$buf30 ),
    .D(_7476_),
    .Y(_7479_)
);

AOI21X1 _18151_ (
    .A(_7425__bF$buf34),
    .B(\datapath.registers.838[14] [1]),
    .C(_7419__bF$buf5),
    .Y(_7480_)
);

OAI21X1 _18152_ (
    .A(_5819_),
    .B(_7425__bF$buf33),
    .C(_7480_),
    .Y(_7481_)
);

NAND2X1 _18153_ (
    .A(\datapath.registers.838[12] [1]),
    .B(_7425__bF$buf32),
    .Y(_7482_)
);

AOI21X1 _18154_ (
    .A(\datapath.registers.838[13] [1]),
    .B(\datapath.idinstr_20_bF$buf31 ),
    .C(\datapath.idinstr_21_bF$buf29 ),
    .Y(_7483_)
);

AOI21X1 _18155_ (
    .A(_7482_),
    .B(_7483_),
    .C(_7420__bF$buf4),
    .Y(_7484_)
);

AOI22X1 _18156_ (
    .A(_7481_),
    .B(_7484_),
    .C(_7420__bF$buf3),
    .D(_7479_),
    .Y(_7485_)
);

NOR2X1 _18157_ (
    .A(\datapath.registers.838[0] [1]),
    .B(\datapath.idinstr_20_bF$buf30 ),
    .Y(_7486_)
);

OAI21X1 _18158_ (
    .A(\datapath.registers.838[1] [1]),
    .B(_7425__bF$buf31),
    .C(_7419__bF$buf4),
    .Y(_7487_)
);

NOR2X1 _18159_ (
    .A(\datapath.registers.838[3] [1]),
    .B(_7425__bF$buf30),
    .Y(_7488_)
);

OAI21X1 _18160_ (
    .A(\datapath.registers.838[2] [1]),
    .B(\datapath.idinstr_20_bF$buf29 ),
    .C(\datapath.idinstr_21_bF$buf28 ),
    .Y(_7489_)
);

OAI22X1 _18161_ (
    .A(_7488_),
    .B(_7489_),
    .C(_7486_),
    .D(_7487_),
    .Y(_7490_)
);

NOR2X1 _18162_ (
    .A(\datapath.idinstr_22_bF$buf31 ),
    .B(_7490_),
    .Y(_7491_)
);

MUX2X1 _18163_ (
    .A(\datapath.registers.838[5] [1]),
    .B(\datapath.registers.838[4] [1]),
    .S(\datapath.idinstr_20_bF$buf28 ),
    .Y(_7492_)
);

NOR2X1 _18164_ (
    .A(\datapath.registers.838[7] [1]),
    .B(_7425__bF$buf29),
    .Y(_7493_)
);

OAI21X1 _18165_ (
    .A(\datapath.registers.838[6] [1]),
    .B(\datapath.idinstr_20_bF$buf27 ),
    .C(\datapath.idinstr_21_bF$buf27 ),
    .Y(_7494_)
);

OAI22X1 _18166_ (
    .A(_7494_),
    .B(_7493_),
    .C(\datapath.idinstr_21_bF$buf26 ),
    .D(_7492_),
    .Y(_7495_)
);

OAI21X1 _18167_ (
    .A(_7420__bF$buf2),
    .B(_7495_),
    .C(_7423__bF$buf4),
    .Y(_7496_)
);

OAI22X1 _18168_ (
    .A(_7423__bF$buf3),
    .B(_7485_),
    .C(_7491_),
    .D(_7496_),
    .Y(_7497_)
);

NAND2X1 _18169_ (
    .A(_7451__bF$buf3),
    .B(_7497_),
    .Y(_7498_)
);

AOI21X1 _18170_ (
    .A(\datapath.registers.838[31] [1]),
    .B(\datapath.idinstr_22_bF$buf30 ),
    .C(_7425__bF$buf28),
    .Y(_7499_)
);

OAI21X1 _18171_ (
    .A(_5839_),
    .B(\datapath.idinstr_22_bF$buf29 ),
    .C(_7499_),
    .Y(_7500_)
);

AOI21X1 _18172_ (
    .A(\datapath.registers.838[30] [1]),
    .B(\datapath.idinstr_22_bF$buf28 ),
    .C(\datapath.idinstr_20_bF$buf26 ),
    .Y(_7501_)
);

OAI21X1 _18173_ (
    .A(_5842_),
    .B(\datapath.idinstr_22_bF$buf27 ),
    .C(_7501_),
    .Y(_7502_)
);

NAND3X1 _18174_ (
    .A(\datapath.idinstr_21_bF$buf25 ),
    .B(_7502_),
    .C(_7500_),
    .Y(_7503_)
);

AOI21X1 _18175_ (
    .A(\datapath.registers.838[29] [1]),
    .B(\datapath.idinstr_22_bF$buf26 ),
    .C(_7425__bF$buf27),
    .Y(_7504_)
);

OAI21X1 _18176_ (
    .A(_5846_),
    .B(\datapath.idinstr_22_bF$buf25 ),
    .C(_7504_),
    .Y(_7505_)
);

AOI21X1 _18177_ (
    .A(\datapath.registers.838[28] [1]),
    .B(\datapath.idinstr_22_bF$buf24 ),
    .C(\datapath.idinstr_20_bF$buf25 ),
    .Y(_7506_)
);

OAI21X1 _18178_ (
    .A(_5849_),
    .B(\datapath.idinstr_22_bF$buf23 ),
    .C(_7506_),
    .Y(_7507_)
);

NAND3X1 _18179_ (
    .A(_7419__bF$buf3),
    .B(_7507_),
    .C(_7505_),
    .Y(_7508_)
);

AOI21X1 _18180_ (
    .A(_7503_),
    .B(_7508_),
    .C(_7423__bF$buf2),
    .Y(_7509_)
);

MUX2X1 _18181_ (
    .A(\datapath.registers.838[18] [1]),
    .B(\datapath.registers.838[16] [1]),
    .S(\datapath.idinstr_21_bF$buf24 ),
    .Y(_7510_)
);

NAND2X1 _18182_ (
    .A(_7425__bF$buf26),
    .B(_7510_),
    .Y(_7511_)
);

MUX2X1 _18183_ (
    .A(\datapath.registers.838[19] [1]),
    .B(\datapath.registers.838[17] [1]),
    .S(\datapath.idinstr_21_bF$buf23 ),
    .Y(_7512_)
);

NAND2X1 _18184_ (
    .A(\datapath.idinstr_20_bF$buf24 ),
    .B(_7512_),
    .Y(_7513_)
);

NAND3X1 _18185_ (
    .A(_7420__bF$buf1),
    .B(_7511_),
    .C(_7513_),
    .Y(_7514_)
);

MUX2X1 _18186_ (
    .A(\datapath.registers.838[22] [1]),
    .B(\datapath.registers.838[20] [1]),
    .S(\datapath.idinstr_21_bF$buf22 ),
    .Y(_7515_)
);

NAND2X1 _18187_ (
    .A(_7425__bF$buf25),
    .B(_7515_),
    .Y(_7516_)
);

MUX2X1 _18188_ (
    .A(\datapath.registers.838[23] [1]),
    .B(\datapath.registers.838[21] [1]),
    .S(\datapath.idinstr_21_bF$buf21 ),
    .Y(_7517_)
);

NAND2X1 _18189_ (
    .A(\datapath.idinstr_20_bF$buf23 ),
    .B(_7517_),
    .Y(_7518_)
);

NAND3X1 _18190_ (
    .A(\datapath.idinstr_22_bF$buf22 ),
    .B(_7516_),
    .C(_7518_),
    .Y(_7519_)
);

AOI21X1 _18191_ (
    .A(_7514_),
    .B(_7519_),
    .C(\datapath.idinstr_23_bF$buf5 ),
    .Y(_7520_)
);

OAI21X1 _18192_ (
    .A(_7509_),
    .B(_7520_),
    .C(\datapath.idinstr_24_bF$buf4 ),
    .Y(_7521_)
);

AOI22X1 _18193_ (
    .A(_7418__bF$buf3),
    .B(_7422__bF$buf3),
    .C(_7521_),
    .D(_7498_),
    .Y(\datapath.registers.regb_data [1])
);

NAND2X1 _18194_ (
    .A(\datapath.registers.838[27] [2]),
    .B(\datapath.idinstr_20_bF$buf22 ),
    .Y(_7522_)
);

NAND2X1 _18195_ (
    .A(\datapath.registers.838[26] [2]),
    .B(_7425__bF$buf24),
    .Y(_7523_)
);

NAND3X1 _18196_ (
    .A(\datapath.idinstr_21_bF$buf20 ),
    .B(_7522_),
    .C(_7523_),
    .Y(_7524_)
);

NAND2X1 _18197_ (
    .A(\datapath.registers.838[25] [2]),
    .B(\datapath.idinstr_20_bF$buf21 ),
    .Y(_7525_)
);

AOI21X1 _18198_ (
    .A(_7425__bF$buf23),
    .B(\datapath.registers.838[24] [2]),
    .C(\datapath.idinstr_21_bF$buf19 ),
    .Y(_7526_)
);

NAND2X1 _18199_ (
    .A(_7525_),
    .B(_7526_),
    .Y(_7527_)
);

NAND3X1 _18200_ (
    .A(_7420__bF$buf0),
    .B(_7524_),
    .C(_7527_),
    .Y(_7528_)
);

NAND2X1 _18201_ (
    .A(\datapath.registers.838[31] [2]),
    .B(\datapath.idinstr_20_bF$buf20 ),
    .Y(_7529_)
);

AOI21X1 _18202_ (
    .A(_7425__bF$buf22),
    .B(\datapath.registers.838[30] [2]),
    .C(_7419__bF$buf2),
    .Y(_7530_)
);

NAND2X1 _18203_ (
    .A(_7529_),
    .B(_7530_),
    .Y(_7531_)
);

AOI21X1 _18204_ (
    .A(\datapath.registers.838[29] [2]),
    .B(\datapath.idinstr_20_bF$buf19 ),
    .C(\datapath.idinstr_21_bF$buf18 ),
    .Y(_7532_)
);

OAI21X1 _18205_ (
    .A(_5876_),
    .B(\datapath.idinstr_20_bF$buf18 ),
    .C(_7532_),
    .Y(_7533_)
);

NAND3X1 _18206_ (
    .A(\datapath.idinstr_22_bF$buf21 ),
    .B(_7533_),
    .C(_7531_),
    .Y(_7534_)
);

AOI21X1 _18207_ (
    .A(_7528_),
    .B(_7534_),
    .C(_7423__bF$buf1),
    .Y(_7535_)
);

MUX2X1 _18208_ (
    .A(\datapath.registers.838[18] [2]),
    .B(\datapath.registers.838[16] [2]),
    .S(\datapath.idinstr_21_bF$buf17 ),
    .Y(_7536_)
);

NAND2X1 _18209_ (
    .A(_7425__bF$buf21),
    .B(_7536_),
    .Y(_7537_)
);

MUX2X1 _18210_ (
    .A(\datapath.registers.838[19] [2]),
    .B(\datapath.registers.838[17] [2]),
    .S(\datapath.idinstr_21_bF$buf16 ),
    .Y(_7538_)
);

NAND2X1 _18211_ (
    .A(\datapath.idinstr_20_bF$buf17 ),
    .B(_7538_),
    .Y(_7539_)
);

NAND3X1 _18212_ (
    .A(_7420__bF$buf10),
    .B(_7537_),
    .C(_7539_),
    .Y(_7540_)
);

MUX2X1 _18213_ (
    .A(\datapath.registers.838[22] [2]),
    .B(\datapath.registers.838[20] [2]),
    .S(\datapath.idinstr_21_bF$buf15 ),
    .Y(_7541_)
);

NAND2X1 _18214_ (
    .A(_7425__bF$buf20),
    .B(_7541_),
    .Y(_7542_)
);

MUX2X1 _18215_ (
    .A(\datapath.registers.838[23] [2]),
    .B(\datapath.registers.838[21] [2]),
    .S(\datapath.idinstr_21_bF$buf14 ),
    .Y(_7543_)
);

NAND2X1 _18216_ (
    .A(\datapath.idinstr_20_bF$buf16 ),
    .B(_7543_),
    .Y(_7544_)
);

NAND3X1 _18217_ (
    .A(\datapath.idinstr_22_bF$buf20 ),
    .B(_7542_),
    .C(_7544_),
    .Y(_7545_)
);

AOI21X1 _18218_ (
    .A(_7540_),
    .B(_7545_),
    .C(\datapath.idinstr_23_bF$buf4 ),
    .Y(_7546_)
);

OAI21X1 _18219_ (
    .A(_7546_),
    .B(_7535_),
    .C(\datapath.idinstr_24_bF$buf3 ),
    .Y(_7547_)
);

AOI21X1 _18220_ (
    .A(\datapath.registers.838[13] [2]),
    .B(\datapath.idinstr_22_bF$buf19 ),
    .C(_7425__bF$buf19),
    .Y(_7548_)
);

OAI21X1 _18221_ (
    .A(_5267_),
    .B(\datapath.idinstr_22_bF$buf18 ),
    .C(_7548_),
    .Y(_7549_)
);

INVX1 _18222_ (
    .A(\datapath.registers.838[8] [2]),
    .Y(_7550_)
);

AOI21X1 _18223_ (
    .A(\datapath.registers.838[12] [2]),
    .B(\datapath.idinstr_22_bF$buf17 ),
    .C(\datapath.idinstr_20_bF$buf15 ),
    .Y(_7551_)
);

OAI21X1 _18224_ (
    .A(_7550_),
    .B(\datapath.idinstr_22_bF$buf16 ),
    .C(_7551_),
    .Y(_7552_)
);

NAND3X1 _18225_ (
    .A(_7419__bF$buf1),
    .B(_7552_),
    .C(_7549_),
    .Y(_7553_)
);

INVX1 _18226_ (
    .A(\datapath.registers.838[11] [2]),
    .Y(_7554_)
);

AOI21X1 _18227_ (
    .A(\datapath.registers.838[15] [2]),
    .B(\datapath.idinstr_22_bF$buf15 ),
    .C(_7425__bF$buf18),
    .Y(_7555_)
);

OAI21X1 _18228_ (
    .A(_7554_),
    .B(\datapath.idinstr_22_bF$buf14 ),
    .C(_7555_),
    .Y(_7556_)
);

AOI21X1 _18229_ (
    .A(\datapath.registers.838[14] [2]),
    .B(\datapath.idinstr_22_bF$buf13 ),
    .C(\datapath.idinstr_20_bF$buf14 ),
    .Y(_7557_)
);

OAI21X1 _18230_ (
    .A(_5223_),
    .B(\datapath.idinstr_22_bF$buf12 ),
    .C(_7557_),
    .Y(_7558_)
);

NAND3X1 _18231_ (
    .A(\datapath.idinstr_21_bF$buf13 ),
    .B(_7558_),
    .C(_7556_),
    .Y(_7559_)
);

AOI21X1 _18232_ (
    .A(_7553_),
    .B(_7559_),
    .C(_7423__bF$buf0),
    .Y(_7560_)
);

MUX2X1 _18233_ (
    .A(\datapath.registers.838[1] [2]),
    .B(\datapath.registers.838[0] [2]),
    .S(\datapath.idinstr_20_bF$buf13 ),
    .Y(_7561_)
);

NOR2X1 _18234_ (
    .A(\datapath.registers.838[3] [2]),
    .B(_7425__bF$buf17),
    .Y(_7562_)
);

OAI21X1 _18235_ (
    .A(\datapath.registers.838[2] [2]),
    .B(\datapath.idinstr_20_bF$buf12 ),
    .C(\datapath.idinstr_21_bF$buf12 ),
    .Y(_7563_)
);

OAI22X1 _18236_ (
    .A(_7563_),
    .B(_7562_),
    .C(\datapath.idinstr_21_bF$buf11 ),
    .D(_7561_),
    .Y(_7564_)
);

NAND2X1 _18237_ (
    .A(_7420__bF$buf9),
    .B(_7564_),
    .Y(_7565_)
);

MUX2X1 _18238_ (
    .A(\datapath.registers.838[5] [2]),
    .B(\datapath.registers.838[4] [2]),
    .S(\datapath.idinstr_20_bF$buf11 ),
    .Y(_7566_)
);

NOR2X1 _18239_ (
    .A(\datapath.registers.838[7] [2]),
    .B(_7425__bF$buf16),
    .Y(_7567_)
);

OAI21X1 _18240_ (
    .A(\datapath.registers.838[6] [2]),
    .B(\datapath.idinstr_20_bF$buf10 ),
    .C(\datapath.idinstr_21_bF$buf10 ),
    .Y(_7568_)
);

OAI22X1 _18241_ (
    .A(_7568_),
    .B(_7567_),
    .C(\datapath.idinstr_21_bF$buf9 ),
    .D(_7566_),
    .Y(_7569_)
);

NAND2X1 _18242_ (
    .A(\datapath.idinstr_22_bF$buf11 ),
    .B(_7569_),
    .Y(_7570_)
);

AOI21X1 _18243_ (
    .A(_7565_),
    .B(_7570_),
    .C(\datapath.idinstr_23_bF$buf3 ),
    .Y(_7571_)
);

OAI21X1 _18244_ (
    .A(_7560_),
    .B(_7571_),
    .C(_7451__bF$buf2),
    .Y(_7572_)
);

AOI22X1 _18245_ (
    .A(_7418__bF$buf2),
    .B(_7422__bF$buf2),
    .C(_7547_),
    .D(_7572_),
    .Y(\datapath.registers.regb_data [2])
);

NAND2X1 _18246_ (
    .A(\datapath.registers.838[27] [3]),
    .B(\datapath.idinstr_20_bF$buf9 ),
    .Y(_7573_)
);

NAND2X1 _18247_ (
    .A(\datapath.registers.838[26] [3]),
    .B(_7425__bF$buf15),
    .Y(_7574_)
);

NAND3X1 _18248_ (
    .A(\datapath.idinstr_21_bF$buf8 ),
    .B(_7573_),
    .C(_7574_),
    .Y(_7575_)
);

NAND2X1 _18249_ (
    .A(\datapath.registers.838[25] [3]),
    .B(\datapath.idinstr_20_bF$buf8 ),
    .Y(_7576_)
);

AOI21X1 _18250_ (
    .A(_7425__bF$buf14),
    .B(\datapath.registers.838[24] [3]),
    .C(\datapath.idinstr_21_bF$buf7 ),
    .Y(_7577_)
);

NAND2X1 _18251_ (
    .A(_7576_),
    .B(_7577_),
    .Y(_7578_)
);

NAND3X1 _18252_ (
    .A(_7420__bF$buf8),
    .B(_7575_),
    .C(_7578_),
    .Y(_7579_)
);

NAND2X1 _18253_ (
    .A(\datapath.registers.838[31] [3]),
    .B(\datapath.idinstr_20_bF$buf7 ),
    .Y(_7580_)
);

AOI21X1 _18254_ (
    .A(_7425__bF$buf13),
    .B(\datapath.registers.838[30] [3]),
    .C(_7419__bF$buf0),
    .Y(_7581_)
);

NAND2X1 _18255_ (
    .A(_7580_),
    .B(_7581_),
    .Y(_7582_)
);

INVX1 _18256_ (
    .A(\datapath.registers.838[28] [3]),
    .Y(_7583_)
);

AOI21X1 _18257_ (
    .A(\datapath.registers.838[29] [3]),
    .B(\datapath.idinstr_20_bF$buf6 ),
    .C(\datapath.idinstr_21_bF$buf6 ),
    .Y(_7584_)
);

OAI21X1 _18258_ (
    .A(_7583_),
    .B(\datapath.idinstr_20_bF$buf5 ),
    .C(_7584_),
    .Y(_7585_)
);

NAND3X1 _18259_ (
    .A(\datapath.idinstr_22_bF$buf10 ),
    .B(_7585_),
    .C(_7582_),
    .Y(_7586_)
);

AOI21X1 _18260_ (
    .A(_7579_),
    .B(_7586_),
    .C(_7423__bF$buf7),
    .Y(_7587_)
);

MUX2X1 _18261_ (
    .A(\datapath.registers.838[18] [3]),
    .B(\datapath.registers.838[16] [3]),
    .S(\datapath.idinstr_21_bF$buf5 ),
    .Y(_7588_)
);

NAND2X1 _18262_ (
    .A(_7425__bF$buf12),
    .B(_7588_),
    .Y(_7589_)
);

MUX2X1 _18263_ (
    .A(\datapath.registers.838[19] [3]),
    .B(\datapath.registers.838[17] [3]),
    .S(\datapath.idinstr_21_bF$buf4 ),
    .Y(_7590_)
);

NAND2X1 _18264_ (
    .A(\datapath.idinstr_20_bF$buf4 ),
    .B(_7590_),
    .Y(_7591_)
);

NAND3X1 _18265_ (
    .A(_7420__bF$buf7),
    .B(_7589_),
    .C(_7591_),
    .Y(_7592_)
);

MUX2X1 _18266_ (
    .A(\datapath.registers.838[22] [3]),
    .B(\datapath.registers.838[20] [3]),
    .S(\datapath.idinstr_21_bF$buf3 ),
    .Y(_7593_)
);

NAND2X1 _18267_ (
    .A(_7425__bF$buf11),
    .B(_7593_),
    .Y(_7594_)
);

MUX2X1 _18268_ (
    .A(\datapath.registers.838[23] [3]),
    .B(\datapath.registers.838[21] [3]),
    .S(\datapath.idinstr_21_bF$buf2 ),
    .Y(_7595_)
);

NAND2X1 _18269_ (
    .A(\datapath.idinstr_20_bF$buf3 ),
    .B(_7595_),
    .Y(_7596_)
);

NAND3X1 _18270_ (
    .A(\datapath.idinstr_22_bF$buf9 ),
    .B(_7594_),
    .C(_7596_),
    .Y(_7597_)
);

AOI21X1 _18271_ (
    .A(_7592_),
    .B(_7597_),
    .C(\datapath.idinstr_23_bF$buf2 ),
    .Y(_7598_)
);

OAI21X1 _18272_ (
    .A(_7598_),
    .B(_7587_),
    .C(\datapath.idinstr_24_bF$buf2 ),
    .Y(_7599_)
);

MUX2X1 _18273_ (
    .A(\datapath.registers.838[9] [3]),
    .B(\datapath.registers.838[8] [3]),
    .S(\datapath.idinstr_20_bF$buf2 ),
    .Y(_7600_)
);

NOR2X1 _18274_ (
    .A(\datapath.registers.838[11] [3]),
    .B(_7425__bF$buf10),
    .Y(_7601_)
);

OAI21X1 _18275_ (
    .A(\datapath.registers.838[10] [3]),
    .B(\datapath.idinstr_20_bF$buf1 ),
    .C(\datapath.idinstr_21_bF$buf1 ),
    .Y(_7602_)
);

OAI22X1 _18276_ (
    .A(_7602_),
    .B(_7601_),
    .C(\datapath.idinstr_21_bF$buf0 ),
    .D(_7600_),
    .Y(_7603_)
);

INVX1 _18277_ (
    .A(\datapath.registers.838[15] [3]),
    .Y(_7604_)
);

AOI21X1 _18278_ (
    .A(_7425__bF$buf9),
    .B(\datapath.registers.838[14] [3]),
    .C(_7419__bF$buf9),
    .Y(_7605_)
);

OAI21X1 _18279_ (
    .A(_7604_),
    .B(_7425__bF$buf8),
    .C(_7605_),
    .Y(_7606_)
);

NAND2X1 _18280_ (
    .A(\datapath.registers.838[12] [3]),
    .B(_7425__bF$buf7),
    .Y(_7607_)
);

AOI21X1 _18281_ (
    .A(\datapath.registers.838[13] [3]),
    .B(\datapath.idinstr_20_bF$buf0 ),
    .C(\datapath.idinstr_21_bF$buf51 ),
    .Y(_7608_)
);

AOI21X1 _18282_ (
    .A(_7607_),
    .B(_7608_),
    .C(_7420__bF$buf6),
    .Y(_7609_)
);

AOI22X1 _18283_ (
    .A(_7606_),
    .B(_7609_),
    .C(_7420__bF$buf5),
    .D(_7603_),
    .Y(_7610_)
);

NOR2X1 _18284_ (
    .A(\datapath.registers.838[0] [3]),
    .B(\datapath.idinstr_20_bF$buf55 ),
    .Y(_7611_)
);

OAI21X1 _18285_ (
    .A(\datapath.registers.838[1] [3]),
    .B(_7425__bF$buf6),
    .C(_7419__bF$buf8),
    .Y(_7612_)
);

NOR2X1 _18286_ (
    .A(\datapath.registers.838[3] [3]),
    .B(_7425__bF$buf5),
    .Y(_7613_)
);

OAI21X1 _18287_ (
    .A(\datapath.registers.838[2] [3]),
    .B(\datapath.idinstr_20_bF$buf54 ),
    .C(\datapath.idinstr_21_bF$buf50 ),
    .Y(_7614_)
);

OAI22X1 _18288_ (
    .A(_7613_),
    .B(_7614_),
    .C(_7611_),
    .D(_7612_),
    .Y(_7615_)
);

NOR2X1 _18289_ (
    .A(\datapath.idinstr_22_bF$buf8 ),
    .B(_7615_),
    .Y(_7616_)
);

MUX2X1 _18290_ (
    .A(\datapath.registers.838[5] [3]),
    .B(\datapath.registers.838[4] [3]),
    .S(\datapath.idinstr_20_bF$buf53 ),
    .Y(_7617_)
);

NOR2X1 _18291_ (
    .A(\datapath.registers.838[7] [3]),
    .B(_7425__bF$buf4),
    .Y(_7618_)
);

OAI21X1 _18292_ (
    .A(\datapath.registers.838[6] [3]),
    .B(\datapath.idinstr_20_bF$buf52 ),
    .C(\datapath.idinstr_21_bF$buf49 ),
    .Y(_7619_)
);

OAI22X1 _18293_ (
    .A(_7619_),
    .B(_7618_),
    .C(\datapath.idinstr_21_bF$buf48 ),
    .D(_7617_),
    .Y(_7620_)
);

OAI21X1 _18294_ (
    .A(_7420__bF$buf4),
    .B(_7620_),
    .C(_7423__bF$buf6),
    .Y(_7621_)
);

OAI22X1 _18295_ (
    .A(_7423__bF$buf5),
    .B(_7610_),
    .C(_7616_),
    .D(_7621_),
    .Y(_7622_)
);

NAND2X1 _18296_ (
    .A(_7451__bF$buf1),
    .B(_7622_),
    .Y(_7623_)
);

AOI22X1 _18297_ (
    .A(_7418__bF$buf1),
    .B(_7422__bF$buf1),
    .C(_7599_),
    .D(_7623_),
    .Y(\datapath.registers.regb_data [3])
);

MUX2X1 _18298_ (
    .A(\datapath.registers.838[9] [4]),
    .B(\datapath.registers.838[8] [4]),
    .S(\datapath.idinstr_20_bF$buf51 ),
    .Y(_7624_)
);

NOR2X1 _18299_ (
    .A(\datapath.registers.838[11] [4]),
    .B(_7425__bF$buf3),
    .Y(_7625_)
);

OAI21X1 _18300_ (
    .A(\datapath.registers.838[10] [4]),
    .B(\datapath.idinstr_20_bF$buf50 ),
    .C(\datapath.idinstr_21_bF$buf47 ),
    .Y(_7626_)
);

OAI22X1 _18301_ (
    .A(_7626_),
    .B(_7625_),
    .C(\datapath.idinstr_21_bF$buf46 ),
    .D(_7624_),
    .Y(_7627_)
);

AOI21X1 _18302_ (
    .A(_7425__bF$buf2),
    .B(\datapath.registers.838[14] [4]),
    .C(_7419__bF$buf7),
    .Y(_7628_)
);

OAI21X1 _18303_ (
    .A(_5998_),
    .B(_7425__bF$buf1),
    .C(_7628_),
    .Y(_7629_)
);

NAND2X1 _18304_ (
    .A(\datapath.registers.838[12] [4]),
    .B(_7425__bF$buf0),
    .Y(_7630_)
);

AOI21X1 _18305_ (
    .A(\datapath.registers.838[13] [4]),
    .B(\datapath.idinstr_20_bF$buf49 ),
    .C(\datapath.idinstr_21_bF$buf45 ),
    .Y(_7631_)
);

AOI21X1 _18306_ (
    .A(_7630_),
    .B(_7631_),
    .C(_7420__bF$buf3),
    .Y(_7632_)
);

AOI22X1 _18307_ (
    .A(_7629_),
    .B(_7632_),
    .C(_7420__bF$buf2),
    .D(_7627_),
    .Y(_7633_)
);

NOR2X1 _18308_ (
    .A(\datapath.registers.838[0] [4]),
    .B(\datapath.idinstr_20_bF$buf48 ),
    .Y(_7634_)
);

OAI21X1 _18309_ (
    .A(\datapath.registers.838[1] [4]),
    .B(_7425__bF$buf47),
    .C(_7419__bF$buf6),
    .Y(_7635_)
);

NOR2X1 _18310_ (
    .A(\datapath.registers.838[3] [4]),
    .B(_7425__bF$buf46),
    .Y(_7636_)
);

OAI21X1 _18311_ (
    .A(\datapath.registers.838[2] [4]),
    .B(\datapath.idinstr_20_bF$buf47 ),
    .C(\datapath.idinstr_21_bF$buf44 ),
    .Y(_7637_)
);

OAI22X1 _18312_ (
    .A(_7636_),
    .B(_7637_),
    .C(_7634_),
    .D(_7635_),
    .Y(_7638_)
);

NOR2X1 _18313_ (
    .A(\datapath.idinstr_22_bF$buf7 ),
    .B(_7638_),
    .Y(_7639_)
);

MUX2X1 _18314_ (
    .A(\datapath.registers.838[5] [4]),
    .B(\datapath.registers.838[4] [4]),
    .S(\datapath.idinstr_20_bF$buf46 ),
    .Y(_7640_)
);

NOR2X1 _18315_ (
    .A(\datapath.registers.838[7] [4]),
    .B(_7425__bF$buf45),
    .Y(_7641_)
);

OAI21X1 _18316_ (
    .A(\datapath.registers.838[6] [4]),
    .B(\datapath.idinstr_20_bF$buf45 ),
    .C(\datapath.idinstr_21_bF$buf43 ),
    .Y(_7642_)
);

OAI22X1 _18317_ (
    .A(_7642_),
    .B(_7641_),
    .C(\datapath.idinstr_21_bF$buf42 ),
    .D(_7640_),
    .Y(_7643_)
);

OAI21X1 _18318_ (
    .A(_7420__bF$buf1),
    .B(_7643_),
    .C(_7423__bF$buf4),
    .Y(_7644_)
);

OAI22X1 _18319_ (
    .A(_7423__bF$buf3),
    .B(_7633_),
    .C(_7639_),
    .D(_7644_),
    .Y(_7645_)
);

NAND2X1 _18320_ (
    .A(_7451__bF$buf0),
    .B(_7645_),
    .Y(_7646_)
);

INVX1 _18321_ (
    .A(\datapath.registers.838[19] [4]),
    .Y(_7647_)
);

AOI21X1 _18322_ (
    .A(\datapath.registers.838[23] [4]),
    .B(\datapath.idinstr_22_bF$buf6 ),
    .C(_7425__bF$buf44),
    .Y(_7648_)
);

OAI21X1 _18323_ (
    .A(_7647_),
    .B(\datapath.idinstr_22_bF$buf5 ),
    .C(_7648_),
    .Y(_7649_)
);

NAND2X1 _18324_ (
    .A(\datapath.registers.838[18] [4]),
    .B(_7420__bF$buf0),
    .Y(_7650_)
);

AOI21X1 _18325_ (
    .A(\datapath.registers.838[22] [4]),
    .B(\datapath.idinstr_22_bF$buf4 ),
    .C(\datapath.idinstr_20_bF$buf44 ),
    .Y(_7651_)
);

AOI21X1 _18326_ (
    .A(_7650_),
    .B(_7651_),
    .C(_7419__bF$buf5),
    .Y(_7652_)
);

AOI21X1 _18327_ (
    .A(\datapath.registers.838[21] [4]),
    .B(\datapath.idinstr_22_bF$buf3 ),
    .C(_7425__bF$buf43),
    .Y(_7653_)
);

OAI21X1 _18328_ (
    .A(_4975_),
    .B(\datapath.idinstr_22_bF$buf2 ),
    .C(_7653_),
    .Y(_7654_)
);

NAND2X1 _18329_ (
    .A(\datapath.registers.838[16] [4]),
    .B(_7420__bF$buf10),
    .Y(_7655_)
);

AOI21X1 _18330_ (
    .A(\datapath.registers.838[20] [4]),
    .B(\datapath.idinstr_22_bF$buf1 ),
    .C(\datapath.idinstr_20_bF$buf43 ),
    .Y(_7656_)
);

AOI21X1 _18331_ (
    .A(_7655_),
    .B(_7656_),
    .C(\datapath.idinstr_21_bF$buf41 ),
    .Y(_7657_)
);

AOI22X1 _18332_ (
    .A(_7652_),
    .B(_7649_),
    .C(_7654_),
    .D(_7657_),
    .Y(_7658_)
);

NOR2X1 _18333_ (
    .A(\datapath.registers.838[24] [4]),
    .B(\datapath.idinstr_20_bF$buf42 ),
    .Y(_7659_)
);

OAI21X1 _18334_ (
    .A(\datapath.registers.838[25] [4]),
    .B(_7425__bF$buf42),
    .C(_7419__bF$buf4),
    .Y(_7660_)
);

NOR2X1 _18335_ (
    .A(\datapath.registers.838[27] [4]),
    .B(_7425__bF$buf41),
    .Y(_7661_)
);

OAI21X1 _18336_ (
    .A(\datapath.registers.838[26] [4]),
    .B(\datapath.idinstr_20_bF$buf41 ),
    .C(\datapath.idinstr_21_bF$buf40 ),
    .Y(_7662_)
);

OAI22X1 _18337_ (
    .A(_7661_),
    .B(_7662_),
    .C(_7659_),
    .D(_7660_),
    .Y(_7663_)
);

NOR2X1 _18338_ (
    .A(\datapath.idinstr_22_bF$buf0 ),
    .B(_7663_),
    .Y(_7664_)
);

MUX2X1 _18339_ (
    .A(\datapath.registers.838[29] [4]),
    .B(\datapath.registers.838[28] [4]),
    .S(\datapath.idinstr_20_bF$buf40 ),
    .Y(_7665_)
);

NOR2X1 _18340_ (
    .A(\datapath.registers.838[31] [4]),
    .B(_7425__bF$buf40),
    .Y(_7666_)
);

OAI21X1 _18341_ (
    .A(\datapath.registers.838[30] [4]),
    .B(\datapath.idinstr_20_bF$buf39 ),
    .C(\datapath.idinstr_21_bF$buf39 ),
    .Y(_7667_)
);

OAI22X1 _18342_ (
    .A(_7667_),
    .B(_7666_),
    .C(\datapath.idinstr_21_bF$buf38 ),
    .D(_7665_),
    .Y(_7668_)
);

OAI21X1 _18343_ (
    .A(_7420__bF$buf9),
    .B(_7668_),
    .C(\datapath.idinstr_23_bF$buf1 ),
    .Y(_7669_)
);

OAI22X1 _18344_ (
    .A(\datapath.idinstr_23_bF$buf0 ),
    .B(_7658_),
    .C(_7664_),
    .D(_7669_),
    .Y(_7670_)
);

NAND2X1 _18345_ (
    .A(\datapath.idinstr_24_bF$buf1 ),
    .B(_7670_),
    .Y(_7671_)
);

AOI22X1 _18346_ (
    .A(_7418__bF$buf0),
    .B(_7422__bF$buf0),
    .C(_7671_),
    .D(_7646_),
    .Y(\datapath.registers.regb_data [4])
);

MUX2X1 _18347_ (
    .A(\datapath.registers.838[9] [5]),
    .B(\datapath.registers.838[8] [5]),
    .S(\datapath.idinstr_20_bF$buf38 ),
    .Y(_7672_)
);

NOR2X1 _18348_ (
    .A(\datapath.registers.838[11] [5]),
    .B(_7425__bF$buf39),
    .Y(_7673_)
);

OAI21X1 _18349_ (
    .A(\datapath.registers.838[10] [5]),
    .B(\datapath.idinstr_20_bF$buf37 ),
    .C(\datapath.idinstr_21_bF$buf37 ),
    .Y(_7674_)
);

OAI22X1 _18350_ (
    .A(_7674_),
    .B(_7673_),
    .C(\datapath.idinstr_21_bF$buf36 ),
    .D(_7672_),
    .Y(_7675_)
);

AOI21X1 _18351_ (
    .A(_7425__bF$buf38),
    .B(\datapath.registers.838[14] [5]),
    .C(_7419__bF$buf3),
    .Y(_7676_)
);

OAI21X1 _18352_ (
    .A(_6022_),
    .B(_7425__bF$buf37),
    .C(_7676_),
    .Y(_7677_)
);

NAND2X1 _18353_ (
    .A(\datapath.registers.838[12] [5]),
    .B(_7425__bF$buf36),
    .Y(_7678_)
);

AOI21X1 _18354_ (
    .A(\datapath.registers.838[13] [5]),
    .B(\datapath.idinstr_20_bF$buf36 ),
    .C(\datapath.idinstr_21_bF$buf35 ),
    .Y(_7679_)
);

AOI21X1 _18355_ (
    .A(_7678_),
    .B(_7679_),
    .C(_7420__bF$buf8),
    .Y(_7680_)
);

AOI22X1 _18356_ (
    .A(_7677_),
    .B(_7680_),
    .C(_7420__bF$buf7),
    .D(_7675_),
    .Y(_7681_)
);

NOR2X1 _18357_ (
    .A(\datapath.registers.838[0] [5]),
    .B(\datapath.idinstr_20_bF$buf35 ),
    .Y(_7682_)
);

OAI21X1 _18358_ (
    .A(\datapath.registers.838[1] [5]),
    .B(_7425__bF$buf35),
    .C(_7419__bF$buf2),
    .Y(_7683_)
);

NOR2X1 _18359_ (
    .A(\datapath.registers.838[3] [5]),
    .B(_7425__bF$buf34),
    .Y(_7684_)
);

OAI21X1 _18360_ (
    .A(\datapath.registers.838[2] [5]),
    .B(\datapath.idinstr_20_bF$buf34 ),
    .C(\datapath.idinstr_21_bF$buf34 ),
    .Y(_7685_)
);

OAI22X1 _18361_ (
    .A(_7684_),
    .B(_7685_),
    .C(_7682_),
    .D(_7683_),
    .Y(_7686_)
);

NOR2X1 _18362_ (
    .A(\datapath.idinstr_22_bF$buf41 ),
    .B(_7686_),
    .Y(_7687_)
);

MUX2X1 _18363_ (
    .A(\datapath.registers.838[5] [5]),
    .B(\datapath.registers.838[4] [5]),
    .S(\datapath.idinstr_20_bF$buf33 ),
    .Y(_7688_)
);

NOR2X1 _18364_ (
    .A(\datapath.registers.838[7] [5]),
    .B(_7425__bF$buf33),
    .Y(_7689_)
);

OAI21X1 _18365_ (
    .A(\datapath.registers.838[6] [5]),
    .B(\datapath.idinstr_20_bF$buf32 ),
    .C(\datapath.idinstr_21_bF$buf33 ),
    .Y(_7690_)
);

OAI22X1 _18366_ (
    .A(_7690_),
    .B(_7689_),
    .C(\datapath.idinstr_21_bF$buf32 ),
    .D(_7688_),
    .Y(_7691_)
);

OAI21X1 _18367_ (
    .A(_7420__bF$buf6),
    .B(_7691_),
    .C(_7423__bF$buf2),
    .Y(_7692_)
);

OAI22X1 _18368_ (
    .A(_7423__bF$buf1),
    .B(_7681_),
    .C(_7687_),
    .D(_7692_),
    .Y(_7693_)
);

NAND2X1 _18369_ (
    .A(_7451__bF$buf4),
    .B(_7693_),
    .Y(_7694_)
);

INVX1 _18370_ (
    .A(\datapath.registers.838[19] [5]),
    .Y(_7695_)
);

AOI21X1 _18371_ (
    .A(\datapath.registers.838[23] [5]),
    .B(\datapath.idinstr_22_bF$buf40 ),
    .C(_7425__bF$buf32),
    .Y(_7696_)
);

OAI21X1 _18372_ (
    .A(_7695_),
    .B(\datapath.idinstr_22_bF$buf39 ),
    .C(_7696_),
    .Y(_7697_)
);

NAND2X1 _18373_ (
    .A(\datapath.registers.838[18] [5]),
    .B(_7420__bF$buf5),
    .Y(_7698_)
);

AOI21X1 _18374_ (
    .A(\datapath.registers.838[22] [5]),
    .B(\datapath.idinstr_22_bF$buf38 ),
    .C(\datapath.idinstr_20_bF$buf31 ),
    .Y(_7699_)
);

AOI21X1 _18375_ (
    .A(_7698_),
    .B(_7699_),
    .C(_7419__bF$buf1),
    .Y(_7700_)
);

AOI21X1 _18376_ (
    .A(\datapath.registers.838[21] [5]),
    .B(\datapath.idinstr_22_bF$buf37 ),
    .C(_7425__bF$buf31),
    .Y(_7701_)
);

OAI21X1 _18377_ (
    .A(_4977_),
    .B(\datapath.idinstr_22_bF$buf36 ),
    .C(_7701_),
    .Y(_7702_)
);

NAND2X1 _18378_ (
    .A(\datapath.registers.838[16] [5]),
    .B(_7420__bF$buf4),
    .Y(_7703_)
);

AOI21X1 _18379_ (
    .A(\datapath.registers.838[20] [5]),
    .B(\datapath.idinstr_22_bF$buf35 ),
    .C(\datapath.idinstr_20_bF$buf30 ),
    .Y(_7704_)
);

AOI21X1 _18380_ (
    .A(_7703_),
    .B(_7704_),
    .C(\datapath.idinstr_21_bF$buf31 ),
    .Y(_7705_)
);

AOI22X1 _18381_ (
    .A(_7700_),
    .B(_7697_),
    .C(_7702_),
    .D(_7705_),
    .Y(_7706_)
);

NOR2X1 _18382_ (
    .A(\datapath.registers.838[24] [5]),
    .B(\datapath.idinstr_20_bF$buf29 ),
    .Y(_7707_)
);

OAI21X1 _18383_ (
    .A(\datapath.registers.838[25] [5]),
    .B(_7425__bF$buf30),
    .C(_7419__bF$buf0),
    .Y(_7708_)
);

NOR2X1 _18384_ (
    .A(\datapath.registers.838[27] [5]),
    .B(_7425__bF$buf29),
    .Y(_7709_)
);

OAI21X1 _18385_ (
    .A(\datapath.registers.838[26] [5]),
    .B(\datapath.idinstr_20_bF$buf28 ),
    .C(\datapath.idinstr_21_bF$buf30 ),
    .Y(_7710_)
);

OAI22X1 _18386_ (
    .A(_7709_),
    .B(_7710_),
    .C(_7707_),
    .D(_7708_),
    .Y(_7711_)
);

NOR2X1 _18387_ (
    .A(\datapath.idinstr_22_bF$buf34 ),
    .B(_7711_),
    .Y(_7712_)
);

MUX2X1 _18388_ (
    .A(\datapath.registers.838[29] [5]),
    .B(\datapath.registers.838[28] [5]),
    .S(\datapath.idinstr_20_bF$buf27 ),
    .Y(_7713_)
);

NOR2X1 _18389_ (
    .A(\datapath.registers.838[31] [5]),
    .B(_7425__bF$buf28),
    .Y(_7714_)
);

OAI21X1 _18390_ (
    .A(\datapath.registers.838[30] [5]),
    .B(\datapath.idinstr_20_bF$buf26 ),
    .C(\datapath.idinstr_21_bF$buf29 ),
    .Y(_7715_)
);

OAI22X1 _18391_ (
    .A(_7715_),
    .B(_7714_),
    .C(\datapath.idinstr_21_bF$buf28 ),
    .D(_7713_),
    .Y(_7716_)
);

OAI21X1 _18392_ (
    .A(_7420__bF$buf3),
    .B(_7716_),
    .C(\datapath.idinstr_23_bF$buf6 ),
    .Y(_7717_)
);

OAI22X1 _18393_ (
    .A(\datapath.idinstr_23_bF$buf5 ),
    .B(_7706_),
    .C(_7712_),
    .D(_7717_),
    .Y(_7718_)
);

NAND2X1 _18394_ (
    .A(\datapath.idinstr_24_bF$buf0 ),
    .B(_7718_),
    .Y(_7719_)
);

AOI22X1 _18395_ (
    .A(_7418__bF$buf4),
    .B(_7422__bF$buf4),
    .C(_7719_),
    .D(_7694_),
    .Y(\datapath.registers.regb_data [5])
);

MUX2X1 _18396_ (
    .A(\datapath.registers.838[2] [6]),
    .B(\datapath.registers.838[0] [6]),
    .S(\datapath.idinstr_21_bF$buf27 ),
    .Y(_7720_)
);

NAND2X1 _18397_ (
    .A(_7425__bF$buf27),
    .B(_7720_),
    .Y(_7721_)
);

MUX2X1 _18398_ (
    .A(\datapath.registers.838[3] [6]),
    .B(\datapath.registers.838[1] [6]),
    .S(\datapath.idinstr_21_bF$buf26 ),
    .Y(_7722_)
);

NAND2X1 _18399_ (
    .A(\datapath.idinstr_20_bF$buf25 ),
    .B(_7722_),
    .Y(_7723_)
);

NAND3X1 _18400_ (
    .A(_7420__bF$buf2),
    .B(_7721_),
    .C(_7723_),
    .Y(_7724_)
);

MUX2X1 _18401_ (
    .A(\datapath.registers.838[6] [6]),
    .B(\datapath.registers.838[4] [6]),
    .S(\datapath.idinstr_21_bF$buf25 ),
    .Y(_7725_)
);

NAND2X1 _18402_ (
    .A(_7425__bF$buf26),
    .B(_7725_),
    .Y(_7726_)
);

MUX2X1 _18403_ (
    .A(\datapath.registers.838[7] [6]),
    .B(\datapath.registers.838[5] [6]),
    .S(\datapath.idinstr_21_bF$buf24 ),
    .Y(_7727_)
);

NAND2X1 _18404_ (
    .A(\datapath.idinstr_20_bF$buf24 ),
    .B(_7727_),
    .Y(_7728_)
);

NAND3X1 _18405_ (
    .A(\datapath.idinstr_22_bF$buf33 ),
    .B(_7726_),
    .C(_7728_),
    .Y(_7729_)
);

AOI21X1 _18406_ (
    .A(_7724_),
    .B(_7729_),
    .C(\datapath.idinstr_23_bF$buf4 ),
    .Y(_7730_)
);

AOI21X1 _18407_ (
    .A(\datapath.registers.838[13] [6]),
    .B(\datapath.idinstr_22_bF$buf32 ),
    .C(_7425__bF$buf25),
    .Y(_7731_)
);

OAI21X1 _18408_ (
    .A(_5273_),
    .B(\datapath.idinstr_22_bF$buf31 ),
    .C(_7731_),
    .Y(_7732_)
);

AOI21X1 _18409_ (
    .A(\datapath.registers.838[12] [6]),
    .B(\datapath.idinstr_22_bF$buf30 ),
    .C(\datapath.idinstr_20_bF$buf23 ),
    .Y(_7733_)
);

OAI21X1 _18410_ (
    .A(_6082_),
    .B(\datapath.idinstr_22_bF$buf29 ),
    .C(_7733_),
    .Y(_7734_)
);

NAND3X1 _18411_ (
    .A(_7419__bF$buf9),
    .B(_7734_),
    .C(_7732_),
    .Y(_7735_)
);

AOI21X1 _18412_ (
    .A(\datapath.registers.838[15] [6]),
    .B(\datapath.idinstr_22_bF$buf28 ),
    .C(_7425__bF$buf24),
    .Y(_7736_)
);

OAI21X1 _18413_ (
    .A(_6086_),
    .B(\datapath.idinstr_22_bF$buf27 ),
    .C(_7736_),
    .Y(_7737_)
);

AOI21X1 _18414_ (
    .A(\datapath.registers.838[14] [6]),
    .B(\datapath.idinstr_22_bF$buf26 ),
    .C(\datapath.idinstr_20_bF$buf22 ),
    .Y(_7738_)
);

OAI21X1 _18415_ (
    .A(_5229_),
    .B(\datapath.idinstr_22_bF$buf25 ),
    .C(_7738_),
    .Y(_7739_)
);

NAND3X1 _18416_ (
    .A(\datapath.idinstr_21_bF$buf23 ),
    .B(_7739_),
    .C(_7737_),
    .Y(_7740_)
);

AOI21X1 _18417_ (
    .A(_7735_),
    .B(_7740_),
    .C(_7423__bF$buf0),
    .Y(_7741_)
);

OAI21X1 _18418_ (
    .A(_7741_),
    .B(_7730_),
    .C(_7451__bF$buf3),
    .Y(_7742_)
);

NOR2X1 _18419_ (
    .A(\datapath.registers.838[24] [6]),
    .B(\datapath.idinstr_20_bF$buf21 ),
    .Y(_7743_)
);

OAI21X1 _18420_ (
    .A(\datapath.registers.838[25] [6]),
    .B(_7425__bF$buf23),
    .C(_7419__bF$buf8),
    .Y(_7744_)
);

NOR2X1 _18421_ (
    .A(\datapath.registers.838[27] [6]),
    .B(_7425__bF$buf22),
    .Y(_7745_)
);

OAI21X1 _18422_ (
    .A(\datapath.registers.838[26] [6]),
    .B(\datapath.idinstr_20_bF$buf20 ),
    .C(\datapath.idinstr_21_bF$buf22 ),
    .Y(_7746_)
);

OAI22X1 _18423_ (
    .A(_7745_),
    .B(_7746_),
    .C(_7743_),
    .D(_7744_),
    .Y(_7747_)
);

NOR2X1 _18424_ (
    .A(\datapath.idinstr_22_bF$buf24 ),
    .B(_7747_),
    .Y(_7748_)
);

MUX2X1 _18425_ (
    .A(\datapath.registers.838[29] [6]),
    .B(\datapath.registers.838[28] [6]),
    .S(\datapath.idinstr_20_bF$buf19 ),
    .Y(_7749_)
);

NOR2X1 _18426_ (
    .A(\datapath.registers.838[31] [6]),
    .B(_7425__bF$buf21),
    .Y(_7750_)
);

OAI21X1 _18427_ (
    .A(\datapath.registers.838[30] [6]),
    .B(\datapath.idinstr_20_bF$buf18 ),
    .C(\datapath.idinstr_21_bF$buf21 ),
    .Y(_7751_)
);

OAI22X1 _18428_ (
    .A(_7751_),
    .B(_7750_),
    .C(\datapath.idinstr_21_bF$buf20 ),
    .D(_7749_),
    .Y(_7752_)
);

OAI21X1 _18429_ (
    .A(_7420__bF$buf1),
    .B(_7752_),
    .C(\datapath.idinstr_23_bF$buf3 ),
    .Y(_7753_)
);

AOI21X1 _18430_ (
    .A(\datapath.registers.838[23] [6]),
    .B(\datapath.idinstr_22_bF$buf23 ),
    .C(_7425__bF$buf20),
    .Y(_7754_)
);

OAI21X1 _18431_ (
    .A(_6105_),
    .B(\datapath.idinstr_22_bF$buf22 ),
    .C(_7754_),
    .Y(_7755_)
);

NAND2X1 _18432_ (
    .A(\datapath.registers.838[18] [6]),
    .B(_7420__bF$buf0),
    .Y(_7756_)
);

AOI21X1 _18433_ (
    .A(\datapath.registers.838[22] [6]),
    .B(\datapath.idinstr_22_bF$buf21 ),
    .C(\datapath.idinstr_20_bF$buf17 ),
    .Y(_7757_)
);

AOI21X1 _18434_ (
    .A(_7756_),
    .B(_7757_),
    .C(_7419__bF$buf7),
    .Y(_7758_)
);

AOI21X1 _18435_ (
    .A(\datapath.registers.838[21] [6]),
    .B(\datapath.idinstr_22_bF$buf20 ),
    .C(_7425__bF$buf19),
    .Y(_7759_)
);

OAI21X1 _18436_ (
    .A(_4979_),
    .B(\datapath.idinstr_22_bF$buf19 ),
    .C(_7759_),
    .Y(_7760_)
);

NAND2X1 _18437_ (
    .A(\datapath.registers.838[16] [6]),
    .B(_7420__bF$buf10),
    .Y(_7761_)
);

AOI21X1 _18438_ (
    .A(\datapath.registers.838[20] [6]),
    .B(\datapath.idinstr_22_bF$buf18 ),
    .C(\datapath.idinstr_20_bF$buf16 ),
    .Y(_7762_)
);

AOI21X1 _18439_ (
    .A(_7761_),
    .B(_7762_),
    .C(\datapath.idinstr_21_bF$buf19 ),
    .Y(_7763_)
);

AOI22X1 _18440_ (
    .A(_7758_),
    .B(_7755_),
    .C(_7760_),
    .D(_7763_),
    .Y(_7764_)
);

OAI22X1 _18441_ (
    .A(\datapath.idinstr_23_bF$buf2 ),
    .B(_7764_),
    .C(_7748_),
    .D(_7753_),
    .Y(_7765_)
);

NAND2X1 _18442_ (
    .A(\datapath.idinstr_24_bF$buf5 ),
    .B(_7765_),
    .Y(_7766_)
);

AOI22X1 _18443_ (
    .A(_7418__bF$buf3),
    .B(_7422__bF$buf3),
    .C(_7742_),
    .D(_7766_),
    .Y(\datapath.registers.regb_data [6])
);

NAND2X1 _18444_ (
    .A(\datapath.registers.838[27] [7]),
    .B(\datapath.idinstr_20_bF$buf15 ),
    .Y(_7767_)
);

NAND2X1 _18445_ (
    .A(\datapath.registers.838[26] [7]),
    .B(_7425__bF$buf18),
    .Y(_7768_)
);

NAND3X1 _18446_ (
    .A(\datapath.idinstr_21_bF$buf18 ),
    .B(_7767_),
    .C(_7768_),
    .Y(_7769_)
);

NAND2X1 _18447_ (
    .A(\datapath.registers.838[25] [7]),
    .B(\datapath.idinstr_20_bF$buf14 ),
    .Y(_7770_)
);

AOI21X1 _18448_ (
    .A(_7425__bF$buf17),
    .B(\datapath.registers.838[24] [7]),
    .C(\datapath.idinstr_21_bF$buf17 ),
    .Y(_7771_)
);

NAND2X1 _18449_ (
    .A(_7770_),
    .B(_7771_),
    .Y(_7772_)
);

NAND3X1 _18450_ (
    .A(_7420__bF$buf9),
    .B(_7769_),
    .C(_7772_),
    .Y(_7773_)
);

NAND2X1 _18451_ (
    .A(\datapath.registers.838[31] [7]),
    .B(\datapath.idinstr_20_bF$buf13 ),
    .Y(_7774_)
);

AOI21X1 _18452_ (
    .A(_7425__bF$buf16),
    .B(\datapath.registers.838[30] [7]),
    .C(_7419__bF$buf6),
    .Y(_7775_)
);

NAND2X1 _18453_ (
    .A(_7774_),
    .B(_7775_),
    .Y(_7776_)
);

INVX1 _18454_ (
    .A(\datapath.registers.838[28] [7]),
    .Y(_7777_)
);

AOI21X1 _18455_ (
    .A(\datapath.registers.838[29] [7]),
    .B(\datapath.idinstr_20_bF$buf12 ),
    .C(\datapath.idinstr_21_bF$buf16 ),
    .Y(_7778_)
);

OAI21X1 _18456_ (
    .A(_7777_),
    .B(\datapath.idinstr_20_bF$buf11 ),
    .C(_7778_),
    .Y(_7779_)
);

NAND3X1 _18457_ (
    .A(\datapath.idinstr_22_bF$buf17 ),
    .B(_7779_),
    .C(_7776_),
    .Y(_7780_)
);

AOI21X1 _18458_ (
    .A(_7773_),
    .B(_7780_),
    .C(_7423__bF$buf7),
    .Y(_7781_)
);

MUX2X1 _18459_ (
    .A(\datapath.registers.838[18] [7]),
    .B(\datapath.registers.838[16] [7]),
    .S(\datapath.idinstr_21_bF$buf15 ),
    .Y(_7782_)
);

NAND2X1 _18460_ (
    .A(_7425__bF$buf15),
    .B(_7782_),
    .Y(_7783_)
);

MUX2X1 _18461_ (
    .A(\datapath.registers.838[19] [7]),
    .B(\datapath.registers.838[17] [7]),
    .S(\datapath.idinstr_21_bF$buf14 ),
    .Y(_7784_)
);

NAND2X1 _18462_ (
    .A(\datapath.idinstr_20_bF$buf10 ),
    .B(_7784_),
    .Y(_7785_)
);

NAND3X1 _18463_ (
    .A(_7420__bF$buf8),
    .B(_7783_),
    .C(_7785_),
    .Y(_7786_)
);

MUX2X1 _18464_ (
    .A(\datapath.registers.838[22] [7]),
    .B(\datapath.registers.838[20] [7]),
    .S(\datapath.idinstr_21_bF$buf13 ),
    .Y(_7787_)
);

NAND2X1 _18465_ (
    .A(_7425__bF$buf14),
    .B(_7787_),
    .Y(_7788_)
);

MUX2X1 _18466_ (
    .A(\datapath.registers.838[23] [7]),
    .B(\datapath.registers.838[21] [7]),
    .S(\datapath.idinstr_21_bF$buf12 ),
    .Y(_7789_)
);

NAND2X1 _18467_ (
    .A(\datapath.idinstr_20_bF$buf9 ),
    .B(_7789_),
    .Y(_7790_)
);

NAND3X1 _18468_ (
    .A(\datapath.idinstr_22_bF$buf16 ),
    .B(_7788_),
    .C(_7790_),
    .Y(_7791_)
);

AOI21X1 _18469_ (
    .A(_7786_),
    .B(_7791_),
    .C(\datapath.idinstr_23_bF$buf1 ),
    .Y(_7792_)
);

OAI21X1 _18470_ (
    .A(_7792_),
    .B(_7781_),
    .C(\datapath.idinstr_24_bF$buf4 ),
    .Y(_7793_)
);

MUX2X1 _18471_ (
    .A(\datapath.registers.838[9] [7]),
    .B(\datapath.registers.838[8] [7]),
    .S(\datapath.idinstr_20_bF$buf8 ),
    .Y(_7794_)
);

NOR2X1 _18472_ (
    .A(\datapath.registers.838[11] [7]),
    .B(_7425__bF$buf13),
    .Y(_7795_)
);

OAI21X1 _18473_ (
    .A(\datapath.registers.838[10] [7]),
    .B(\datapath.idinstr_20_bF$buf7 ),
    .C(\datapath.idinstr_21_bF$buf11 ),
    .Y(_7796_)
);

OAI22X1 _18474_ (
    .A(_7796_),
    .B(_7795_),
    .C(\datapath.idinstr_21_bF$buf10 ),
    .D(_7794_),
    .Y(_7797_)
);

AOI21X1 _18475_ (
    .A(_7425__bF$buf12),
    .B(\datapath.registers.838[14] [7]),
    .C(_7419__bF$buf5),
    .Y(_7798_)
);

OAI21X1 _18476_ (
    .A(_6123_),
    .B(_7425__bF$buf11),
    .C(_7798_),
    .Y(_7799_)
);

NAND2X1 _18477_ (
    .A(\datapath.registers.838[12] [7]),
    .B(_7425__bF$buf10),
    .Y(_7800_)
);

AOI21X1 _18478_ (
    .A(\datapath.registers.838[13] [7]),
    .B(\datapath.idinstr_20_bF$buf6 ),
    .C(\datapath.idinstr_21_bF$buf9 ),
    .Y(_7801_)
);

AOI21X1 _18479_ (
    .A(_7800_),
    .B(_7801_),
    .C(_7420__bF$buf7),
    .Y(_7802_)
);

AOI22X1 _18480_ (
    .A(_7799_),
    .B(_7802_),
    .C(_7420__bF$buf6),
    .D(_7797_),
    .Y(_7803_)
);

NOR2X1 _18481_ (
    .A(\datapath.registers.838[0] [7]),
    .B(\datapath.idinstr_20_bF$buf5 ),
    .Y(_7804_)
);

OAI21X1 _18482_ (
    .A(\datapath.registers.838[1] [7]),
    .B(_7425__bF$buf9),
    .C(_7419__bF$buf4),
    .Y(_7805_)
);

NOR2X1 _18483_ (
    .A(\datapath.registers.838[3] [7]),
    .B(_7425__bF$buf8),
    .Y(_7806_)
);

OAI21X1 _18484_ (
    .A(\datapath.registers.838[2] [7]),
    .B(\datapath.idinstr_20_bF$buf4 ),
    .C(\datapath.idinstr_21_bF$buf8 ),
    .Y(_7807_)
);

OAI22X1 _18485_ (
    .A(_7806_),
    .B(_7807_),
    .C(_7804_),
    .D(_7805_),
    .Y(_7808_)
);

NOR2X1 _18486_ (
    .A(\datapath.idinstr_22_bF$buf15 ),
    .B(_7808_),
    .Y(_7809_)
);

MUX2X1 _18487_ (
    .A(\datapath.registers.838[5] [7]),
    .B(\datapath.registers.838[4] [7]),
    .S(\datapath.idinstr_20_bF$buf3 ),
    .Y(_7810_)
);

NOR2X1 _18488_ (
    .A(\datapath.registers.838[7] [7]),
    .B(_7425__bF$buf7),
    .Y(_7811_)
);

OAI21X1 _18489_ (
    .A(\datapath.registers.838[6] [7]),
    .B(\datapath.idinstr_20_bF$buf2 ),
    .C(\datapath.idinstr_21_bF$buf7 ),
    .Y(_7812_)
);

OAI22X1 _18490_ (
    .A(_7812_),
    .B(_7811_),
    .C(\datapath.idinstr_21_bF$buf6 ),
    .D(_7810_),
    .Y(_7813_)
);

OAI21X1 _18491_ (
    .A(_7420__bF$buf5),
    .B(_7813_),
    .C(_7423__bF$buf6),
    .Y(_7814_)
);

OAI22X1 _18492_ (
    .A(_7423__bF$buf5),
    .B(_7803_),
    .C(_7809_),
    .D(_7814_),
    .Y(_7815_)
);

NAND2X1 _18493_ (
    .A(_7451__bF$buf2),
    .B(_7815_),
    .Y(_7816_)
);

AOI22X1 _18494_ (
    .A(_7418__bF$buf2),
    .B(_7422__bF$buf2),
    .C(_7793_),
    .D(_7816_),
    .Y(\datapath.registers.regb_data [7])
);

AOI21X1 _18495_ (
    .A(\datapath.registers.838[5] [8]),
    .B(\datapath.idinstr_22_bF$buf14 ),
    .C(_7425__bF$buf6),
    .Y(_7817_)
);

OAI21X1 _18496_ (
    .A(_6212_),
    .B(\datapath.idinstr_22_bF$buf13 ),
    .C(_7817_),
    .Y(_7818_)
);

AOI21X1 _18497_ (
    .A(\datapath.registers.838[4] [8]),
    .B(\datapath.idinstr_22_bF$buf12 ),
    .C(\datapath.idinstr_20_bF$buf1 ),
    .Y(_7819_)
);

OAI21X1 _18498_ (
    .A(_6215_),
    .B(\datapath.idinstr_22_bF$buf11 ),
    .C(_7819_),
    .Y(_7820_)
);

NAND3X1 _18499_ (
    .A(_7419__bF$buf3),
    .B(_7820_),
    .C(_7818_),
    .Y(_7821_)
);

AOI21X1 _18500_ (
    .A(\datapath.registers.838[7] [8]),
    .B(\datapath.idinstr_22_bF$buf10 ),
    .C(_7425__bF$buf5),
    .Y(_7822_)
);

OAI21X1 _18501_ (
    .A(_5519_),
    .B(\datapath.idinstr_22_bF$buf9 ),
    .C(_7822_),
    .Y(_7823_)
);

AOI21X1 _18502_ (
    .A(\datapath.registers.838[6] [8]),
    .B(\datapath.idinstr_22_bF$buf8 ),
    .C(\datapath.idinstr_20_bF$buf0 ),
    .Y(_7824_)
);

OAI21X1 _18503_ (
    .A(_6221_),
    .B(\datapath.idinstr_22_bF$buf7 ),
    .C(_7824_),
    .Y(_7825_)
);

NAND3X1 _18504_ (
    .A(\datapath.idinstr_21_bF$buf5 ),
    .B(_7825_),
    .C(_7823_),
    .Y(_7826_)
);

AOI21X1 _18505_ (
    .A(_7821_),
    .B(_7826_),
    .C(\datapath.idinstr_23_bF$buf0 ),
    .Y(_7827_)
);

NAND2X1 _18506_ (
    .A(\datapath.registers.838[11] [8]),
    .B(\datapath.idinstr_21_bF$buf4 ),
    .Y(_7828_)
);

NAND2X1 _18507_ (
    .A(\datapath.registers.838[9] [8]),
    .B(_7419__bF$buf2),
    .Y(_7829_)
);

NAND3X1 _18508_ (
    .A(\datapath.idinstr_20_bF$buf55 ),
    .B(_7828_),
    .C(_7829_),
    .Y(_7830_)
);

NAND2X1 _18509_ (
    .A(\datapath.registers.838[10] [8]),
    .B(\datapath.idinstr_21_bF$buf3 ),
    .Y(_7831_)
);

AOI21X1 _18510_ (
    .A(_7419__bF$buf1),
    .B(\datapath.registers.838[8] [8]),
    .C(\datapath.idinstr_20_bF$buf54 ),
    .Y(_7832_)
);

NAND2X1 _18511_ (
    .A(_7831_),
    .B(_7832_),
    .Y(_7833_)
);

NAND3X1 _18512_ (
    .A(_7420__bF$buf4),
    .B(_7830_),
    .C(_7833_),
    .Y(_7834_)
);

NAND2X1 _18513_ (
    .A(\datapath.registers.838[15] [8]),
    .B(\datapath.idinstr_21_bF$buf2 ),
    .Y(_7835_)
);

NAND2X1 _18514_ (
    .A(\datapath.registers.838[13] [8]),
    .B(_7419__bF$buf0),
    .Y(_7836_)
);

NAND3X1 _18515_ (
    .A(\datapath.idinstr_20_bF$buf53 ),
    .B(_7835_),
    .C(_7836_),
    .Y(_7837_)
);

NAND2X1 _18516_ (
    .A(\datapath.registers.838[14] [8]),
    .B(\datapath.idinstr_21_bF$buf1 ),
    .Y(_7838_)
);

AOI21X1 _18517_ (
    .A(_7419__bF$buf9),
    .B(\datapath.registers.838[12] [8]),
    .C(\datapath.idinstr_20_bF$buf52 ),
    .Y(_7839_)
);

NAND2X1 _18518_ (
    .A(_7838_),
    .B(_7839_),
    .Y(_7840_)
);

NAND3X1 _18519_ (
    .A(\datapath.idinstr_22_bF$buf6 ),
    .B(_7837_),
    .C(_7840_),
    .Y(_7841_)
);

AOI21X1 _18520_ (
    .A(_7834_),
    .B(_7841_),
    .C(_7423__bF$buf4),
    .Y(_7842_)
);

OAI21X1 _18521_ (
    .A(_7827_),
    .B(_7842_),
    .C(_7451__bF$buf1),
    .Y(_7843_)
);

MUX2X1 _18522_ (
    .A(\datapath.registers.838[17] [8]),
    .B(\datapath.registers.838[16] [8]),
    .S(\datapath.idinstr_20_bF$buf51 ),
    .Y(_7844_)
);

NOR2X1 _18523_ (
    .A(\datapath.registers.838[19] [8]),
    .B(_7425__bF$buf4),
    .Y(_7845_)
);

OAI21X1 _18524_ (
    .A(\datapath.registers.838[18] [8]),
    .B(\datapath.idinstr_20_bF$buf50 ),
    .C(\datapath.idinstr_21_bF$buf0 ),
    .Y(_7846_)
);

OAI22X1 _18525_ (
    .A(_7846_),
    .B(_7845_),
    .C(\datapath.idinstr_21_bF$buf51 ),
    .D(_7844_),
    .Y(_7847_)
);

NAND2X1 _18526_ (
    .A(_7420__bF$buf3),
    .B(_7847_),
    .Y(_7848_)
);

MUX2X1 _18527_ (
    .A(\datapath.registers.838[21] [8]),
    .B(\datapath.registers.838[20] [8]),
    .S(\datapath.idinstr_20_bF$buf49 ),
    .Y(_7849_)
);

NOR2X1 _18528_ (
    .A(\datapath.registers.838[23] [8]),
    .B(_7425__bF$buf3),
    .Y(_7850_)
);

OAI21X1 _18529_ (
    .A(\datapath.registers.838[22] [8]),
    .B(\datapath.idinstr_20_bF$buf48 ),
    .C(\datapath.idinstr_21_bF$buf50 ),
    .Y(_7851_)
);

OAI22X1 _18530_ (
    .A(_7851_),
    .B(_7850_),
    .C(\datapath.idinstr_21_bF$buf49 ),
    .D(_7849_),
    .Y(_7852_)
);

NAND2X1 _18531_ (
    .A(\datapath.idinstr_22_bF$buf5 ),
    .B(_7852_),
    .Y(_7853_)
);

AOI21X1 _18532_ (
    .A(_7848_),
    .B(_7853_),
    .C(\datapath.idinstr_23_bF$buf6 ),
    .Y(_7854_)
);

INVX1 _18533_ (
    .A(\datapath.registers.838[27] [8]),
    .Y(_7855_)
);

AOI21X1 _18534_ (
    .A(\datapath.registers.838[31] [8]),
    .B(\datapath.idinstr_22_bF$buf4 ),
    .C(_7425__bF$buf2),
    .Y(_7856_)
);

OAI21X1 _18535_ (
    .A(_7855_),
    .B(\datapath.idinstr_22_bF$buf3 ),
    .C(_7856_),
    .Y(_7857_)
);

INVX1 _18536_ (
    .A(\datapath.registers.838[26] [8]),
    .Y(_7858_)
);

AOI21X1 _18537_ (
    .A(\datapath.registers.838[30] [8]),
    .B(\datapath.idinstr_22_bF$buf2 ),
    .C(\datapath.idinstr_20_bF$buf47 ),
    .Y(_7859_)
);

OAI21X1 _18538_ (
    .A(_7858_),
    .B(\datapath.idinstr_22_bF$buf1 ),
    .C(_7859_),
    .Y(_7860_)
);

NAND3X1 _18539_ (
    .A(\datapath.idinstr_21_bF$buf48 ),
    .B(_7860_),
    .C(_7857_),
    .Y(_7861_)
);

INVX1 _18540_ (
    .A(\datapath.registers.838[25] [8]),
    .Y(_7862_)
);

AOI21X1 _18541_ (
    .A(\datapath.registers.838[29] [8]),
    .B(\datapath.idinstr_22_bF$buf0 ),
    .C(_7425__bF$buf1),
    .Y(_7863_)
);

OAI21X1 _18542_ (
    .A(_7862_),
    .B(\datapath.idinstr_22_bF$buf41 ),
    .C(_7863_),
    .Y(_7864_)
);

INVX1 _18543_ (
    .A(\datapath.registers.838[24] [8]),
    .Y(_7865_)
);

AOI21X1 _18544_ (
    .A(\datapath.registers.838[28] [8]),
    .B(\datapath.idinstr_22_bF$buf40 ),
    .C(\datapath.idinstr_20_bF$buf46 ),
    .Y(_7866_)
);

OAI21X1 _18545_ (
    .A(_7865_),
    .B(\datapath.idinstr_22_bF$buf39 ),
    .C(_7866_),
    .Y(_7867_)
);

NAND3X1 _18546_ (
    .A(_7419__bF$buf8),
    .B(_7867_),
    .C(_7864_),
    .Y(_7868_)
);

AOI21X1 _18547_ (
    .A(_7861_),
    .B(_7868_),
    .C(_7423__bF$buf3),
    .Y(_7869_)
);

OAI21X1 _18548_ (
    .A(_7869_),
    .B(_7854_),
    .C(\datapath.idinstr_24_bF$buf3 ),
    .Y(_7870_)
);

AOI22X1 _18549_ (
    .A(_7418__bF$buf1),
    .B(_7422__bF$buf1),
    .C(_7843_),
    .D(_7870_),
    .Y(\datapath.registers.regb_data [8])
);

NAND2X1 _18550_ (
    .A(\datapath.registers.838[11] [9]),
    .B(\datapath.idinstr_21_bF$buf47 ),
    .Y(_7871_)
);

NAND2X1 _18551_ (
    .A(\datapath.registers.838[9] [9]),
    .B(_7419__bF$buf7),
    .Y(_7872_)
);

NAND3X1 _18552_ (
    .A(\datapath.idinstr_20_bF$buf45 ),
    .B(_7871_),
    .C(_7872_),
    .Y(_7873_)
);

NAND2X1 _18553_ (
    .A(\datapath.registers.838[10] [9]),
    .B(\datapath.idinstr_21_bF$buf46 ),
    .Y(_7874_)
);

AOI21X1 _18554_ (
    .A(_7419__bF$buf6),
    .B(\datapath.registers.838[8] [9]),
    .C(\datapath.idinstr_20_bF$buf44 ),
    .Y(_7875_)
);

NAND2X1 _18555_ (
    .A(_7874_),
    .B(_7875_),
    .Y(_7876_)
);

NAND3X1 _18556_ (
    .A(_7420__bF$buf2),
    .B(_7873_),
    .C(_7876_),
    .Y(_7877_)
);

NAND2X1 _18557_ (
    .A(\datapath.registers.838[15] [9]),
    .B(\datapath.idinstr_21_bF$buf45 ),
    .Y(_7878_)
);

NAND2X1 _18558_ (
    .A(\datapath.registers.838[13] [9]),
    .B(_7419__bF$buf5),
    .Y(_7879_)
);

NAND3X1 _18559_ (
    .A(\datapath.idinstr_20_bF$buf43 ),
    .B(_7878_),
    .C(_7879_),
    .Y(_7880_)
);

NAND2X1 _18560_ (
    .A(\datapath.registers.838[14] [9]),
    .B(\datapath.idinstr_21_bF$buf44 ),
    .Y(_7881_)
);

AOI21X1 _18561_ (
    .A(_7419__bF$buf4),
    .B(\datapath.registers.838[12] [9]),
    .C(\datapath.idinstr_20_bF$buf42 ),
    .Y(_7882_)
);

NAND2X1 _18562_ (
    .A(_7881_),
    .B(_7882_),
    .Y(_7883_)
);

NAND3X1 _18563_ (
    .A(\datapath.idinstr_22_bF$buf38 ),
    .B(_7880_),
    .C(_7883_),
    .Y(_7884_)
);

AOI21X1 _18564_ (
    .A(_7877_),
    .B(_7884_),
    .C(_7423__bF$buf2),
    .Y(_7885_)
);

INVX1 _18565_ (
    .A(\datapath.registers.838[1] [9]),
    .Y(_7886_)
);

AOI21X1 _18566_ (
    .A(\datapath.registers.838[5] [9]),
    .B(\datapath.idinstr_22_bF$buf37 ),
    .C(_7425__bF$buf0),
    .Y(_7887_)
);

OAI21X1 _18567_ (
    .A(_7886_),
    .B(\datapath.idinstr_22_bF$buf36 ),
    .C(_7887_),
    .Y(_7888_)
);

INVX1 _18568_ (
    .A(\datapath.registers.838[0] [9]),
    .Y(_7889_)
);

AOI21X1 _18569_ (
    .A(\datapath.registers.838[4] [9]),
    .B(\datapath.idinstr_22_bF$buf35 ),
    .C(\datapath.idinstr_20_bF$buf41 ),
    .Y(_7890_)
);

OAI21X1 _18570_ (
    .A(_7889_),
    .B(\datapath.idinstr_22_bF$buf34 ),
    .C(_7890_),
    .Y(_7891_)
);

NAND3X1 _18571_ (
    .A(_7419__bF$buf3),
    .B(_7891_),
    .C(_7888_),
    .Y(_7892_)
);

AOI21X1 _18572_ (
    .A(\datapath.registers.838[7] [9]),
    .B(\datapath.idinstr_22_bF$buf33 ),
    .C(_7425__bF$buf47),
    .Y(_7893_)
);

OAI21X1 _18573_ (
    .A(_5521_),
    .B(\datapath.idinstr_22_bF$buf32 ),
    .C(_7893_),
    .Y(_7894_)
);

INVX1 _18574_ (
    .A(\datapath.registers.838[2] [9]),
    .Y(_7895_)
);

AOI21X1 _18575_ (
    .A(\datapath.registers.838[6] [9]),
    .B(\datapath.idinstr_22_bF$buf31 ),
    .C(\datapath.idinstr_20_bF$buf40 ),
    .Y(_7896_)
);

OAI21X1 _18576_ (
    .A(_7895_),
    .B(\datapath.idinstr_22_bF$buf30 ),
    .C(_7896_),
    .Y(_7897_)
);

NAND3X1 _18577_ (
    .A(\datapath.idinstr_21_bF$buf43 ),
    .B(_7897_),
    .C(_7894_),
    .Y(_7898_)
);

AOI21X1 _18578_ (
    .A(_7892_),
    .B(_7898_),
    .C(\datapath.idinstr_23_bF$buf5 ),
    .Y(_7899_)
);

OAI21X1 _18579_ (
    .A(_7899_),
    .B(_7885_),
    .C(_7451__bF$buf0),
    .Y(_7900_)
);

INVX1 _18580_ (
    .A(\datapath.registers.838[19] [9]),
    .Y(_7901_)
);

AOI21X1 _18581_ (
    .A(\datapath.registers.838[23] [9]),
    .B(\datapath.idinstr_22_bF$buf29 ),
    .C(_7425__bF$buf46),
    .Y(_7902_)
);

OAI21X1 _18582_ (
    .A(_7901_),
    .B(\datapath.idinstr_22_bF$buf28 ),
    .C(_7902_),
    .Y(_7903_)
);

NAND2X1 _18583_ (
    .A(\datapath.registers.838[18] [9]),
    .B(_7420__bF$buf1),
    .Y(_7904_)
);

AOI21X1 _18584_ (
    .A(\datapath.registers.838[22] [9]),
    .B(\datapath.idinstr_22_bF$buf27 ),
    .C(\datapath.idinstr_20_bF$buf39 ),
    .Y(_7905_)
);

AOI21X1 _18585_ (
    .A(_7904_),
    .B(_7905_),
    .C(_7419__bF$buf2),
    .Y(_7906_)
);

AOI21X1 _18586_ (
    .A(\datapath.registers.838[21] [9]),
    .B(\datapath.idinstr_22_bF$buf26 ),
    .C(_7425__bF$buf45),
    .Y(_7907_)
);

OAI21X1 _18587_ (
    .A(_4983_),
    .B(\datapath.idinstr_22_bF$buf25 ),
    .C(_7907_),
    .Y(_7908_)
);

NAND2X1 _18588_ (
    .A(\datapath.registers.838[16] [9]),
    .B(_7420__bF$buf0),
    .Y(_7909_)
);

AOI21X1 _18589_ (
    .A(\datapath.registers.838[20] [9]),
    .B(\datapath.idinstr_22_bF$buf24 ),
    .C(\datapath.idinstr_20_bF$buf38 ),
    .Y(_7910_)
);

AOI21X1 _18590_ (
    .A(_7909_),
    .B(_7910_),
    .C(\datapath.idinstr_21_bF$buf42 ),
    .Y(_7911_)
);

AOI22X1 _18591_ (
    .A(_7906_),
    .B(_7903_),
    .C(_7908_),
    .D(_7911_),
    .Y(_7912_)
);

NOR2X1 _18592_ (
    .A(\datapath.registers.838[24] [9]),
    .B(\datapath.idinstr_20_bF$buf37 ),
    .Y(_7913_)
);

OAI21X1 _18593_ (
    .A(\datapath.registers.838[25] [9]),
    .B(_7425__bF$buf44),
    .C(_7419__bF$buf1),
    .Y(_7914_)
);

NOR2X1 _18594_ (
    .A(\datapath.registers.838[27] [9]),
    .B(_7425__bF$buf43),
    .Y(_7915_)
);

OAI21X1 _18595_ (
    .A(\datapath.registers.838[26] [9]),
    .B(\datapath.idinstr_20_bF$buf36 ),
    .C(\datapath.idinstr_21_bF$buf41 ),
    .Y(_7916_)
);

OAI22X1 _18596_ (
    .A(_7915_),
    .B(_7916_),
    .C(_7913_),
    .D(_7914_),
    .Y(_7917_)
);

NOR2X1 _18597_ (
    .A(\datapath.idinstr_22_bF$buf23 ),
    .B(_7917_),
    .Y(_7918_)
);

MUX2X1 _18598_ (
    .A(\datapath.registers.838[29] [9]),
    .B(\datapath.registers.838[28] [9]),
    .S(\datapath.idinstr_20_bF$buf35 ),
    .Y(_7919_)
);

NOR2X1 _18599_ (
    .A(\datapath.registers.838[31] [9]),
    .B(_7425__bF$buf42),
    .Y(_7920_)
);

OAI21X1 _18600_ (
    .A(\datapath.registers.838[30] [9]),
    .B(\datapath.idinstr_20_bF$buf34 ),
    .C(\datapath.idinstr_21_bF$buf40 ),
    .Y(_7921_)
);

OAI22X1 _18601_ (
    .A(_7921_),
    .B(_7920_),
    .C(\datapath.idinstr_21_bF$buf39 ),
    .D(_7919_),
    .Y(_7922_)
);

OAI21X1 _18602_ (
    .A(_7420__bF$buf10),
    .B(_7922_),
    .C(\datapath.idinstr_23_bF$buf4 ),
    .Y(_7923_)
);

OAI22X1 _18603_ (
    .A(\datapath.idinstr_23_bF$buf3 ),
    .B(_7912_),
    .C(_7918_),
    .D(_7923_),
    .Y(_7924_)
);

NAND2X1 _18604_ (
    .A(\datapath.idinstr_24_bF$buf2 ),
    .B(_7924_),
    .Y(_7925_)
);

AOI22X1 _18605_ (
    .A(_7418__bF$buf0),
    .B(_7422__bF$buf0),
    .C(_7900_),
    .D(_7925_),
    .Y(\datapath.registers.regb_data [9])
);

NAND2X1 _18606_ (
    .A(\datapath.registers.838[27] [10]),
    .B(\datapath.idinstr_20_bF$buf33 ),
    .Y(_7926_)
);

NAND2X1 _18607_ (
    .A(\datapath.registers.838[26] [10]),
    .B(_7425__bF$buf41),
    .Y(_7927_)
);

NAND3X1 _18608_ (
    .A(\datapath.idinstr_21_bF$buf38 ),
    .B(_7926_),
    .C(_7927_),
    .Y(_7928_)
);

NAND2X1 _18609_ (
    .A(\datapath.registers.838[25] [10]),
    .B(\datapath.idinstr_20_bF$buf32 ),
    .Y(_7929_)
);

AOI21X1 _18610_ (
    .A(_7425__bF$buf40),
    .B(\datapath.registers.838[24] [10]),
    .C(\datapath.idinstr_21_bF$buf37 ),
    .Y(_7930_)
);

NAND2X1 _18611_ (
    .A(_7929_),
    .B(_7930_),
    .Y(_7931_)
);

NAND3X1 _18612_ (
    .A(_7420__bF$buf9),
    .B(_7928_),
    .C(_7931_),
    .Y(_7932_)
);

NAND2X1 _18613_ (
    .A(\datapath.registers.838[31] [10]),
    .B(\datapath.idinstr_20_bF$buf31 ),
    .Y(_7933_)
);

AOI21X1 _18614_ (
    .A(_7425__bF$buf39),
    .B(\datapath.registers.838[30] [10]),
    .C(_7419__bF$buf0),
    .Y(_7934_)
);

NAND2X1 _18615_ (
    .A(_7933_),
    .B(_7934_),
    .Y(_7935_)
);

INVX1 _18616_ (
    .A(\datapath.registers.838[28] [10]),
    .Y(_7936_)
);

AOI21X1 _18617_ (
    .A(\datapath.registers.838[29] [10]),
    .B(\datapath.idinstr_20_bF$buf30 ),
    .C(\datapath.idinstr_21_bF$buf36 ),
    .Y(_7937_)
);

OAI21X1 _18618_ (
    .A(_7936_),
    .B(\datapath.idinstr_20_bF$buf29 ),
    .C(_7937_),
    .Y(_7938_)
);

NAND3X1 _18619_ (
    .A(\datapath.idinstr_22_bF$buf22 ),
    .B(_7938_),
    .C(_7935_),
    .Y(_7939_)
);

AOI21X1 _18620_ (
    .A(_7932_),
    .B(_7939_),
    .C(_7423__bF$buf1),
    .Y(_7940_)
);

MUX2X1 _18621_ (
    .A(\datapath.registers.838[18] [10]),
    .B(\datapath.registers.838[16] [10]),
    .S(\datapath.idinstr_21_bF$buf35 ),
    .Y(_7941_)
);

NAND2X1 _18622_ (
    .A(_7425__bF$buf38),
    .B(_7941_),
    .Y(_7942_)
);

MUX2X1 _18623_ (
    .A(\datapath.registers.838[19] [10]),
    .B(\datapath.registers.838[17] [10]),
    .S(\datapath.idinstr_21_bF$buf34 ),
    .Y(_7943_)
);

NAND2X1 _18624_ (
    .A(\datapath.idinstr_20_bF$buf28 ),
    .B(_7943_),
    .Y(_7944_)
);

NAND3X1 _18625_ (
    .A(_7420__bF$buf8),
    .B(_7942_),
    .C(_7944_),
    .Y(_7945_)
);

MUX2X1 _18626_ (
    .A(\datapath.registers.838[22] [10]),
    .B(\datapath.registers.838[20] [10]),
    .S(\datapath.idinstr_21_bF$buf33 ),
    .Y(_7946_)
);

NAND2X1 _18627_ (
    .A(_7425__bF$buf37),
    .B(_7946_),
    .Y(_7947_)
);

MUX2X1 _18628_ (
    .A(\datapath.registers.838[23] [10]),
    .B(\datapath.registers.838[21] [10]),
    .S(\datapath.idinstr_21_bF$buf32 ),
    .Y(_7948_)
);

NAND2X1 _18629_ (
    .A(\datapath.idinstr_20_bF$buf27 ),
    .B(_7948_),
    .Y(_7949_)
);

NAND3X1 _18630_ (
    .A(\datapath.idinstr_22_bF$buf21 ),
    .B(_7947_),
    .C(_7949_),
    .Y(_7950_)
);

AOI21X1 _18631_ (
    .A(_7945_),
    .B(_7950_),
    .C(\datapath.idinstr_23_bF$buf2 ),
    .Y(_7951_)
);

OAI21X1 _18632_ (
    .A(_7951_),
    .B(_7940_),
    .C(\datapath.idinstr_24_bF$buf1 ),
    .Y(_7952_)
);

MUX2X1 _18633_ (
    .A(\datapath.registers.838[9] [10]),
    .B(\datapath.registers.838[8] [10]),
    .S(\datapath.idinstr_20_bF$buf26 ),
    .Y(_7953_)
);

NOR2X1 _18634_ (
    .A(\datapath.registers.838[11] [10]),
    .B(_7425__bF$buf36),
    .Y(_7954_)
);

OAI21X1 _18635_ (
    .A(\datapath.registers.838[10] [10]),
    .B(\datapath.idinstr_20_bF$buf25 ),
    .C(\datapath.idinstr_21_bF$buf31 ),
    .Y(_7955_)
);

OAI22X1 _18636_ (
    .A(_7955_),
    .B(_7954_),
    .C(\datapath.idinstr_21_bF$buf30 ),
    .D(_7953_),
    .Y(_7956_)
);

INVX1 _18637_ (
    .A(\datapath.registers.838[15] [10]),
    .Y(_7957_)
);

AOI21X1 _18638_ (
    .A(_7425__bF$buf35),
    .B(\datapath.registers.838[14] [10]),
    .C(_7419__bF$buf9),
    .Y(_7958_)
);

OAI21X1 _18639_ (
    .A(_7957_),
    .B(_7425__bF$buf34),
    .C(_7958_),
    .Y(_7959_)
);

NAND2X1 _18640_ (
    .A(\datapath.registers.838[12] [10]),
    .B(_7425__bF$buf33),
    .Y(_7960_)
);

AOI21X1 _18641_ (
    .A(\datapath.registers.838[13] [10]),
    .B(\datapath.idinstr_20_bF$buf24 ),
    .C(\datapath.idinstr_21_bF$buf29 ),
    .Y(_7961_)
);

AOI21X1 _18642_ (
    .A(_7960_),
    .B(_7961_),
    .C(_7420__bF$buf7),
    .Y(_7962_)
);

AOI22X1 _18643_ (
    .A(_7959_),
    .B(_7962_),
    .C(_7420__bF$buf6),
    .D(_7956_),
    .Y(_7963_)
);

NOR2X1 _18644_ (
    .A(\datapath.registers.838[0] [10]),
    .B(\datapath.idinstr_20_bF$buf23 ),
    .Y(_7964_)
);

OAI21X1 _18645_ (
    .A(\datapath.registers.838[1] [10]),
    .B(_7425__bF$buf32),
    .C(_7419__bF$buf8),
    .Y(_7965_)
);

NOR2X1 _18646_ (
    .A(\datapath.registers.838[3] [10]),
    .B(_7425__bF$buf31),
    .Y(_7966_)
);

OAI21X1 _18647_ (
    .A(\datapath.registers.838[2] [10]),
    .B(\datapath.idinstr_20_bF$buf22 ),
    .C(\datapath.idinstr_21_bF$buf28 ),
    .Y(_7967_)
);

OAI22X1 _18648_ (
    .A(_7966_),
    .B(_7967_),
    .C(_7964_),
    .D(_7965_),
    .Y(_7968_)
);

NOR2X1 _18649_ (
    .A(\datapath.idinstr_22_bF$buf20 ),
    .B(_7968_),
    .Y(_7969_)
);

MUX2X1 _18650_ (
    .A(\datapath.registers.838[5] [10]),
    .B(\datapath.registers.838[4] [10]),
    .S(\datapath.idinstr_20_bF$buf21 ),
    .Y(_7970_)
);

NOR2X1 _18651_ (
    .A(\datapath.registers.838[7] [10]),
    .B(_7425__bF$buf30),
    .Y(_7971_)
);

OAI21X1 _18652_ (
    .A(\datapath.registers.838[6] [10]),
    .B(\datapath.idinstr_20_bF$buf20 ),
    .C(\datapath.idinstr_21_bF$buf27 ),
    .Y(_7972_)
);

OAI22X1 _18653_ (
    .A(_7972_),
    .B(_7971_),
    .C(\datapath.idinstr_21_bF$buf26 ),
    .D(_7970_),
    .Y(_7973_)
);

OAI21X1 _18654_ (
    .A(_7420__bF$buf5),
    .B(_7973_),
    .C(_7423__bF$buf0),
    .Y(_7974_)
);

OAI22X1 _18655_ (
    .A(_7423__bF$buf7),
    .B(_7963_),
    .C(_7969_),
    .D(_7974_),
    .Y(_7975_)
);

NAND2X1 _18656_ (
    .A(_7451__bF$buf4),
    .B(_7975_),
    .Y(_7976_)
);

AOI22X1 _18657_ (
    .A(_7418__bF$buf4),
    .B(_7422__bF$buf4),
    .C(_7952_),
    .D(_7976_),
    .Y(\datapath.registers.regb_data [10])
);

NAND2X1 _18658_ (
    .A(\datapath.registers.838[27] [11]),
    .B(\datapath.idinstr_20_bF$buf19 ),
    .Y(_7977_)
);

NAND2X1 _18659_ (
    .A(\datapath.registers.838[26] [11]),
    .B(_7425__bF$buf29),
    .Y(_7978_)
);

NAND3X1 _18660_ (
    .A(\datapath.idinstr_21_bF$buf25 ),
    .B(_7977_),
    .C(_7978_),
    .Y(_7979_)
);

NAND2X1 _18661_ (
    .A(\datapath.registers.838[25] [11]),
    .B(\datapath.idinstr_20_bF$buf18 ),
    .Y(_7980_)
);

AOI21X1 _18662_ (
    .A(_7425__bF$buf28),
    .B(\datapath.registers.838[24] [11]),
    .C(\datapath.idinstr_21_bF$buf24 ),
    .Y(_7981_)
);

NAND2X1 _18663_ (
    .A(_7980_),
    .B(_7981_),
    .Y(_7982_)
);

NAND3X1 _18664_ (
    .A(_7420__bF$buf4),
    .B(_7979_),
    .C(_7982_),
    .Y(_7983_)
);

NAND2X1 _18665_ (
    .A(\datapath.registers.838[31] [11]),
    .B(\datapath.idinstr_20_bF$buf17 ),
    .Y(_7984_)
);

AOI21X1 _18666_ (
    .A(_7425__bF$buf27),
    .B(\datapath.registers.838[30] [11]),
    .C(_7419__bF$buf7),
    .Y(_7985_)
);

NAND2X1 _18667_ (
    .A(_7984_),
    .B(_7985_),
    .Y(_7986_)
);

AOI21X1 _18668_ (
    .A(\datapath.registers.838[29] [11]),
    .B(\datapath.idinstr_20_bF$buf16 ),
    .C(\datapath.idinstr_21_bF$buf23 ),
    .Y(_7987_)
);

OAI21X1 _18669_ (
    .A(_6344_),
    .B(\datapath.idinstr_20_bF$buf15 ),
    .C(_7987_),
    .Y(_7988_)
);

NAND3X1 _18670_ (
    .A(\datapath.idinstr_22_bF$buf19 ),
    .B(_7988_),
    .C(_7986_),
    .Y(_7989_)
);

AOI21X1 _18671_ (
    .A(_7983_),
    .B(_7989_),
    .C(_7423__bF$buf6),
    .Y(_7990_)
);

MUX2X1 _18672_ (
    .A(\datapath.registers.838[18] [11]),
    .B(\datapath.registers.838[16] [11]),
    .S(\datapath.idinstr_21_bF$buf22 ),
    .Y(_7991_)
);

NAND2X1 _18673_ (
    .A(_7425__bF$buf26),
    .B(_7991_),
    .Y(_7992_)
);

MUX2X1 _18674_ (
    .A(\datapath.registers.838[19] [11]),
    .B(\datapath.registers.838[17] [11]),
    .S(\datapath.idinstr_21_bF$buf21 ),
    .Y(_7993_)
);

NAND2X1 _18675_ (
    .A(\datapath.idinstr_20_bF$buf14 ),
    .B(_7993_),
    .Y(_7994_)
);

NAND3X1 _18676_ (
    .A(_7420__bF$buf3),
    .B(_7992_),
    .C(_7994_),
    .Y(_7995_)
);

MUX2X1 _18677_ (
    .A(\datapath.registers.838[22] [11]),
    .B(\datapath.registers.838[20] [11]),
    .S(\datapath.idinstr_21_bF$buf20 ),
    .Y(_7996_)
);

NAND2X1 _18678_ (
    .A(_7425__bF$buf25),
    .B(_7996_),
    .Y(_7997_)
);

MUX2X1 _18679_ (
    .A(\datapath.registers.838[23] [11]),
    .B(\datapath.registers.838[21] [11]),
    .S(\datapath.idinstr_21_bF$buf19 ),
    .Y(_7998_)
);

NAND2X1 _18680_ (
    .A(\datapath.idinstr_20_bF$buf13 ),
    .B(_7998_),
    .Y(_7999_)
);

NAND3X1 _18681_ (
    .A(\datapath.idinstr_22_bF$buf18 ),
    .B(_7997_),
    .C(_7999_),
    .Y(_8000_)
);

AOI21X1 _18682_ (
    .A(_7995_),
    .B(_8000_),
    .C(\datapath.idinstr_23_bF$buf1 ),
    .Y(_8001_)
);

OAI21X1 _18683_ (
    .A(_8001_),
    .B(_7990_),
    .C(\datapath.idinstr_24_bF$buf0 ),
    .Y(_8002_)
);

MUX2X1 _18684_ (
    .A(\datapath.registers.838[9] [11]),
    .B(\datapath.registers.838[8] [11]),
    .S(\datapath.idinstr_20_bF$buf12 ),
    .Y(_8003_)
);

NOR2X1 _18685_ (
    .A(\datapath.registers.838[11] [11]),
    .B(_7425__bF$buf24),
    .Y(_8004_)
);

OAI21X1 _18686_ (
    .A(\datapath.registers.838[10] [11]),
    .B(\datapath.idinstr_20_bF$buf11 ),
    .C(\datapath.idinstr_21_bF$buf18 ),
    .Y(_8005_)
);

OAI22X1 _18687_ (
    .A(_8005_),
    .B(_8004_),
    .C(\datapath.idinstr_21_bF$buf17 ),
    .D(_8003_),
    .Y(_8006_)
);

AOI21X1 _18688_ (
    .A(_7425__bF$buf23),
    .B(\datapath.registers.838[14] [11]),
    .C(_7419__bF$buf6),
    .Y(_8007_)
);

OAI21X1 _18689_ (
    .A(_6365_),
    .B(_7425__bF$buf22),
    .C(_8007_),
    .Y(_8008_)
);

NAND2X1 _18690_ (
    .A(\datapath.registers.838[12] [11]),
    .B(_7425__bF$buf21),
    .Y(_8009_)
);

AOI21X1 _18691_ (
    .A(\datapath.registers.838[13] [11]),
    .B(\datapath.idinstr_20_bF$buf10 ),
    .C(\datapath.idinstr_21_bF$buf16 ),
    .Y(_8010_)
);

AOI21X1 _18692_ (
    .A(_8009_),
    .B(_8010_),
    .C(_7420__bF$buf2),
    .Y(_8011_)
);

AOI22X1 _18693_ (
    .A(_8008_),
    .B(_8011_),
    .C(_7420__bF$buf1),
    .D(_8006_),
    .Y(_8012_)
);

NOR2X1 _18694_ (
    .A(\datapath.registers.838[0] [11]),
    .B(\datapath.idinstr_20_bF$buf9 ),
    .Y(_8013_)
);

OAI21X1 _18695_ (
    .A(\datapath.registers.838[1] [11]),
    .B(_7425__bF$buf20),
    .C(_7419__bF$buf5),
    .Y(_8014_)
);

NOR2X1 _18696_ (
    .A(\datapath.registers.838[3] [11]),
    .B(_7425__bF$buf19),
    .Y(_8015_)
);

OAI21X1 _18697_ (
    .A(\datapath.registers.838[2] [11]),
    .B(\datapath.idinstr_20_bF$buf8 ),
    .C(\datapath.idinstr_21_bF$buf15 ),
    .Y(_8016_)
);

OAI22X1 _18698_ (
    .A(_8015_),
    .B(_8016_),
    .C(_8013_),
    .D(_8014_),
    .Y(_8017_)
);

NOR2X1 _18699_ (
    .A(\datapath.idinstr_22_bF$buf17 ),
    .B(_8017_),
    .Y(_8018_)
);

MUX2X1 _18700_ (
    .A(\datapath.registers.838[5] [11]),
    .B(\datapath.registers.838[4] [11]),
    .S(\datapath.idinstr_20_bF$buf7 ),
    .Y(_8019_)
);

NOR2X1 _18701_ (
    .A(\datapath.registers.838[7] [11]),
    .B(_7425__bF$buf18),
    .Y(_8020_)
);

OAI21X1 _18702_ (
    .A(\datapath.registers.838[6] [11]),
    .B(\datapath.idinstr_20_bF$buf6 ),
    .C(\datapath.idinstr_21_bF$buf14 ),
    .Y(_8021_)
);

OAI22X1 _18703_ (
    .A(_8021_),
    .B(_8020_),
    .C(\datapath.idinstr_21_bF$buf13 ),
    .D(_8019_),
    .Y(_8022_)
);

OAI21X1 _18704_ (
    .A(_7420__bF$buf0),
    .B(_8022_),
    .C(_7423__bF$buf5),
    .Y(_8023_)
);

OAI22X1 _18705_ (
    .A(_7423__bF$buf4),
    .B(_8012_),
    .C(_8018_),
    .D(_8023_),
    .Y(_8024_)
);

NAND2X1 _18706_ (
    .A(_7451__bF$buf3),
    .B(_8024_),
    .Y(_8025_)
);

AOI22X1 _18707_ (
    .A(_7418__bF$buf3),
    .B(_7422__bF$buf3),
    .C(_8002_),
    .D(_8025_),
    .Y(\datapath.registers.regb_data [11])
);

NAND2X1 _18708_ (
    .A(\datapath.registers.838[27] [12]),
    .B(\datapath.idinstr_20_bF$buf5 ),
    .Y(_8026_)
);

NAND2X1 _18709_ (
    .A(\datapath.registers.838[26] [12]),
    .B(_7425__bF$buf17),
    .Y(_8027_)
);

NAND3X1 _18710_ (
    .A(\datapath.idinstr_21_bF$buf12 ),
    .B(_8026_),
    .C(_8027_),
    .Y(_8028_)
);

NAND2X1 _18711_ (
    .A(\datapath.registers.838[25] [12]),
    .B(\datapath.idinstr_20_bF$buf4 ),
    .Y(_8029_)
);

AOI21X1 _18712_ (
    .A(_7425__bF$buf16),
    .B(\datapath.registers.838[24] [12]),
    .C(\datapath.idinstr_21_bF$buf11 ),
    .Y(_8030_)
);

NAND2X1 _18713_ (
    .A(_8029_),
    .B(_8030_),
    .Y(_8031_)
);

NAND3X1 _18714_ (
    .A(_7420__bF$buf10),
    .B(_8028_),
    .C(_8031_),
    .Y(_8032_)
);

NAND2X1 _18715_ (
    .A(\datapath.registers.838[31] [12]),
    .B(\datapath.idinstr_20_bF$buf3 ),
    .Y(_8033_)
);

AOI21X1 _18716_ (
    .A(_7425__bF$buf15),
    .B(\datapath.registers.838[30] [12]),
    .C(_7419__bF$buf4),
    .Y(_8034_)
);

NAND2X1 _18717_ (
    .A(_8033_),
    .B(_8034_),
    .Y(_8035_)
);

AOI21X1 _18718_ (
    .A(\datapath.registers.838[29] [12]),
    .B(\datapath.idinstr_20_bF$buf2 ),
    .C(\datapath.idinstr_21_bF$buf10 ),
    .Y(_8036_)
);

OAI21X1 _18719_ (
    .A(_6395_),
    .B(\datapath.idinstr_20_bF$buf1 ),
    .C(_8036_),
    .Y(_8037_)
);

NAND3X1 _18720_ (
    .A(\datapath.idinstr_22_bF$buf16 ),
    .B(_8037_),
    .C(_8035_),
    .Y(_8038_)
);

AOI21X1 _18721_ (
    .A(_8032_),
    .B(_8038_),
    .C(_7423__bF$buf3),
    .Y(_8039_)
);

MUX2X1 _18722_ (
    .A(\datapath.registers.838[18] [12]),
    .B(\datapath.registers.838[16] [12]),
    .S(\datapath.idinstr_21_bF$buf9 ),
    .Y(_8040_)
);

NAND2X1 _18723_ (
    .A(_7425__bF$buf14),
    .B(_8040_),
    .Y(_8041_)
);

MUX2X1 _18724_ (
    .A(\datapath.registers.838[19] [12]),
    .B(\datapath.registers.838[17] [12]),
    .S(\datapath.idinstr_21_bF$buf8 ),
    .Y(_8042_)
);

NAND2X1 _18725_ (
    .A(\datapath.idinstr_20_bF$buf0 ),
    .B(_8042_),
    .Y(_8043_)
);

NAND3X1 _18726_ (
    .A(_7420__bF$buf9),
    .B(_8041_),
    .C(_8043_),
    .Y(_8044_)
);

MUX2X1 _18727_ (
    .A(\datapath.registers.838[22] [12]),
    .B(\datapath.registers.838[20] [12]),
    .S(\datapath.idinstr_21_bF$buf7 ),
    .Y(_8045_)
);

NAND2X1 _18728_ (
    .A(_7425__bF$buf13),
    .B(_8045_),
    .Y(_8046_)
);

MUX2X1 _18729_ (
    .A(\datapath.registers.838[23] [12]),
    .B(\datapath.registers.838[21] [12]),
    .S(\datapath.idinstr_21_bF$buf6 ),
    .Y(_8047_)
);

NAND2X1 _18730_ (
    .A(\datapath.idinstr_20_bF$buf55 ),
    .B(_8047_),
    .Y(_8048_)
);

NAND3X1 _18731_ (
    .A(\datapath.idinstr_22_bF$buf15 ),
    .B(_8046_),
    .C(_8048_),
    .Y(_8049_)
);

AOI21X1 _18732_ (
    .A(_8044_),
    .B(_8049_),
    .C(\datapath.idinstr_23_bF$buf0 ),
    .Y(_8050_)
);

OAI21X1 _18733_ (
    .A(_8050_),
    .B(_8039_),
    .C(\datapath.idinstr_24_bF$buf5 ),
    .Y(_8051_)
);

AOI21X1 _18734_ (
    .A(\datapath.registers.838[13] [12]),
    .B(\datapath.idinstr_22_bF$buf14 ),
    .C(_7425__bF$buf12),
    .Y(_8052_)
);

OAI21X1 _18735_ (
    .A(_5281_),
    .B(\datapath.idinstr_22_bF$buf13 ),
    .C(_8052_),
    .Y(_8053_)
);

INVX1 _18736_ (
    .A(\datapath.registers.838[8] [12]),
    .Y(_8054_)
);

AOI21X1 _18737_ (
    .A(\datapath.registers.838[12] [12]),
    .B(\datapath.idinstr_22_bF$buf12 ),
    .C(\datapath.idinstr_20_bF$buf54 ),
    .Y(_8055_)
);

OAI21X1 _18738_ (
    .A(_8054_),
    .B(\datapath.idinstr_22_bF$buf11 ),
    .C(_8055_),
    .Y(_8056_)
);

NAND3X1 _18739_ (
    .A(_7419__bF$buf3),
    .B(_8056_),
    .C(_8053_),
    .Y(_8057_)
);

INVX1 _18740_ (
    .A(\datapath.registers.838[11] [12]),
    .Y(_8058_)
);

AOI21X1 _18741_ (
    .A(\datapath.registers.838[15] [12]),
    .B(\datapath.idinstr_22_bF$buf10 ),
    .C(_7425__bF$buf11),
    .Y(_8059_)
);

OAI21X1 _18742_ (
    .A(_8058_),
    .B(\datapath.idinstr_22_bF$buf9 ),
    .C(_8059_),
    .Y(_8060_)
);

AOI21X1 _18743_ (
    .A(\datapath.registers.838[14] [12]),
    .B(\datapath.idinstr_22_bF$buf8 ),
    .C(\datapath.idinstr_20_bF$buf53 ),
    .Y(_8061_)
);

OAI21X1 _18744_ (
    .A(_5237_),
    .B(\datapath.idinstr_22_bF$buf7 ),
    .C(_8061_),
    .Y(_8062_)
);

NAND3X1 _18745_ (
    .A(\datapath.idinstr_21_bF$buf5 ),
    .B(_8062_),
    .C(_8060_),
    .Y(_8063_)
);

AOI21X1 _18746_ (
    .A(_8057_),
    .B(_8063_),
    .C(_7423__bF$buf2),
    .Y(_8064_)
);

MUX2X1 _18747_ (
    .A(\datapath.registers.838[1] [12]),
    .B(\datapath.registers.838[0] [12]),
    .S(\datapath.idinstr_20_bF$buf52 ),
    .Y(_8065_)
);

NOR2X1 _18748_ (
    .A(\datapath.registers.838[3] [12]),
    .B(_7425__bF$buf10),
    .Y(_8066_)
);

OAI21X1 _18749_ (
    .A(\datapath.registers.838[2] [12]),
    .B(\datapath.idinstr_20_bF$buf51 ),
    .C(\datapath.idinstr_21_bF$buf4 ),
    .Y(_8067_)
);

OAI22X1 _18750_ (
    .A(_8067_),
    .B(_8066_),
    .C(\datapath.idinstr_21_bF$buf3 ),
    .D(_8065_),
    .Y(_8068_)
);

NAND2X1 _18751_ (
    .A(_7420__bF$buf8),
    .B(_8068_),
    .Y(_8069_)
);

MUX2X1 _18752_ (
    .A(\datapath.registers.838[5] [12]),
    .B(\datapath.registers.838[4] [12]),
    .S(\datapath.idinstr_20_bF$buf50 ),
    .Y(_8070_)
);

NOR2X1 _18753_ (
    .A(\datapath.registers.838[7] [12]),
    .B(_7425__bF$buf9),
    .Y(_8071_)
);

OAI21X1 _18754_ (
    .A(\datapath.registers.838[6] [12]),
    .B(\datapath.idinstr_20_bF$buf49 ),
    .C(\datapath.idinstr_21_bF$buf2 ),
    .Y(_8072_)
);

OAI22X1 _18755_ (
    .A(_8072_),
    .B(_8071_),
    .C(\datapath.idinstr_21_bF$buf1 ),
    .D(_8070_),
    .Y(_8073_)
);

NAND2X1 _18756_ (
    .A(\datapath.idinstr_22_bF$buf6 ),
    .B(_8073_),
    .Y(_8074_)
);

AOI21X1 _18757_ (
    .A(_8069_),
    .B(_8074_),
    .C(\datapath.idinstr_23_bF$buf6 ),
    .Y(_8075_)
);

OAI21X1 _18758_ (
    .A(_8064_),
    .B(_8075_),
    .C(_7451__bF$buf2),
    .Y(_8076_)
);

AOI22X1 _18759_ (
    .A(_7418__bF$buf2),
    .B(_7422__bF$buf2),
    .C(_8051_),
    .D(_8076_),
    .Y(\datapath.registers.regb_data [12])
);

NAND2X1 _18760_ (
    .A(\datapath.registers.838[27] [13]),
    .B(\datapath.idinstr_20_bF$buf48 ),
    .Y(_8077_)
);

NAND2X1 _18761_ (
    .A(\datapath.registers.838[26] [13]),
    .B(_7425__bF$buf8),
    .Y(_8078_)
);

NAND3X1 _18762_ (
    .A(\datapath.idinstr_21_bF$buf0 ),
    .B(_8077_),
    .C(_8078_),
    .Y(_8079_)
);

NAND2X1 _18763_ (
    .A(\datapath.registers.838[25] [13]),
    .B(\datapath.idinstr_20_bF$buf47 ),
    .Y(_8080_)
);

AOI21X1 _18764_ (
    .A(_7425__bF$buf7),
    .B(\datapath.registers.838[24] [13]),
    .C(\datapath.idinstr_21_bF$buf51 ),
    .Y(_8081_)
);

NAND2X1 _18765_ (
    .A(_8080_),
    .B(_8081_),
    .Y(_8082_)
);

NAND3X1 _18766_ (
    .A(_7420__bF$buf7),
    .B(_8079_),
    .C(_8082_),
    .Y(_8083_)
);

NAND2X1 _18767_ (
    .A(\datapath.registers.838[31] [13]),
    .B(\datapath.idinstr_20_bF$buf46 ),
    .Y(_8084_)
);

AOI21X1 _18768_ (
    .A(_7425__bF$buf6),
    .B(\datapath.registers.838[30] [13]),
    .C(_7419__bF$buf2),
    .Y(_8085_)
);

NAND2X1 _18769_ (
    .A(_8084_),
    .B(_8085_),
    .Y(_8086_)
);

AOI21X1 _18770_ (
    .A(\datapath.registers.838[29] [13]),
    .B(\datapath.idinstr_20_bF$buf45 ),
    .C(\datapath.idinstr_21_bF$buf50 ),
    .Y(_8087_)
);

OAI21X1 _18771_ (
    .A(_6452_),
    .B(\datapath.idinstr_20_bF$buf44 ),
    .C(_8087_),
    .Y(_8088_)
);

NAND3X1 _18772_ (
    .A(\datapath.idinstr_22_bF$buf5 ),
    .B(_8088_),
    .C(_8086_),
    .Y(_8089_)
);

AOI21X1 _18773_ (
    .A(_8083_),
    .B(_8089_),
    .C(_7423__bF$buf1),
    .Y(_8090_)
);

MUX2X1 _18774_ (
    .A(\datapath.registers.838[18] [13]),
    .B(\datapath.registers.838[16] [13]),
    .S(\datapath.idinstr_21_bF$buf49 ),
    .Y(_8091_)
);

NAND2X1 _18775_ (
    .A(_7425__bF$buf5),
    .B(_8091_),
    .Y(_8092_)
);

MUX2X1 _18776_ (
    .A(\datapath.registers.838[19] [13]),
    .B(\datapath.registers.838[17] [13]),
    .S(\datapath.idinstr_21_bF$buf48 ),
    .Y(_8093_)
);

NAND2X1 _18777_ (
    .A(\datapath.idinstr_20_bF$buf43 ),
    .B(_8093_),
    .Y(_8094_)
);

NAND3X1 _18778_ (
    .A(_7420__bF$buf6),
    .B(_8092_),
    .C(_8094_),
    .Y(_8095_)
);

MUX2X1 _18779_ (
    .A(\datapath.registers.838[22] [13]),
    .B(\datapath.registers.838[20] [13]),
    .S(\datapath.idinstr_21_bF$buf47 ),
    .Y(_8096_)
);

NAND2X1 _18780_ (
    .A(_7425__bF$buf4),
    .B(_8096_),
    .Y(_8097_)
);

MUX2X1 _18781_ (
    .A(\datapath.registers.838[23] [13]),
    .B(\datapath.registers.838[21] [13]),
    .S(\datapath.idinstr_21_bF$buf46 ),
    .Y(_8098_)
);

NAND2X1 _18782_ (
    .A(\datapath.idinstr_20_bF$buf42 ),
    .B(_8098_),
    .Y(_8099_)
);

NAND3X1 _18783_ (
    .A(\datapath.idinstr_22_bF$buf4 ),
    .B(_8097_),
    .C(_8099_),
    .Y(_8100_)
);

AOI21X1 _18784_ (
    .A(_8095_),
    .B(_8100_),
    .C(\datapath.idinstr_23_bF$buf5 ),
    .Y(_8101_)
);

OAI21X1 _18785_ (
    .A(_8101_),
    .B(_8090_),
    .C(\datapath.idinstr_24_bF$buf4 ),
    .Y(_8102_)
);

MUX2X1 _18786_ (
    .A(\datapath.registers.838[9] [13]),
    .B(\datapath.registers.838[8] [13]),
    .S(\datapath.idinstr_20_bF$buf41 ),
    .Y(_8103_)
);

NOR2X1 _18787_ (
    .A(\datapath.registers.838[11] [13]),
    .B(_7425__bF$buf3),
    .Y(_8104_)
);

OAI21X1 _18788_ (
    .A(\datapath.registers.838[10] [13]),
    .B(\datapath.idinstr_20_bF$buf40 ),
    .C(\datapath.idinstr_21_bF$buf45 ),
    .Y(_8105_)
);

OAI22X1 _18789_ (
    .A(_8105_),
    .B(_8104_),
    .C(\datapath.idinstr_21_bF$buf44 ),
    .D(_8103_),
    .Y(_8106_)
);

AOI21X1 _18790_ (
    .A(_7425__bF$buf2),
    .B(\datapath.registers.838[14] [13]),
    .C(_7419__bF$buf1),
    .Y(_8107_)
);

OAI21X1 _18791_ (
    .A(_6473_),
    .B(_7425__bF$buf1),
    .C(_8107_),
    .Y(_8108_)
);

NAND2X1 _18792_ (
    .A(\datapath.registers.838[12] [13]),
    .B(_7425__bF$buf0),
    .Y(_8109_)
);

AOI21X1 _18793_ (
    .A(\datapath.registers.838[13] [13]),
    .B(\datapath.idinstr_20_bF$buf39 ),
    .C(\datapath.idinstr_21_bF$buf43 ),
    .Y(_8110_)
);

AOI21X1 _18794_ (
    .A(_8109_),
    .B(_8110_),
    .C(_7420__bF$buf5),
    .Y(_8111_)
);

AOI22X1 _18795_ (
    .A(_8108_),
    .B(_8111_),
    .C(_7420__bF$buf4),
    .D(_8106_),
    .Y(_8112_)
);

NOR2X1 _18796_ (
    .A(\datapath.registers.838[0] [13]),
    .B(\datapath.idinstr_20_bF$buf38 ),
    .Y(_8113_)
);

OAI21X1 _18797_ (
    .A(\datapath.registers.838[1] [13]),
    .B(_7425__bF$buf47),
    .C(_7419__bF$buf0),
    .Y(_8114_)
);

NOR2X1 _18798_ (
    .A(\datapath.registers.838[3] [13]),
    .B(_7425__bF$buf46),
    .Y(_8115_)
);

OAI21X1 _18799_ (
    .A(\datapath.registers.838[2] [13]),
    .B(\datapath.idinstr_20_bF$buf37 ),
    .C(\datapath.idinstr_21_bF$buf42 ),
    .Y(_8116_)
);

OAI22X1 _18800_ (
    .A(_8115_),
    .B(_8116_),
    .C(_8113_),
    .D(_8114_),
    .Y(_8117_)
);

NOR2X1 _18801_ (
    .A(\datapath.idinstr_22_bF$buf3 ),
    .B(_8117_),
    .Y(_8118_)
);

MUX2X1 _18802_ (
    .A(\datapath.registers.838[5] [13]),
    .B(\datapath.registers.838[4] [13]),
    .S(\datapath.idinstr_20_bF$buf36 ),
    .Y(_8119_)
);

NOR2X1 _18803_ (
    .A(\datapath.registers.838[7] [13]),
    .B(_7425__bF$buf45),
    .Y(_8120_)
);

OAI21X1 _18804_ (
    .A(\datapath.registers.838[6] [13]),
    .B(\datapath.idinstr_20_bF$buf35 ),
    .C(\datapath.idinstr_21_bF$buf41 ),
    .Y(_8121_)
);

OAI22X1 _18805_ (
    .A(_8121_),
    .B(_8120_),
    .C(\datapath.idinstr_21_bF$buf40 ),
    .D(_8119_),
    .Y(_8122_)
);

OAI21X1 _18806_ (
    .A(_7420__bF$buf3),
    .B(_8122_),
    .C(_7423__bF$buf0),
    .Y(_8123_)
);

OAI22X1 _18807_ (
    .A(_7423__bF$buf7),
    .B(_8112_),
    .C(_8118_),
    .D(_8123_),
    .Y(_8124_)
);

NAND2X1 _18808_ (
    .A(_7451__bF$buf1),
    .B(_8124_),
    .Y(_8125_)
);

AOI22X1 _18809_ (
    .A(_7418__bF$buf1),
    .B(_7422__bF$buf1),
    .C(_8102_),
    .D(_8125_),
    .Y(\datapath.registers.regb_data [13])
);

MUX2X1 _18810_ (
    .A(\datapath.registers.838[9] [14]),
    .B(\datapath.registers.838[8] [14]),
    .S(\datapath.idinstr_20_bF$buf34 ),
    .Y(_8126_)
);

NOR2X1 _18811_ (
    .A(\datapath.registers.838[11] [14]),
    .B(_7425__bF$buf44),
    .Y(_8127_)
);

OAI21X1 _18812_ (
    .A(\datapath.registers.838[10] [14]),
    .B(\datapath.idinstr_20_bF$buf33 ),
    .C(\datapath.idinstr_21_bF$buf39 ),
    .Y(_8128_)
);

OAI22X1 _18813_ (
    .A(_8128_),
    .B(_8127_),
    .C(\datapath.idinstr_21_bF$buf38 ),
    .D(_8126_),
    .Y(_8129_)
);

AOI21X1 _18814_ (
    .A(_7425__bF$buf43),
    .B(\datapath.registers.838[14] [14]),
    .C(_7419__bF$buf9),
    .Y(_8130_)
);

OAI21X1 _18815_ (
    .A(_6524_),
    .B(_7425__bF$buf42),
    .C(_8130_),
    .Y(_8131_)
);

NAND2X1 _18816_ (
    .A(\datapath.registers.838[12] [14]),
    .B(_7425__bF$buf41),
    .Y(_8132_)
);

AOI21X1 _18817_ (
    .A(\datapath.registers.838[13] [14]),
    .B(\datapath.idinstr_20_bF$buf32 ),
    .C(\datapath.idinstr_21_bF$buf37 ),
    .Y(_8133_)
);

AOI21X1 _18818_ (
    .A(_8132_),
    .B(_8133_),
    .C(_7420__bF$buf2),
    .Y(_8134_)
);

AOI22X1 _18819_ (
    .A(_8131_),
    .B(_8134_),
    .C(_7420__bF$buf1),
    .D(_8129_),
    .Y(_8135_)
);

NOR2X1 _18820_ (
    .A(\datapath.registers.838[0] [14]),
    .B(\datapath.idinstr_20_bF$buf31 ),
    .Y(_8136_)
);

OAI21X1 _18821_ (
    .A(\datapath.registers.838[1] [14]),
    .B(_7425__bF$buf40),
    .C(_7419__bF$buf8),
    .Y(_8137_)
);

NOR2X1 _18822_ (
    .A(\datapath.registers.838[3] [14]),
    .B(_7425__bF$buf39),
    .Y(_8138_)
);

OAI21X1 _18823_ (
    .A(\datapath.registers.838[2] [14]),
    .B(\datapath.idinstr_20_bF$buf30 ),
    .C(\datapath.idinstr_21_bF$buf36 ),
    .Y(_8139_)
);

OAI22X1 _18824_ (
    .A(_8138_),
    .B(_8139_),
    .C(_8136_),
    .D(_8137_),
    .Y(_8140_)
);

NOR2X1 _18825_ (
    .A(\datapath.idinstr_22_bF$buf2 ),
    .B(_8140_),
    .Y(_8141_)
);

MUX2X1 _18826_ (
    .A(\datapath.registers.838[5] [14]),
    .B(\datapath.registers.838[4] [14]),
    .S(\datapath.idinstr_20_bF$buf29 ),
    .Y(_8142_)
);

NOR2X1 _18827_ (
    .A(\datapath.registers.838[7] [14]),
    .B(_7425__bF$buf38),
    .Y(_8143_)
);

OAI21X1 _18828_ (
    .A(\datapath.registers.838[6] [14]),
    .B(\datapath.idinstr_20_bF$buf28 ),
    .C(\datapath.idinstr_21_bF$buf35 ),
    .Y(_8144_)
);

OAI22X1 _18829_ (
    .A(_8144_),
    .B(_8143_),
    .C(\datapath.idinstr_21_bF$buf34 ),
    .D(_8142_),
    .Y(_8145_)
);

OAI21X1 _18830_ (
    .A(_7420__bF$buf0),
    .B(_8145_),
    .C(_7423__bF$buf6),
    .Y(_8146_)
);

OAI22X1 _18831_ (
    .A(_7423__bF$buf5),
    .B(_8135_),
    .C(_8141_),
    .D(_8146_),
    .Y(_8147_)
);

NAND2X1 _18832_ (
    .A(_7451__bF$buf0),
    .B(_8147_),
    .Y(_8148_)
);

INVX1 _18833_ (
    .A(\datapath.registers.838[27] [14]),
    .Y(_8149_)
);

AOI21X1 _18834_ (
    .A(\datapath.registers.838[31] [14]),
    .B(\datapath.idinstr_22_bF$buf1 ),
    .C(_7425__bF$buf37),
    .Y(_8150_)
);

OAI21X1 _18835_ (
    .A(_8149_),
    .B(\datapath.idinstr_22_bF$buf0 ),
    .C(_8150_),
    .Y(_8151_)
);

INVX1 _18836_ (
    .A(\datapath.registers.838[26] [14]),
    .Y(_8152_)
);

AOI21X1 _18837_ (
    .A(\datapath.registers.838[30] [14]),
    .B(\datapath.idinstr_22_bF$buf41 ),
    .C(\datapath.idinstr_20_bF$buf27 ),
    .Y(_8153_)
);

OAI21X1 _18838_ (
    .A(_8152_),
    .B(\datapath.idinstr_22_bF$buf40 ),
    .C(_8153_),
    .Y(_8154_)
);

NAND3X1 _18839_ (
    .A(\datapath.idinstr_21_bF$buf33 ),
    .B(_8154_),
    .C(_8151_),
    .Y(_8155_)
);

INVX1 _18840_ (
    .A(\datapath.registers.838[25] [14]),
    .Y(_8156_)
);

AOI21X1 _18841_ (
    .A(\datapath.registers.838[29] [14]),
    .B(\datapath.idinstr_22_bF$buf39 ),
    .C(_7425__bF$buf36),
    .Y(_8157_)
);

OAI21X1 _18842_ (
    .A(_8156_),
    .B(\datapath.idinstr_22_bF$buf38 ),
    .C(_8157_),
    .Y(_8158_)
);

INVX1 _18843_ (
    .A(\datapath.registers.838[24] [14]),
    .Y(_8159_)
);

AOI21X1 _18844_ (
    .A(\datapath.registers.838[28] [14]),
    .B(\datapath.idinstr_22_bF$buf37 ),
    .C(\datapath.idinstr_20_bF$buf26 ),
    .Y(_8160_)
);

OAI21X1 _18845_ (
    .A(_8159_),
    .B(\datapath.idinstr_22_bF$buf36 ),
    .C(_8160_),
    .Y(_8161_)
);

NAND3X1 _18846_ (
    .A(_7419__bF$buf7),
    .B(_8161_),
    .C(_8158_),
    .Y(_8162_)
);

AOI21X1 _18847_ (
    .A(_8155_),
    .B(_8162_),
    .C(_7423__bF$buf4),
    .Y(_8163_)
);

MUX2X1 _18848_ (
    .A(\datapath.registers.838[18] [14]),
    .B(\datapath.registers.838[16] [14]),
    .S(\datapath.idinstr_21_bF$buf32 ),
    .Y(_8164_)
);

NAND2X1 _18849_ (
    .A(_7425__bF$buf35),
    .B(_8164_),
    .Y(_8165_)
);

MUX2X1 _18850_ (
    .A(\datapath.registers.838[19] [14]),
    .B(\datapath.registers.838[17] [14]),
    .S(\datapath.idinstr_21_bF$buf31 ),
    .Y(_8166_)
);

NAND2X1 _18851_ (
    .A(\datapath.idinstr_20_bF$buf25 ),
    .B(_8166_),
    .Y(_8167_)
);

NAND3X1 _18852_ (
    .A(_7420__bF$buf10),
    .B(_8165_),
    .C(_8167_),
    .Y(_8168_)
);

MUX2X1 _18853_ (
    .A(\datapath.registers.838[22] [14]),
    .B(\datapath.registers.838[20] [14]),
    .S(\datapath.idinstr_21_bF$buf30 ),
    .Y(_8169_)
);

NAND2X1 _18854_ (
    .A(_7425__bF$buf34),
    .B(_8169_),
    .Y(_8170_)
);

MUX2X1 _18855_ (
    .A(\datapath.registers.838[23] [14]),
    .B(\datapath.registers.838[21] [14]),
    .S(\datapath.idinstr_21_bF$buf29 ),
    .Y(_8171_)
);

NAND2X1 _18856_ (
    .A(\datapath.idinstr_20_bF$buf24 ),
    .B(_8171_),
    .Y(_8172_)
);

NAND3X1 _18857_ (
    .A(\datapath.idinstr_22_bF$buf35 ),
    .B(_8170_),
    .C(_8172_),
    .Y(_8173_)
);

AOI21X1 _18858_ (
    .A(_8168_),
    .B(_8173_),
    .C(\datapath.idinstr_23_bF$buf4 ),
    .Y(_8174_)
);

OAI21X1 _18859_ (
    .A(_8163_),
    .B(_8174_),
    .C(\datapath.idinstr_24_bF$buf3 ),
    .Y(_8175_)
);

AOI22X1 _18860_ (
    .A(_7418__bF$buf0),
    .B(_7422__bF$buf0),
    .C(_8175_),
    .D(_8148_),
    .Y(\datapath.registers.regb_data [14])
);

MUX2X1 _18861_ (
    .A(\datapath.registers.838[9] [15]),
    .B(\datapath.registers.838[8] [15]),
    .S(\datapath.idinstr_20_bF$buf23 ),
    .Y(_8176_)
);

NOR2X1 _18862_ (
    .A(\datapath.registers.838[11] [15]),
    .B(_7425__bF$buf33),
    .Y(_8177_)
);

OAI21X1 _18863_ (
    .A(\datapath.registers.838[10] [15]),
    .B(\datapath.idinstr_20_bF$buf22 ),
    .C(\datapath.idinstr_21_bF$buf28 ),
    .Y(_8178_)
);

OAI22X1 _18864_ (
    .A(_8178_),
    .B(_8177_),
    .C(\datapath.idinstr_21_bF$buf27 ),
    .D(_8176_),
    .Y(_8179_)
);

AOI21X1 _18865_ (
    .A(_7425__bF$buf32),
    .B(\datapath.registers.838[14] [15]),
    .C(_7419__bF$buf6),
    .Y(_8180_)
);

OAI21X1 _18866_ (
    .A(_6548_),
    .B(_7425__bF$buf31),
    .C(_8180_),
    .Y(_8181_)
);

NAND2X1 _18867_ (
    .A(\datapath.registers.838[12] [15]),
    .B(_7425__bF$buf30),
    .Y(_8182_)
);

AOI21X1 _18868_ (
    .A(\datapath.registers.838[13] [15]),
    .B(\datapath.idinstr_20_bF$buf21 ),
    .C(\datapath.idinstr_21_bF$buf26 ),
    .Y(_8183_)
);

AOI21X1 _18869_ (
    .A(_8182_),
    .B(_8183_),
    .C(_7420__bF$buf9),
    .Y(_8184_)
);

AOI22X1 _18870_ (
    .A(_8181_),
    .B(_8184_),
    .C(_7420__bF$buf8),
    .D(_8179_),
    .Y(_8185_)
);

NOR2X1 _18871_ (
    .A(\datapath.registers.838[0] [15]),
    .B(\datapath.idinstr_20_bF$buf20 ),
    .Y(_8186_)
);

OAI21X1 _18872_ (
    .A(\datapath.registers.838[1] [15]),
    .B(_7425__bF$buf29),
    .C(_7419__bF$buf5),
    .Y(_8187_)
);

NOR2X1 _18873_ (
    .A(\datapath.registers.838[3] [15]),
    .B(_7425__bF$buf28),
    .Y(_8188_)
);

OAI21X1 _18874_ (
    .A(\datapath.registers.838[2] [15]),
    .B(\datapath.idinstr_20_bF$buf19 ),
    .C(\datapath.idinstr_21_bF$buf25 ),
    .Y(_8189_)
);

OAI22X1 _18875_ (
    .A(_8188_),
    .B(_8189_),
    .C(_8186_),
    .D(_8187_),
    .Y(_8190_)
);

NOR2X1 _18876_ (
    .A(\datapath.idinstr_22_bF$buf34 ),
    .B(_8190_),
    .Y(_8191_)
);

MUX2X1 _18877_ (
    .A(\datapath.registers.838[5] [15]),
    .B(\datapath.registers.838[4] [15]),
    .S(\datapath.idinstr_20_bF$buf18 ),
    .Y(_8192_)
);

NOR2X1 _18878_ (
    .A(\datapath.registers.838[7] [15]),
    .B(_7425__bF$buf27),
    .Y(_8193_)
);

OAI21X1 _18879_ (
    .A(\datapath.registers.838[6] [15]),
    .B(\datapath.idinstr_20_bF$buf17 ),
    .C(\datapath.idinstr_21_bF$buf24 ),
    .Y(_8194_)
);

OAI22X1 _18880_ (
    .A(_8194_),
    .B(_8193_),
    .C(\datapath.idinstr_21_bF$buf23 ),
    .D(_8192_),
    .Y(_8195_)
);

OAI21X1 _18881_ (
    .A(_7420__bF$buf7),
    .B(_8195_),
    .C(_7423__bF$buf3),
    .Y(_8196_)
);

OAI22X1 _18882_ (
    .A(_7423__bF$buf2),
    .B(_8185_),
    .C(_8191_),
    .D(_8196_),
    .Y(_8197_)
);

NAND2X1 _18883_ (
    .A(_7451__bF$buf4),
    .B(_8197_),
    .Y(_8198_)
);

AOI21X1 _18884_ (
    .A(\datapath.registers.838[31] [15]),
    .B(\datapath.idinstr_22_bF$buf33 ),
    .C(_7425__bF$buf26),
    .Y(_8199_)
);

OAI21X1 _18885_ (
    .A(_6568_),
    .B(\datapath.idinstr_22_bF$buf32 ),
    .C(_8199_),
    .Y(_8200_)
);

AOI21X1 _18886_ (
    .A(\datapath.registers.838[30] [15]),
    .B(\datapath.idinstr_22_bF$buf31 ),
    .C(\datapath.idinstr_20_bF$buf16 ),
    .Y(_8201_)
);

OAI21X1 _18887_ (
    .A(_6571_),
    .B(\datapath.idinstr_22_bF$buf30 ),
    .C(_8201_),
    .Y(_8202_)
);

NAND3X1 _18888_ (
    .A(\datapath.idinstr_21_bF$buf22 ),
    .B(_8202_),
    .C(_8200_),
    .Y(_8203_)
);

AOI21X1 _18889_ (
    .A(\datapath.registers.838[29] [15]),
    .B(\datapath.idinstr_22_bF$buf29 ),
    .C(_7425__bF$buf25),
    .Y(_8204_)
);

OAI21X1 _18890_ (
    .A(_6575_),
    .B(\datapath.idinstr_22_bF$buf28 ),
    .C(_8204_),
    .Y(_8205_)
);

AOI21X1 _18891_ (
    .A(\datapath.registers.838[28] [15]),
    .B(\datapath.idinstr_22_bF$buf27 ),
    .C(\datapath.idinstr_20_bF$buf15 ),
    .Y(_8206_)
);

OAI21X1 _18892_ (
    .A(_6578_),
    .B(\datapath.idinstr_22_bF$buf26 ),
    .C(_8206_),
    .Y(_8207_)
);

NAND3X1 _18893_ (
    .A(_7419__bF$buf4),
    .B(_8207_),
    .C(_8205_),
    .Y(_8208_)
);

AOI21X1 _18894_ (
    .A(_8203_),
    .B(_8208_),
    .C(_7423__bF$buf1),
    .Y(_8209_)
);

MUX2X1 _18895_ (
    .A(\datapath.registers.838[18] [15]),
    .B(\datapath.registers.838[16] [15]),
    .S(\datapath.idinstr_21_bF$buf21 ),
    .Y(_8210_)
);

NAND2X1 _18896_ (
    .A(_7425__bF$buf24),
    .B(_8210_),
    .Y(_8211_)
);

MUX2X1 _18897_ (
    .A(\datapath.registers.838[19] [15]),
    .B(\datapath.registers.838[17] [15]),
    .S(\datapath.idinstr_21_bF$buf20 ),
    .Y(_8212_)
);

NAND2X1 _18898_ (
    .A(\datapath.idinstr_20_bF$buf14 ),
    .B(_8212_),
    .Y(_8213_)
);

NAND3X1 _18899_ (
    .A(_7420__bF$buf6),
    .B(_8211_),
    .C(_8213_),
    .Y(_8214_)
);

MUX2X1 _18900_ (
    .A(\datapath.registers.838[22] [15]),
    .B(\datapath.registers.838[20] [15]),
    .S(\datapath.idinstr_21_bF$buf19 ),
    .Y(_8215_)
);

NAND2X1 _18901_ (
    .A(_7425__bF$buf23),
    .B(_8215_),
    .Y(_8216_)
);

MUX2X1 _18902_ (
    .A(\datapath.registers.838[23] [15]),
    .B(\datapath.registers.838[21] [15]),
    .S(\datapath.idinstr_21_bF$buf18 ),
    .Y(_8217_)
);

NAND2X1 _18903_ (
    .A(\datapath.idinstr_20_bF$buf13 ),
    .B(_8217_),
    .Y(_8218_)
);

NAND3X1 _18904_ (
    .A(\datapath.idinstr_22_bF$buf25 ),
    .B(_8216_),
    .C(_8218_),
    .Y(_8219_)
);

AOI21X1 _18905_ (
    .A(_8214_),
    .B(_8219_),
    .C(\datapath.idinstr_23_bF$buf3 ),
    .Y(_8220_)
);

OAI21X1 _18906_ (
    .A(_8209_),
    .B(_8220_),
    .C(\datapath.idinstr_24_bF$buf2 ),
    .Y(_8221_)
);

AOI22X1 _18907_ (
    .A(_7418__bF$buf4),
    .B(_7422__bF$buf4),
    .C(_8221_),
    .D(_8198_),
    .Y(\datapath.registers.regb_data [15])
);

MUX2X1 _18908_ (
    .A(\datapath.registers.838[9] [16]),
    .B(\datapath.registers.838[8] [16]),
    .S(\datapath.idinstr_20_bF$buf12 ),
    .Y(_8222_)
);

NOR2X1 _18909_ (
    .A(\datapath.registers.838[11] [16]),
    .B(_7425__bF$buf22),
    .Y(_8223_)
);

OAI21X1 _18910_ (
    .A(\datapath.registers.838[10] [16]),
    .B(\datapath.idinstr_20_bF$buf11 ),
    .C(\datapath.idinstr_21_bF$buf17 ),
    .Y(_8224_)
);

OAI22X1 _18911_ (
    .A(_8224_),
    .B(_8223_),
    .C(\datapath.idinstr_21_bF$buf16 ),
    .D(_8222_),
    .Y(_8225_)
);

AOI21X1 _18912_ (
    .A(_7425__bF$buf21),
    .B(\datapath.registers.838[14] [16]),
    .C(_7419__bF$buf3),
    .Y(_8226_)
);

OAI21X1 _18913_ (
    .A(_6599_),
    .B(_7425__bF$buf20),
    .C(_8226_),
    .Y(_8227_)
);

NAND2X1 _18914_ (
    .A(\datapath.registers.838[12] [16]),
    .B(_7425__bF$buf19),
    .Y(_8228_)
);

AOI21X1 _18915_ (
    .A(\datapath.registers.838[13] [16]),
    .B(\datapath.idinstr_20_bF$buf10 ),
    .C(\datapath.idinstr_21_bF$buf15 ),
    .Y(_8229_)
);

AOI21X1 _18916_ (
    .A(_8228_),
    .B(_8229_),
    .C(_7420__bF$buf5),
    .Y(_8230_)
);

AOI22X1 _18917_ (
    .A(_8227_),
    .B(_8230_),
    .C(_7420__bF$buf4),
    .D(_8225_),
    .Y(_8231_)
);

NOR2X1 _18918_ (
    .A(\datapath.registers.838[0] [16]),
    .B(\datapath.idinstr_20_bF$buf9 ),
    .Y(_8232_)
);

OAI21X1 _18919_ (
    .A(\datapath.registers.838[1] [16]),
    .B(_7425__bF$buf18),
    .C(_7419__bF$buf2),
    .Y(_8233_)
);

NOR2X1 _18920_ (
    .A(\datapath.registers.838[3] [16]),
    .B(_7425__bF$buf17),
    .Y(_8234_)
);

OAI21X1 _18921_ (
    .A(\datapath.registers.838[2] [16]),
    .B(\datapath.idinstr_20_bF$buf8 ),
    .C(\datapath.idinstr_21_bF$buf14 ),
    .Y(_8235_)
);

OAI22X1 _18922_ (
    .A(_8234_),
    .B(_8235_),
    .C(_8232_),
    .D(_8233_),
    .Y(_8236_)
);

NOR2X1 _18923_ (
    .A(\datapath.idinstr_22_bF$buf24 ),
    .B(_8236_),
    .Y(_8237_)
);

MUX2X1 _18924_ (
    .A(\datapath.registers.838[5] [16]),
    .B(\datapath.registers.838[4] [16]),
    .S(\datapath.idinstr_20_bF$buf7 ),
    .Y(_8238_)
);

NOR2X1 _18925_ (
    .A(\datapath.registers.838[7] [16]),
    .B(_7425__bF$buf16),
    .Y(_8239_)
);

OAI21X1 _18926_ (
    .A(\datapath.registers.838[6] [16]),
    .B(\datapath.idinstr_20_bF$buf6 ),
    .C(\datapath.idinstr_21_bF$buf13 ),
    .Y(_8240_)
);

OAI22X1 _18927_ (
    .A(_8240_),
    .B(_8239_),
    .C(\datapath.idinstr_21_bF$buf12 ),
    .D(_8238_),
    .Y(_8241_)
);

OAI21X1 _18928_ (
    .A(_7420__bF$buf3),
    .B(_8241_),
    .C(_7423__bF$buf0),
    .Y(_8242_)
);

OAI22X1 _18929_ (
    .A(_7423__bF$buf7),
    .B(_8231_),
    .C(_8237_),
    .D(_8242_),
    .Y(_8243_)
);

NAND2X1 _18930_ (
    .A(_7451__bF$buf3),
    .B(_8243_),
    .Y(_8244_)
);

AOI21X1 _18931_ (
    .A(\datapath.registers.838[31] [16]),
    .B(\datapath.idinstr_22_bF$buf23 ),
    .C(_7425__bF$buf15),
    .Y(_8245_)
);

OAI21X1 _18932_ (
    .A(_6619_),
    .B(\datapath.idinstr_22_bF$buf22 ),
    .C(_8245_),
    .Y(_8246_)
);

AOI21X1 _18933_ (
    .A(\datapath.registers.838[30] [16]),
    .B(\datapath.idinstr_22_bF$buf21 ),
    .C(\datapath.idinstr_20_bF$buf5 ),
    .Y(_8247_)
);

OAI21X1 _18934_ (
    .A(_6622_),
    .B(\datapath.idinstr_22_bF$buf20 ),
    .C(_8247_),
    .Y(_8248_)
);

NAND3X1 _18935_ (
    .A(\datapath.idinstr_21_bF$buf11 ),
    .B(_8248_),
    .C(_8246_),
    .Y(_8249_)
);

AOI21X1 _18936_ (
    .A(\datapath.registers.838[29] [16]),
    .B(\datapath.idinstr_22_bF$buf19 ),
    .C(_7425__bF$buf14),
    .Y(_8250_)
);

OAI21X1 _18937_ (
    .A(_6626_),
    .B(\datapath.idinstr_22_bF$buf18 ),
    .C(_8250_),
    .Y(_8251_)
);

AOI21X1 _18938_ (
    .A(\datapath.registers.838[28] [16]),
    .B(\datapath.idinstr_22_bF$buf17 ),
    .C(\datapath.idinstr_20_bF$buf4 ),
    .Y(_8252_)
);

OAI21X1 _18939_ (
    .A(_6629_),
    .B(\datapath.idinstr_22_bF$buf16 ),
    .C(_8252_),
    .Y(_8253_)
);

NAND3X1 _18940_ (
    .A(_7419__bF$buf1),
    .B(_8253_),
    .C(_8251_),
    .Y(_8254_)
);

AOI21X1 _18941_ (
    .A(_8249_),
    .B(_8254_),
    .C(_7423__bF$buf6),
    .Y(_8255_)
);

MUX2X1 _18942_ (
    .A(\datapath.registers.838[18] [16]),
    .B(\datapath.registers.838[16] [16]),
    .S(\datapath.idinstr_21_bF$buf10 ),
    .Y(_8256_)
);

NAND2X1 _18943_ (
    .A(_7425__bF$buf13),
    .B(_8256_),
    .Y(_8257_)
);

MUX2X1 _18944_ (
    .A(\datapath.registers.838[19] [16]),
    .B(\datapath.registers.838[17] [16]),
    .S(\datapath.idinstr_21_bF$buf9 ),
    .Y(_8258_)
);

NAND2X1 _18945_ (
    .A(\datapath.idinstr_20_bF$buf3 ),
    .B(_8258_),
    .Y(_8259_)
);

NAND3X1 _18946_ (
    .A(_7420__bF$buf2),
    .B(_8257_),
    .C(_8259_),
    .Y(_8260_)
);

MUX2X1 _18947_ (
    .A(\datapath.registers.838[22] [16]),
    .B(\datapath.registers.838[20] [16]),
    .S(\datapath.idinstr_21_bF$buf8 ),
    .Y(_8261_)
);

NAND2X1 _18948_ (
    .A(_7425__bF$buf12),
    .B(_8261_),
    .Y(_8262_)
);

MUX2X1 _18949_ (
    .A(\datapath.registers.838[23] [16]),
    .B(\datapath.registers.838[21] [16]),
    .S(\datapath.idinstr_21_bF$buf7 ),
    .Y(_8263_)
);

NAND2X1 _18950_ (
    .A(\datapath.idinstr_20_bF$buf2 ),
    .B(_8263_),
    .Y(_8264_)
);

NAND3X1 _18951_ (
    .A(\datapath.idinstr_22_bF$buf15 ),
    .B(_8262_),
    .C(_8264_),
    .Y(_8265_)
);

AOI21X1 _18952_ (
    .A(_8260_),
    .B(_8265_),
    .C(\datapath.idinstr_23_bF$buf2 ),
    .Y(_8266_)
);

OAI21X1 _18953_ (
    .A(_8255_),
    .B(_8266_),
    .C(\datapath.idinstr_24_bF$buf1 ),
    .Y(_8267_)
);

AOI22X1 _18954_ (
    .A(_7418__bF$buf3),
    .B(_7422__bF$buf3),
    .C(_8267_),
    .D(_8244_),
    .Y(\datapath.registers.regb_data [16])
);

NAND2X1 _18955_ (
    .A(\datapath.registers.838[27] [17]),
    .B(\datapath.idinstr_20_bF$buf1 ),
    .Y(_8268_)
);

NAND2X1 _18956_ (
    .A(\datapath.registers.838[26] [17]),
    .B(_7425__bF$buf11),
    .Y(_8269_)
);

NAND3X1 _18957_ (
    .A(\datapath.idinstr_21_bF$buf6 ),
    .B(_8268_),
    .C(_8269_),
    .Y(_8270_)
);

NAND2X1 _18958_ (
    .A(\datapath.registers.838[25] [17]),
    .B(\datapath.idinstr_20_bF$buf0 ),
    .Y(_8271_)
);

AOI21X1 _18959_ (
    .A(_7425__bF$buf10),
    .B(\datapath.registers.838[24] [17]),
    .C(\datapath.idinstr_21_bF$buf5 ),
    .Y(_8272_)
);

NAND2X1 _18960_ (
    .A(_8271_),
    .B(_8272_),
    .Y(_8273_)
);

NAND3X1 _18961_ (
    .A(_7420__bF$buf1),
    .B(_8270_),
    .C(_8273_),
    .Y(_8274_)
);

NAND2X1 _18962_ (
    .A(\datapath.registers.838[31] [17]),
    .B(\datapath.idinstr_20_bF$buf55 ),
    .Y(_8275_)
);

AOI21X1 _18963_ (
    .A(_7425__bF$buf9),
    .B(\datapath.registers.838[30] [17]),
    .C(_7419__bF$buf0),
    .Y(_8276_)
);

NAND2X1 _18964_ (
    .A(_8275_),
    .B(_8276_),
    .Y(_8277_)
);

AOI21X1 _18965_ (
    .A(\datapath.registers.838[29] [17]),
    .B(\datapath.idinstr_20_bF$buf54 ),
    .C(\datapath.idinstr_21_bF$buf4 ),
    .Y(_8278_)
);

OAI21X1 _18966_ (
    .A(_6656_),
    .B(\datapath.idinstr_20_bF$buf53 ),
    .C(_8278_),
    .Y(_8279_)
);

NAND3X1 _18967_ (
    .A(\datapath.idinstr_22_bF$buf14 ),
    .B(_8279_),
    .C(_8277_),
    .Y(_8280_)
);

AOI21X1 _18968_ (
    .A(_8274_),
    .B(_8280_),
    .C(_7423__bF$buf5),
    .Y(_8281_)
);

MUX2X1 _18969_ (
    .A(\datapath.registers.838[18] [17]),
    .B(\datapath.registers.838[16] [17]),
    .S(\datapath.idinstr_21_bF$buf3 ),
    .Y(_8282_)
);

NAND2X1 _18970_ (
    .A(_7425__bF$buf8),
    .B(_8282_),
    .Y(_8283_)
);

MUX2X1 _18971_ (
    .A(\datapath.registers.838[19] [17]),
    .B(\datapath.registers.838[17] [17]),
    .S(\datapath.idinstr_21_bF$buf2 ),
    .Y(_8284_)
);

NAND2X1 _18972_ (
    .A(\datapath.idinstr_20_bF$buf52 ),
    .B(_8284_),
    .Y(_8285_)
);

NAND3X1 _18973_ (
    .A(_7420__bF$buf0),
    .B(_8283_),
    .C(_8285_),
    .Y(_8286_)
);

MUX2X1 _18974_ (
    .A(\datapath.registers.838[22] [17]),
    .B(\datapath.registers.838[20] [17]),
    .S(\datapath.idinstr_21_bF$buf1 ),
    .Y(_8287_)
);

NAND2X1 _18975_ (
    .A(_7425__bF$buf7),
    .B(_8287_),
    .Y(_8288_)
);

MUX2X1 _18976_ (
    .A(\datapath.registers.838[23] [17]),
    .B(\datapath.registers.838[21] [17]),
    .S(\datapath.idinstr_21_bF$buf0 ),
    .Y(_8289_)
);

NAND2X1 _18977_ (
    .A(\datapath.idinstr_20_bF$buf51 ),
    .B(_8289_),
    .Y(_8290_)
);

NAND3X1 _18978_ (
    .A(\datapath.idinstr_22_bF$buf13 ),
    .B(_8288_),
    .C(_8290_),
    .Y(_8291_)
);

AOI21X1 _18979_ (
    .A(_8286_),
    .B(_8291_),
    .C(\datapath.idinstr_23_bF$buf1 ),
    .Y(_8292_)
);

OAI21X1 _18980_ (
    .A(_8292_),
    .B(_8281_),
    .C(\datapath.idinstr_24_bF$buf0 ),
    .Y(_8293_)
);

AOI21X1 _18981_ (
    .A(\datapath.registers.838[13] [17]),
    .B(\datapath.idinstr_22_bF$buf12 ),
    .C(_7425__bF$buf6),
    .Y(_8294_)
);

OAI21X1 _18982_ (
    .A(_5287_),
    .B(\datapath.idinstr_22_bF$buf11 ),
    .C(_8294_),
    .Y(_8295_)
);

INVX1 _18983_ (
    .A(\datapath.registers.838[8] [17]),
    .Y(_8296_)
);

AOI21X1 _18984_ (
    .A(\datapath.registers.838[12] [17]),
    .B(\datapath.idinstr_22_bF$buf10 ),
    .C(\datapath.idinstr_20_bF$buf50 ),
    .Y(_8297_)
);

OAI21X1 _18985_ (
    .A(_8296_),
    .B(\datapath.idinstr_22_bF$buf9 ),
    .C(_8297_),
    .Y(_8298_)
);

NAND3X1 _18986_ (
    .A(_7419__bF$buf9),
    .B(_8298_),
    .C(_8295_),
    .Y(_8299_)
);

INVX1 _18987_ (
    .A(\datapath.registers.838[11] [17]),
    .Y(_8300_)
);

AOI21X1 _18988_ (
    .A(\datapath.registers.838[15] [17]),
    .B(\datapath.idinstr_22_bF$buf8 ),
    .C(_7425__bF$buf5),
    .Y(_8301_)
);

OAI21X1 _18989_ (
    .A(_8300_),
    .B(\datapath.idinstr_22_bF$buf7 ),
    .C(_8301_),
    .Y(_8302_)
);

AOI21X1 _18990_ (
    .A(\datapath.registers.838[14] [17]),
    .B(\datapath.idinstr_22_bF$buf6 ),
    .C(\datapath.idinstr_20_bF$buf49 ),
    .Y(_8303_)
);

OAI21X1 _18991_ (
    .A(_5243_),
    .B(\datapath.idinstr_22_bF$buf5 ),
    .C(_8303_),
    .Y(_8304_)
);

NAND3X1 _18992_ (
    .A(\datapath.idinstr_21_bF$buf51 ),
    .B(_8304_),
    .C(_8302_),
    .Y(_8305_)
);

AOI21X1 _18993_ (
    .A(_8299_),
    .B(_8305_),
    .C(_7423__bF$buf4),
    .Y(_8306_)
);

MUX2X1 _18994_ (
    .A(\datapath.registers.838[1] [17]),
    .B(\datapath.registers.838[0] [17]),
    .S(\datapath.idinstr_20_bF$buf48 ),
    .Y(_8307_)
);

NOR2X1 _18995_ (
    .A(\datapath.registers.838[3] [17]),
    .B(_7425__bF$buf4),
    .Y(_8308_)
);

OAI21X1 _18996_ (
    .A(\datapath.registers.838[2] [17]),
    .B(\datapath.idinstr_20_bF$buf47 ),
    .C(\datapath.idinstr_21_bF$buf50 ),
    .Y(_8309_)
);

OAI22X1 _18997_ (
    .A(_8309_),
    .B(_8308_),
    .C(\datapath.idinstr_21_bF$buf49 ),
    .D(_8307_),
    .Y(_8310_)
);

NAND2X1 _18998_ (
    .A(_7420__bF$buf10),
    .B(_8310_),
    .Y(_8311_)
);

MUX2X1 _18999_ (
    .A(\datapath.registers.838[5] [17]),
    .B(\datapath.registers.838[4] [17]),
    .S(\datapath.idinstr_20_bF$buf46 ),
    .Y(_8312_)
);

NOR2X1 _19000_ (
    .A(\datapath.registers.838[7] [17]),
    .B(_7425__bF$buf3),
    .Y(_8313_)
);

OAI21X1 _19001_ (
    .A(\datapath.registers.838[6] [17]),
    .B(\datapath.idinstr_20_bF$buf45 ),
    .C(\datapath.idinstr_21_bF$buf48 ),
    .Y(_8314_)
);

OAI22X1 _19002_ (
    .A(_8314_),
    .B(_8313_),
    .C(\datapath.idinstr_21_bF$buf47 ),
    .D(_8312_),
    .Y(_8315_)
);

NAND2X1 _19003_ (
    .A(\datapath.idinstr_22_bF$buf4 ),
    .B(_8315_),
    .Y(_8316_)
);

AOI21X1 _19004_ (
    .A(_8311_),
    .B(_8316_),
    .C(\datapath.idinstr_23_bF$buf0 ),
    .Y(_8317_)
);

OAI21X1 _19005_ (
    .A(_8306_),
    .B(_8317_),
    .C(_7451__bF$buf2),
    .Y(_8318_)
);

AOI22X1 _19006_ (
    .A(_7418__bF$buf2),
    .B(_7422__bF$buf2),
    .C(_8293_),
    .D(_8318_),
    .Y(\datapath.registers.regb_data [17])
);

NAND2X1 _19007_ (
    .A(\datapath.registers.838[27] [18]),
    .B(\datapath.idinstr_20_bF$buf44 ),
    .Y(_8319_)
);

NAND2X1 _19008_ (
    .A(\datapath.registers.838[26] [18]),
    .B(_7425__bF$buf2),
    .Y(_8320_)
);

NAND3X1 _19009_ (
    .A(\datapath.idinstr_21_bF$buf46 ),
    .B(_8319_),
    .C(_8320_),
    .Y(_8321_)
);

NAND2X1 _19010_ (
    .A(\datapath.registers.838[25] [18]),
    .B(\datapath.idinstr_20_bF$buf43 ),
    .Y(_8322_)
);

AOI21X1 _19011_ (
    .A(_7425__bF$buf1),
    .B(\datapath.registers.838[24] [18]),
    .C(\datapath.idinstr_21_bF$buf45 ),
    .Y(_8323_)
);

NAND2X1 _19012_ (
    .A(_8322_),
    .B(_8323_),
    .Y(_8324_)
);

NAND3X1 _19013_ (
    .A(_7420__bF$buf9),
    .B(_8321_),
    .C(_8324_),
    .Y(_8325_)
);

NAND2X1 _19014_ (
    .A(\datapath.registers.838[31] [18]),
    .B(\datapath.idinstr_20_bF$buf42 ),
    .Y(_8326_)
);

AOI21X1 _19015_ (
    .A(_7425__bF$buf0),
    .B(\datapath.registers.838[30] [18]),
    .C(_7419__bF$buf8),
    .Y(_8327_)
);

NAND2X1 _19016_ (
    .A(_8326_),
    .B(_8327_),
    .Y(_8328_)
);

AOI21X1 _19017_ (
    .A(\datapath.registers.838[29] [18]),
    .B(\datapath.idinstr_20_bF$buf41 ),
    .C(\datapath.idinstr_21_bF$buf44 ),
    .Y(_8329_)
);

OAI21X1 _19018_ (
    .A(_6707_),
    .B(\datapath.idinstr_20_bF$buf40 ),
    .C(_8329_),
    .Y(_8330_)
);

NAND3X1 _19019_ (
    .A(\datapath.idinstr_22_bF$buf3 ),
    .B(_8330_),
    .C(_8328_),
    .Y(_8331_)
);

AOI21X1 _19020_ (
    .A(_8325_),
    .B(_8331_),
    .C(_7423__bF$buf3),
    .Y(_8332_)
);

MUX2X1 _19021_ (
    .A(\datapath.registers.838[18] [18]),
    .B(\datapath.registers.838[16] [18]),
    .S(\datapath.idinstr_21_bF$buf43 ),
    .Y(_8333_)
);

NAND2X1 _19022_ (
    .A(_7425__bF$buf47),
    .B(_8333_),
    .Y(_8334_)
);

MUX2X1 _19023_ (
    .A(\datapath.registers.838[19] [18]),
    .B(\datapath.registers.838[17] [18]),
    .S(\datapath.idinstr_21_bF$buf42 ),
    .Y(_8335_)
);

NAND2X1 _19024_ (
    .A(\datapath.idinstr_20_bF$buf39 ),
    .B(_8335_),
    .Y(_8336_)
);

NAND3X1 _19025_ (
    .A(_7420__bF$buf8),
    .B(_8334_),
    .C(_8336_),
    .Y(_8337_)
);

MUX2X1 _19026_ (
    .A(\datapath.registers.838[22] [18]),
    .B(\datapath.registers.838[20] [18]),
    .S(\datapath.idinstr_21_bF$buf41 ),
    .Y(_8338_)
);

NAND2X1 _19027_ (
    .A(_7425__bF$buf46),
    .B(_8338_),
    .Y(_8339_)
);

MUX2X1 _19028_ (
    .A(\datapath.registers.838[23] [18]),
    .B(\datapath.registers.838[21] [18]),
    .S(\datapath.idinstr_21_bF$buf40 ),
    .Y(_8340_)
);

NAND2X1 _19029_ (
    .A(\datapath.idinstr_20_bF$buf38 ),
    .B(_8340_),
    .Y(_8341_)
);

NAND3X1 _19030_ (
    .A(\datapath.idinstr_22_bF$buf2 ),
    .B(_8339_),
    .C(_8341_),
    .Y(_8342_)
);

AOI21X1 _19031_ (
    .A(_8337_),
    .B(_8342_),
    .C(\datapath.idinstr_23_bF$buf6 ),
    .Y(_8343_)
);

OAI21X1 _19032_ (
    .A(_8343_),
    .B(_8332_),
    .C(\datapath.idinstr_24_bF$buf5 ),
    .Y(_8344_)
);

AOI21X1 _19033_ (
    .A(\datapath.registers.838[13] [18]),
    .B(\datapath.idinstr_22_bF$buf1 ),
    .C(_7425__bF$buf45),
    .Y(_8345_)
);

OAI21X1 _19034_ (
    .A(_5289_),
    .B(\datapath.idinstr_22_bF$buf0 ),
    .C(_8345_),
    .Y(_8346_)
);

INVX1 _19035_ (
    .A(\datapath.registers.838[8] [18]),
    .Y(_8347_)
);

AOI21X1 _19036_ (
    .A(\datapath.registers.838[12] [18]),
    .B(\datapath.idinstr_22_bF$buf41 ),
    .C(\datapath.idinstr_20_bF$buf37 ),
    .Y(_8348_)
);

OAI21X1 _19037_ (
    .A(_8347_),
    .B(\datapath.idinstr_22_bF$buf40 ),
    .C(_8348_),
    .Y(_8349_)
);

NAND3X1 _19038_ (
    .A(_7419__bF$buf7),
    .B(_8349_),
    .C(_8346_),
    .Y(_8350_)
);

INVX1 _19039_ (
    .A(\datapath.registers.838[11] [18]),
    .Y(_8351_)
);

AOI21X1 _19040_ (
    .A(\datapath.registers.838[15] [18]),
    .B(\datapath.idinstr_22_bF$buf39 ),
    .C(_7425__bF$buf44),
    .Y(_8352_)
);

OAI21X1 _19041_ (
    .A(_8351_),
    .B(\datapath.idinstr_22_bF$buf38 ),
    .C(_8352_),
    .Y(_8353_)
);

AOI21X1 _19042_ (
    .A(\datapath.registers.838[14] [18]),
    .B(\datapath.idinstr_22_bF$buf37 ),
    .C(\datapath.idinstr_20_bF$buf36 ),
    .Y(_8354_)
);

OAI21X1 _19043_ (
    .A(_5245_),
    .B(\datapath.idinstr_22_bF$buf36 ),
    .C(_8354_),
    .Y(_8355_)
);

NAND3X1 _19044_ (
    .A(\datapath.idinstr_21_bF$buf39 ),
    .B(_8355_),
    .C(_8353_),
    .Y(_8356_)
);

AOI21X1 _19045_ (
    .A(_8350_),
    .B(_8356_),
    .C(_7423__bF$buf2),
    .Y(_8357_)
);

MUX2X1 _19046_ (
    .A(\datapath.registers.838[1] [18]),
    .B(\datapath.registers.838[0] [18]),
    .S(\datapath.idinstr_20_bF$buf35 ),
    .Y(_8358_)
);

NOR2X1 _19047_ (
    .A(\datapath.registers.838[3] [18]),
    .B(_7425__bF$buf43),
    .Y(_8359_)
);

OAI21X1 _19048_ (
    .A(\datapath.registers.838[2] [18]),
    .B(\datapath.idinstr_20_bF$buf34 ),
    .C(\datapath.idinstr_21_bF$buf38 ),
    .Y(_8360_)
);

OAI22X1 _19049_ (
    .A(_8360_),
    .B(_8359_),
    .C(\datapath.idinstr_21_bF$buf37 ),
    .D(_8358_),
    .Y(_8361_)
);

NAND2X1 _19050_ (
    .A(_7420__bF$buf7),
    .B(_8361_),
    .Y(_8362_)
);

MUX2X1 _19051_ (
    .A(\datapath.registers.838[5] [18]),
    .B(\datapath.registers.838[4] [18]),
    .S(\datapath.idinstr_20_bF$buf33 ),
    .Y(_8363_)
);

NOR2X1 _19052_ (
    .A(\datapath.registers.838[7] [18]),
    .B(_7425__bF$buf42),
    .Y(_8364_)
);

OAI21X1 _19053_ (
    .A(\datapath.registers.838[6] [18]),
    .B(\datapath.idinstr_20_bF$buf32 ),
    .C(\datapath.idinstr_21_bF$buf36 ),
    .Y(_8365_)
);

OAI22X1 _19054_ (
    .A(_8365_),
    .B(_8364_),
    .C(\datapath.idinstr_21_bF$buf35 ),
    .D(_8363_),
    .Y(_8366_)
);

NAND2X1 _19055_ (
    .A(\datapath.idinstr_22_bF$buf35 ),
    .B(_8366_),
    .Y(_8367_)
);

AOI21X1 _19056_ (
    .A(_8362_),
    .B(_8367_),
    .C(\datapath.idinstr_23_bF$buf5 ),
    .Y(_8368_)
);

OAI21X1 _19057_ (
    .A(_8357_),
    .B(_8368_),
    .C(_7451__bF$buf1),
    .Y(_8369_)
);

AOI22X1 _19058_ (
    .A(_7418__bF$buf1),
    .B(_7422__bF$buf1),
    .C(_8344_),
    .D(_8369_),
    .Y(\datapath.registers.regb_data [18])
);

MUX2X1 _19059_ (
    .A(\datapath.registers.838[2] [19]),
    .B(\datapath.registers.838[0] [19]),
    .S(\datapath.idinstr_21_bF$buf34 ),
    .Y(_8370_)
);

NAND2X1 _19060_ (
    .A(_7425__bF$buf41),
    .B(_8370_),
    .Y(_8371_)
);

MUX2X1 _19061_ (
    .A(\datapath.registers.838[3] [19]),
    .B(\datapath.registers.838[1] [19]),
    .S(\datapath.idinstr_21_bF$buf33 ),
    .Y(_8372_)
);

NAND2X1 _19062_ (
    .A(\datapath.idinstr_20_bF$buf31 ),
    .B(_8372_),
    .Y(_8373_)
);

NAND3X1 _19063_ (
    .A(_7420__bF$buf6),
    .B(_8371_),
    .C(_8373_),
    .Y(_8374_)
);

MUX2X1 _19064_ (
    .A(\datapath.registers.838[6] [19]),
    .B(\datapath.registers.838[4] [19]),
    .S(\datapath.idinstr_21_bF$buf32 ),
    .Y(_8375_)
);

NAND2X1 _19065_ (
    .A(_7425__bF$buf40),
    .B(_8375_),
    .Y(_8376_)
);

MUX2X1 _19066_ (
    .A(\datapath.registers.838[7] [19]),
    .B(\datapath.registers.838[5] [19]),
    .S(\datapath.idinstr_21_bF$buf31 ),
    .Y(_8377_)
);

NAND2X1 _19067_ (
    .A(\datapath.idinstr_20_bF$buf30 ),
    .B(_8377_),
    .Y(_8378_)
);

NAND3X1 _19068_ (
    .A(\datapath.idinstr_22_bF$buf34 ),
    .B(_8376_),
    .C(_8378_),
    .Y(_8379_)
);

AOI21X1 _19069_ (
    .A(_8374_),
    .B(_8379_),
    .C(\datapath.idinstr_23_bF$buf4 ),
    .Y(_8380_)
);

AOI21X1 _19070_ (
    .A(\datapath.registers.838[13] [19]),
    .B(\datapath.idinstr_22_bF$buf33 ),
    .C(_7425__bF$buf39),
    .Y(_8381_)
);

OAI21X1 _19071_ (
    .A(_5291_),
    .B(\datapath.idinstr_22_bF$buf32 ),
    .C(_8381_),
    .Y(_8382_)
);

INVX1 _19072_ (
    .A(\datapath.registers.838[8] [19]),
    .Y(_8383_)
);

AOI21X1 _19073_ (
    .A(\datapath.registers.838[12] [19]),
    .B(\datapath.idinstr_22_bF$buf31 ),
    .C(\datapath.idinstr_20_bF$buf29 ),
    .Y(_8384_)
);

OAI21X1 _19074_ (
    .A(_8383_),
    .B(\datapath.idinstr_22_bF$buf30 ),
    .C(_8384_),
    .Y(_8385_)
);

NAND3X1 _19075_ (
    .A(_7419__bF$buf6),
    .B(_8385_),
    .C(_8382_),
    .Y(_8386_)
);

INVX1 _19076_ (
    .A(\datapath.registers.838[11] [19]),
    .Y(_8387_)
);

AOI21X1 _19077_ (
    .A(\datapath.registers.838[15] [19]),
    .B(\datapath.idinstr_22_bF$buf29 ),
    .C(_7425__bF$buf38),
    .Y(_8388_)
);

OAI21X1 _19078_ (
    .A(_8387_),
    .B(\datapath.idinstr_22_bF$buf28 ),
    .C(_8388_),
    .Y(_8389_)
);

AOI21X1 _19079_ (
    .A(\datapath.registers.838[14] [19]),
    .B(\datapath.idinstr_22_bF$buf27 ),
    .C(\datapath.idinstr_20_bF$buf28 ),
    .Y(_8390_)
);

OAI21X1 _19080_ (
    .A(_5247_),
    .B(\datapath.idinstr_22_bF$buf26 ),
    .C(_8390_),
    .Y(_8391_)
);

NAND3X1 _19081_ (
    .A(\datapath.idinstr_21_bF$buf30 ),
    .B(_8391_),
    .C(_8389_),
    .Y(_8392_)
);

AOI21X1 _19082_ (
    .A(_8386_),
    .B(_8392_),
    .C(_7423__bF$buf1),
    .Y(_8393_)
);

OAI21X1 _19083_ (
    .A(_8393_),
    .B(_8380_),
    .C(_7451__bF$buf0),
    .Y(_8394_)
);

NOR2X1 _19084_ (
    .A(\datapath.registers.838[24] [19]),
    .B(\datapath.idinstr_20_bF$buf27 ),
    .Y(_8395_)
);

OAI21X1 _19085_ (
    .A(\datapath.registers.838[25] [19]),
    .B(_7425__bF$buf37),
    .C(_7419__bF$buf5),
    .Y(_8396_)
);

NOR2X1 _19086_ (
    .A(\datapath.registers.838[27] [19]),
    .B(_7425__bF$buf36),
    .Y(_8397_)
);

OAI21X1 _19087_ (
    .A(\datapath.registers.838[26] [19]),
    .B(\datapath.idinstr_20_bF$buf26 ),
    .C(\datapath.idinstr_21_bF$buf29 ),
    .Y(_8398_)
);

OAI22X1 _19088_ (
    .A(_8397_),
    .B(_8398_),
    .C(_8395_),
    .D(_8396_),
    .Y(_8399_)
);

NOR2X1 _19089_ (
    .A(\datapath.idinstr_22_bF$buf25 ),
    .B(_8399_),
    .Y(_8400_)
);

MUX2X1 _19090_ (
    .A(\datapath.registers.838[29] [19]),
    .B(\datapath.registers.838[28] [19]),
    .S(\datapath.idinstr_20_bF$buf25 ),
    .Y(_8401_)
);

NOR2X1 _19091_ (
    .A(\datapath.registers.838[31] [19]),
    .B(_7425__bF$buf35),
    .Y(_8402_)
);

OAI21X1 _19092_ (
    .A(\datapath.registers.838[30] [19]),
    .B(\datapath.idinstr_20_bF$buf24 ),
    .C(\datapath.idinstr_21_bF$buf28 ),
    .Y(_8403_)
);

OAI22X1 _19093_ (
    .A(_8403_),
    .B(_8402_),
    .C(\datapath.idinstr_21_bF$buf27 ),
    .D(_8401_),
    .Y(_8404_)
);

OAI21X1 _19094_ (
    .A(_7420__bF$buf5),
    .B(_8404_),
    .C(\datapath.idinstr_23_bF$buf3 ),
    .Y(_8405_)
);

INVX1 _19095_ (
    .A(\datapath.registers.838[19] [19]),
    .Y(_8406_)
);

AOI21X1 _19096_ (
    .A(\datapath.registers.838[23] [19]),
    .B(\datapath.idinstr_22_bF$buf24 ),
    .C(_7425__bF$buf34),
    .Y(_8407_)
);

OAI21X1 _19097_ (
    .A(_8406_),
    .B(\datapath.idinstr_22_bF$buf23 ),
    .C(_8407_),
    .Y(_8408_)
);

NAND2X1 _19098_ (
    .A(\datapath.registers.838[18] [19]),
    .B(_7420__bF$buf4),
    .Y(_8409_)
);

AOI21X1 _19099_ (
    .A(\datapath.registers.838[22] [19]),
    .B(\datapath.idinstr_22_bF$buf22 ),
    .C(\datapath.idinstr_20_bF$buf23 ),
    .Y(_8410_)
);

AOI21X1 _19100_ (
    .A(_8409_),
    .B(_8410_),
    .C(_7419__bF$buf4),
    .Y(_8411_)
);

AOI21X1 _19101_ (
    .A(\datapath.registers.838[21] [19]),
    .B(\datapath.idinstr_22_bF$buf21 ),
    .C(_7425__bF$buf33),
    .Y(_8412_)
);

OAI21X1 _19102_ (
    .A(_4995_),
    .B(\datapath.idinstr_22_bF$buf20 ),
    .C(_8412_),
    .Y(_8413_)
);

NAND2X1 _19103_ (
    .A(\datapath.registers.838[16] [19]),
    .B(_7420__bF$buf3),
    .Y(_8414_)
);

AOI21X1 _19104_ (
    .A(\datapath.registers.838[20] [19]),
    .B(\datapath.idinstr_22_bF$buf19 ),
    .C(\datapath.idinstr_20_bF$buf22 ),
    .Y(_8415_)
);

AOI21X1 _19105_ (
    .A(_8414_),
    .B(_8415_),
    .C(\datapath.idinstr_21_bF$buf26 ),
    .Y(_8416_)
);

AOI22X1 _19106_ (
    .A(_8411_),
    .B(_8408_),
    .C(_8413_),
    .D(_8416_),
    .Y(_8417_)
);

OAI22X1 _19107_ (
    .A(\datapath.idinstr_23_bF$buf2 ),
    .B(_8417_),
    .C(_8400_),
    .D(_8405_),
    .Y(_8418_)
);

NAND2X1 _19108_ (
    .A(\datapath.idinstr_24_bF$buf4 ),
    .B(_8418_),
    .Y(_8419_)
);

AOI22X1 _19109_ (
    .A(_7418__bF$buf0),
    .B(_7422__bF$buf0),
    .C(_8394_),
    .D(_8419_),
    .Y(\datapath.registers.regb_data [19])
);

NAND2X1 _19110_ (
    .A(\datapath.registers.838[27] [20]),
    .B(\datapath.idinstr_20_bF$buf21 ),
    .Y(_8420_)
);

NAND2X1 _19111_ (
    .A(\datapath.registers.838[26] [20]),
    .B(_7425__bF$buf32),
    .Y(_8421_)
);

NAND3X1 _19112_ (
    .A(\datapath.idinstr_21_bF$buf25 ),
    .B(_8420_),
    .C(_8421_),
    .Y(_8422_)
);

NAND2X1 _19113_ (
    .A(\datapath.registers.838[25] [20]),
    .B(\datapath.idinstr_20_bF$buf20 ),
    .Y(_8423_)
);

AOI21X1 _19114_ (
    .A(_7425__bF$buf31),
    .B(\datapath.registers.838[24] [20]),
    .C(\datapath.idinstr_21_bF$buf24 ),
    .Y(_8424_)
);

NAND2X1 _19115_ (
    .A(_8423_),
    .B(_8424_),
    .Y(_8425_)
);

NAND3X1 _19116_ (
    .A(_7420__bF$buf2),
    .B(_8422_),
    .C(_8425_),
    .Y(_8426_)
);

NAND2X1 _19117_ (
    .A(\datapath.registers.838[31] [20]),
    .B(\datapath.idinstr_20_bF$buf19 ),
    .Y(_8427_)
);

AOI21X1 _19118_ (
    .A(_7425__bF$buf30),
    .B(\datapath.registers.838[30] [20]),
    .C(_7419__bF$buf3),
    .Y(_8428_)
);

NAND2X1 _19119_ (
    .A(_8427_),
    .B(_8428_),
    .Y(_8429_)
);

INVX1 _19120_ (
    .A(\datapath.registers.838[28] [20]),
    .Y(_8430_)
);

AOI21X1 _19121_ (
    .A(\datapath.registers.838[29] [20]),
    .B(\datapath.idinstr_20_bF$buf18 ),
    .C(\datapath.idinstr_21_bF$buf23 ),
    .Y(_8431_)
);

OAI21X1 _19122_ (
    .A(_8430_),
    .B(\datapath.idinstr_20_bF$buf17 ),
    .C(_8431_),
    .Y(_8432_)
);

NAND3X1 _19123_ (
    .A(\datapath.idinstr_22_bF$buf18 ),
    .B(_8432_),
    .C(_8429_),
    .Y(_8433_)
);

AOI21X1 _19124_ (
    .A(_8426_),
    .B(_8433_),
    .C(_7423__bF$buf0),
    .Y(_8434_)
);

MUX2X1 _19125_ (
    .A(\datapath.registers.838[18] [20]),
    .B(\datapath.registers.838[16] [20]),
    .S(\datapath.idinstr_21_bF$buf22 ),
    .Y(_8435_)
);

NAND2X1 _19126_ (
    .A(_7425__bF$buf29),
    .B(_8435_),
    .Y(_8436_)
);

MUX2X1 _19127_ (
    .A(\datapath.registers.838[19] [20]),
    .B(\datapath.registers.838[17] [20]),
    .S(\datapath.idinstr_21_bF$buf21 ),
    .Y(_8437_)
);

NAND2X1 _19128_ (
    .A(\datapath.idinstr_20_bF$buf16 ),
    .B(_8437_),
    .Y(_8438_)
);

NAND3X1 _19129_ (
    .A(_7420__bF$buf1),
    .B(_8436_),
    .C(_8438_),
    .Y(_8439_)
);

MUX2X1 _19130_ (
    .A(\datapath.registers.838[22] [20]),
    .B(\datapath.registers.838[20] [20]),
    .S(\datapath.idinstr_21_bF$buf20 ),
    .Y(_8440_)
);

NAND2X1 _19131_ (
    .A(_7425__bF$buf28),
    .B(_8440_),
    .Y(_8441_)
);

MUX2X1 _19132_ (
    .A(\datapath.registers.838[23] [20]),
    .B(\datapath.registers.838[21] [20]),
    .S(\datapath.idinstr_21_bF$buf19 ),
    .Y(_8442_)
);

NAND2X1 _19133_ (
    .A(\datapath.idinstr_20_bF$buf15 ),
    .B(_8442_),
    .Y(_8443_)
);

NAND3X1 _19134_ (
    .A(\datapath.idinstr_22_bF$buf17 ),
    .B(_8441_),
    .C(_8443_),
    .Y(_8444_)
);

AOI21X1 _19135_ (
    .A(_8439_),
    .B(_8444_),
    .C(\datapath.idinstr_23_bF$buf1 ),
    .Y(_8445_)
);

OAI21X1 _19136_ (
    .A(_8445_),
    .B(_8434_),
    .C(\datapath.idinstr_24_bF$buf3 ),
    .Y(_8446_)
);

MUX2X1 _19137_ (
    .A(\datapath.registers.838[9] [20]),
    .B(\datapath.registers.838[8] [20]),
    .S(\datapath.idinstr_20_bF$buf14 ),
    .Y(_8447_)
);

NOR2X1 _19138_ (
    .A(\datapath.registers.838[11] [20]),
    .B(_7425__bF$buf27),
    .Y(_8448_)
);

OAI21X1 _19139_ (
    .A(\datapath.registers.838[10] [20]),
    .B(\datapath.idinstr_20_bF$buf13 ),
    .C(\datapath.idinstr_21_bF$buf18 ),
    .Y(_8449_)
);

OAI22X1 _19140_ (
    .A(_8449_),
    .B(_8448_),
    .C(\datapath.idinstr_21_bF$buf17 ),
    .D(_8447_),
    .Y(_8450_)
);

AOI21X1 _19141_ (
    .A(_7425__bF$buf26),
    .B(\datapath.registers.838[14] [20]),
    .C(_7419__bF$buf2),
    .Y(_8451_)
);

OAI21X1 _19142_ (
    .A(_6803_),
    .B(_7425__bF$buf25),
    .C(_8451_),
    .Y(_8452_)
);

NAND2X1 _19143_ (
    .A(\datapath.registers.838[12] [20]),
    .B(_7425__bF$buf24),
    .Y(_8453_)
);

AOI21X1 _19144_ (
    .A(\datapath.registers.838[13] [20]),
    .B(\datapath.idinstr_20_bF$buf12 ),
    .C(\datapath.idinstr_21_bF$buf16 ),
    .Y(_8454_)
);

AOI21X1 _19145_ (
    .A(_8453_),
    .B(_8454_),
    .C(_7420__bF$buf0),
    .Y(_8455_)
);

AOI22X1 _19146_ (
    .A(_8452_),
    .B(_8455_),
    .C(_7420__bF$buf10),
    .D(_8450_),
    .Y(_8456_)
);

NOR2X1 _19147_ (
    .A(\datapath.registers.838[0] [20]),
    .B(\datapath.idinstr_20_bF$buf11 ),
    .Y(_8457_)
);

OAI21X1 _19148_ (
    .A(\datapath.registers.838[1] [20]),
    .B(_7425__bF$buf23),
    .C(_7419__bF$buf1),
    .Y(_8458_)
);

NOR2X1 _19149_ (
    .A(\datapath.registers.838[3] [20]),
    .B(_7425__bF$buf22),
    .Y(_8459_)
);

OAI21X1 _19150_ (
    .A(\datapath.registers.838[2] [20]),
    .B(\datapath.idinstr_20_bF$buf10 ),
    .C(\datapath.idinstr_21_bF$buf15 ),
    .Y(_8460_)
);

OAI22X1 _19151_ (
    .A(_8459_),
    .B(_8460_),
    .C(_8457_),
    .D(_8458_),
    .Y(_8461_)
);

NOR2X1 _19152_ (
    .A(\datapath.idinstr_22_bF$buf16 ),
    .B(_8461_),
    .Y(_8462_)
);

MUX2X1 _19153_ (
    .A(\datapath.registers.838[5] [20]),
    .B(\datapath.registers.838[4] [20]),
    .S(\datapath.idinstr_20_bF$buf9 ),
    .Y(_8463_)
);

NOR2X1 _19154_ (
    .A(\datapath.registers.838[7] [20]),
    .B(_7425__bF$buf21),
    .Y(_8464_)
);

OAI21X1 _19155_ (
    .A(\datapath.registers.838[6] [20]),
    .B(\datapath.idinstr_20_bF$buf8 ),
    .C(\datapath.idinstr_21_bF$buf14 ),
    .Y(_8465_)
);

OAI22X1 _19156_ (
    .A(_8465_),
    .B(_8464_),
    .C(\datapath.idinstr_21_bF$buf13 ),
    .D(_8463_),
    .Y(_8466_)
);

OAI21X1 _19157_ (
    .A(_7420__bF$buf9),
    .B(_8466_),
    .C(_7423__bF$buf7),
    .Y(_8467_)
);

OAI22X1 _19158_ (
    .A(_7423__bF$buf6),
    .B(_8456_),
    .C(_8462_),
    .D(_8467_),
    .Y(_8468_)
);

NAND2X1 _19159_ (
    .A(_7451__bF$buf4),
    .B(_8468_),
    .Y(_8469_)
);

AOI22X1 _19160_ (
    .A(_7418__bF$buf4),
    .B(_7422__bF$buf4),
    .C(_8446_),
    .D(_8469_),
    .Y(\datapath.registers.regb_data [20])
);

MUX2X1 _19161_ (
    .A(\datapath.registers.838[9] [21]),
    .B(\datapath.registers.838[8] [21]),
    .S(\datapath.idinstr_20_bF$buf7 ),
    .Y(_8470_)
);

NOR2X1 _19162_ (
    .A(\datapath.registers.838[11] [21]),
    .B(_7425__bF$buf20),
    .Y(_8471_)
);

OAI21X1 _19163_ (
    .A(\datapath.registers.838[10] [21]),
    .B(\datapath.idinstr_20_bF$buf6 ),
    .C(\datapath.idinstr_21_bF$buf12 ),
    .Y(_8472_)
);

OAI22X1 _19164_ (
    .A(_8472_),
    .B(_8471_),
    .C(\datapath.idinstr_21_bF$buf11 ),
    .D(_8470_),
    .Y(_8473_)
);

INVX1 _19165_ (
    .A(\datapath.registers.838[15] [21]),
    .Y(_8474_)
);

AOI21X1 _19166_ (
    .A(_7425__bF$buf19),
    .B(\datapath.registers.838[14] [21]),
    .C(_7419__bF$buf0),
    .Y(_8475_)
);

OAI21X1 _19167_ (
    .A(_8474_),
    .B(_7425__bF$buf18),
    .C(_8475_),
    .Y(_8476_)
);

NAND2X1 _19168_ (
    .A(\datapath.registers.838[12] [21]),
    .B(_7425__bF$buf17),
    .Y(_8477_)
);

AOI21X1 _19169_ (
    .A(\datapath.registers.838[13] [21]),
    .B(\datapath.idinstr_20_bF$buf5 ),
    .C(\datapath.idinstr_21_bF$buf10 ),
    .Y(_8478_)
);

AOI21X1 _19170_ (
    .A(_8477_),
    .B(_8478_),
    .C(_7420__bF$buf8),
    .Y(_8479_)
);

AOI22X1 _19171_ (
    .A(_8476_),
    .B(_8479_),
    .C(_7420__bF$buf7),
    .D(_8473_),
    .Y(_8480_)
);

NOR2X1 _19172_ (
    .A(\datapath.registers.838[0] [21]),
    .B(\datapath.idinstr_20_bF$buf4 ),
    .Y(_8481_)
);

OAI21X1 _19173_ (
    .A(\datapath.registers.838[1] [21]),
    .B(_7425__bF$buf16),
    .C(_7419__bF$buf9),
    .Y(_8482_)
);

NOR2X1 _19174_ (
    .A(\datapath.registers.838[3] [21]),
    .B(_7425__bF$buf15),
    .Y(_8483_)
);

OAI21X1 _19175_ (
    .A(\datapath.registers.838[2] [21]),
    .B(\datapath.idinstr_20_bF$buf3 ),
    .C(\datapath.idinstr_21_bF$buf9 ),
    .Y(_8484_)
);

OAI22X1 _19176_ (
    .A(_8483_),
    .B(_8484_),
    .C(_8481_),
    .D(_8482_),
    .Y(_8485_)
);

NOR2X1 _19177_ (
    .A(\datapath.idinstr_22_bF$buf15 ),
    .B(_8485_),
    .Y(_8486_)
);

MUX2X1 _19178_ (
    .A(\datapath.registers.838[5] [21]),
    .B(\datapath.registers.838[4] [21]),
    .S(\datapath.idinstr_20_bF$buf2 ),
    .Y(_8487_)
);

NOR2X1 _19179_ (
    .A(\datapath.registers.838[7] [21]),
    .B(_7425__bF$buf14),
    .Y(_8488_)
);

OAI21X1 _19180_ (
    .A(\datapath.registers.838[6] [21]),
    .B(\datapath.idinstr_20_bF$buf1 ),
    .C(\datapath.idinstr_21_bF$buf8 ),
    .Y(_8489_)
);

OAI22X1 _19181_ (
    .A(_8489_),
    .B(_8488_),
    .C(\datapath.idinstr_21_bF$buf7 ),
    .D(_8487_),
    .Y(_8490_)
);

OAI21X1 _19182_ (
    .A(_7420__bF$buf6),
    .B(_8490_),
    .C(_7423__bF$buf5),
    .Y(_8491_)
);

OAI22X1 _19183_ (
    .A(_7423__bF$buf4),
    .B(_8480_),
    .C(_8486_),
    .D(_8491_),
    .Y(_8492_)
);

NAND2X1 _19184_ (
    .A(_7451__bF$buf3),
    .B(_8492_),
    .Y(_8493_)
);

INVX1 _19185_ (
    .A(\datapath.registers.838[19] [21]),
    .Y(_8494_)
);

AOI21X1 _19186_ (
    .A(\datapath.registers.838[23] [21]),
    .B(\datapath.idinstr_22_bF$buf14 ),
    .C(_7425__bF$buf13),
    .Y(_8495_)
);

OAI21X1 _19187_ (
    .A(_8494_),
    .B(\datapath.idinstr_22_bF$buf13 ),
    .C(_8495_),
    .Y(_8496_)
);

NAND2X1 _19188_ (
    .A(\datapath.registers.838[18] [21]),
    .B(_7420__bF$buf5),
    .Y(_8497_)
);

AOI21X1 _19189_ (
    .A(\datapath.registers.838[22] [21]),
    .B(\datapath.idinstr_22_bF$buf12 ),
    .C(\datapath.idinstr_20_bF$buf0 ),
    .Y(_8498_)
);

AOI21X1 _19190_ (
    .A(_8497_),
    .B(_8498_),
    .C(_7419__bF$buf8),
    .Y(_8499_)
);

AOI21X1 _19191_ (
    .A(\datapath.registers.838[21] [21]),
    .B(\datapath.idinstr_22_bF$buf11 ),
    .C(_7425__bF$buf12),
    .Y(_8500_)
);

OAI21X1 _19192_ (
    .A(_4998_),
    .B(\datapath.idinstr_22_bF$buf10 ),
    .C(_8500_),
    .Y(_8501_)
);

NAND2X1 _19193_ (
    .A(\datapath.registers.838[16] [21]),
    .B(_7420__bF$buf4),
    .Y(_8502_)
);

AOI21X1 _19194_ (
    .A(\datapath.registers.838[20] [21]),
    .B(\datapath.idinstr_22_bF$buf9 ),
    .C(\datapath.idinstr_20_bF$buf55 ),
    .Y(_8503_)
);

AOI21X1 _19195_ (
    .A(_8502_),
    .B(_8503_),
    .C(\datapath.idinstr_21_bF$buf6 ),
    .Y(_8504_)
);

AOI22X1 _19196_ (
    .A(_8499_),
    .B(_8496_),
    .C(_8501_),
    .D(_8504_),
    .Y(_8505_)
);

NOR2X1 _19197_ (
    .A(\datapath.registers.838[24] [21]),
    .B(\datapath.idinstr_20_bF$buf54 ),
    .Y(_8506_)
);

OAI21X1 _19198_ (
    .A(\datapath.registers.838[25] [21]),
    .B(_7425__bF$buf11),
    .C(_7419__bF$buf7),
    .Y(_8507_)
);

NOR2X1 _19199_ (
    .A(\datapath.registers.838[27] [21]),
    .B(_7425__bF$buf10),
    .Y(_8508_)
);

OAI21X1 _19200_ (
    .A(\datapath.registers.838[26] [21]),
    .B(\datapath.idinstr_20_bF$buf53 ),
    .C(\datapath.idinstr_21_bF$buf5 ),
    .Y(_8509_)
);

OAI22X1 _19201_ (
    .A(_8508_),
    .B(_8509_),
    .C(_8506_),
    .D(_8507_),
    .Y(_8510_)
);

NOR2X1 _19202_ (
    .A(\datapath.idinstr_22_bF$buf8 ),
    .B(_8510_),
    .Y(_8511_)
);

MUX2X1 _19203_ (
    .A(\datapath.registers.838[29] [21]),
    .B(\datapath.registers.838[28] [21]),
    .S(\datapath.idinstr_20_bF$buf52 ),
    .Y(_8512_)
);

NOR2X1 _19204_ (
    .A(\datapath.registers.838[31] [21]),
    .B(_7425__bF$buf9),
    .Y(_8513_)
);

OAI21X1 _19205_ (
    .A(\datapath.registers.838[30] [21]),
    .B(\datapath.idinstr_20_bF$buf51 ),
    .C(\datapath.idinstr_21_bF$buf4 ),
    .Y(_8514_)
);

OAI22X1 _19206_ (
    .A(_8514_),
    .B(_8513_),
    .C(\datapath.idinstr_21_bF$buf3 ),
    .D(_8512_),
    .Y(_8515_)
);

OAI21X1 _19207_ (
    .A(_7420__bF$buf3),
    .B(_8515_),
    .C(\datapath.idinstr_23_bF$buf0 ),
    .Y(_8516_)
);

OAI22X1 _19208_ (
    .A(\datapath.idinstr_23_bF$buf6 ),
    .B(_8505_),
    .C(_8511_),
    .D(_8516_),
    .Y(_8517_)
);

NAND2X1 _19209_ (
    .A(\datapath.idinstr_24_bF$buf2 ),
    .B(_8517_),
    .Y(_8518_)
);

AOI22X1 _19210_ (
    .A(_7418__bF$buf3),
    .B(_7422__bF$buf3),
    .C(_8518_),
    .D(_8493_),
    .Y(\datapath.registers.regb_data [21])
);

MUX2X1 _19211_ (
    .A(\datapath.registers.838[9] [22]),
    .B(\datapath.registers.838[8] [22]),
    .S(\datapath.idinstr_20_bF$buf50 ),
    .Y(_8519_)
);

NOR2X1 _19212_ (
    .A(\datapath.registers.838[11] [22]),
    .B(_7425__bF$buf8),
    .Y(_8520_)
);

OAI21X1 _19213_ (
    .A(\datapath.registers.838[10] [22]),
    .B(\datapath.idinstr_20_bF$buf49 ),
    .C(\datapath.idinstr_21_bF$buf2 ),
    .Y(_8521_)
);

OAI22X1 _19214_ (
    .A(_8521_),
    .B(_8520_),
    .C(\datapath.idinstr_21_bF$buf1 ),
    .D(_8519_),
    .Y(_8522_)
);

AOI21X1 _19215_ (
    .A(_7425__bF$buf7),
    .B(\datapath.registers.838[14] [22]),
    .C(_7419__bF$buf6),
    .Y(_8523_)
);

OAI21X1 _19216_ (
    .A(_6911_),
    .B(_7425__bF$buf6),
    .C(_8523_),
    .Y(_8524_)
);

NAND2X1 _19217_ (
    .A(\datapath.registers.838[12] [22]),
    .B(_7425__bF$buf5),
    .Y(_8525_)
);

AOI21X1 _19218_ (
    .A(\datapath.registers.838[13] [22]),
    .B(\datapath.idinstr_20_bF$buf48 ),
    .C(\datapath.idinstr_21_bF$buf0 ),
    .Y(_8526_)
);

AOI21X1 _19219_ (
    .A(_8525_),
    .B(_8526_),
    .C(_7420__bF$buf2),
    .Y(_8527_)
);

AOI22X1 _19220_ (
    .A(_8524_),
    .B(_8527_),
    .C(_7420__bF$buf1),
    .D(_8522_),
    .Y(_8528_)
);

NOR2X1 _19221_ (
    .A(\datapath.registers.838[0] [22]),
    .B(\datapath.idinstr_20_bF$buf47 ),
    .Y(_8529_)
);

OAI21X1 _19222_ (
    .A(\datapath.registers.838[1] [22]),
    .B(_7425__bF$buf4),
    .C(_7419__bF$buf5),
    .Y(_8530_)
);

NOR2X1 _19223_ (
    .A(\datapath.registers.838[3] [22]),
    .B(_7425__bF$buf3),
    .Y(_8531_)
);

OAI21X1 _19224_ (
    .A(\datapath.registers.838[2] [22]),
    .B(\datapath.idinstr_20_bF$buf46 ),
    .C(\datapath.idinstr_21_bF$buf51 ),
    .Y(_8532_)
);

OAI22X1 _19225_ (
    .A(_8531_),
    .B(_8532_),
    .C(_8529_),
    .D(_8530_),
    .Y(_8533_)
);

NOR2X1 _19226_ (
    .A(\datapath.idinstr_22_bF$buf7 ),
    .B(_8533_),
    .Y(_8534_)
);

MUX2X1 _19227_ (
    .A(\datapath.registers.838[5] [22]),
    .B(\datapath.registers.838[4] [22]),
    .S(\datapath.idinstr_20_bF$buf45 ),
    .Y(_8535_)
);

NOR2X1 _19228_ (
    .A(\datapath.registers.838[7] [22]),
    .B(_7425__bF$buf2),
    .Y(_8536_)
);

OAI21X1 _19229_ (
    .A(\datapath.registers.838[6] [22]),
    .B(\datapath.idinstr_20_bF$buf44 ),
    .C(\datapath.idinstr_21_bF$buf50 ),
    .Y(_8537_)
);

OAI22X1 _19230_ (
    .A(_8537_),
    .B(_8536_),
    .C(\datapath.idinstr_21_bF$buf49 ),
    .D(_8535_),
    .Y(_8538_)
);

OAI21X1 _19231_ (
    .A(_7420__bF$buf0),
    .B(_8538_),
    .C(_7423__bF$buf3),
    .Y(_8539_)
);

OAI22X1 _19232_ (
    .A(_7423__bF$buf2),
    .B(_8528_),
    .C(_8534_),
    .D(_8539_),
    .Y(_8540_)
);

NAND2X1 _19233_ (
    .A(_7451__bF$buf2),
    .B(_8540_),
    .Y(_8541_)
);

INVX1 _19234_ (
    .A(\datapath.registers.838[27] [22]),
    .Y(_8542_)
);

AOI21X1 _19235_ (
    .A(\datapath.registers.838[31] [22]),
    .B(\datapath.idinstr_22_bF$buf6 ),
    .C(_7425__bF$buf1),
    .Y(_8543_)
);

OAI21X1 _19236_ (
    .A(_8542_),
    .B(\datapath.idinstr_22_bF$buf5 ),
    .C(_8543_),
    .Y(_8544_)
);

INVX1 _19237_ (
    .A(\datapath.registers.838[26] [22]),
    .Y(_8545_)
);

AOI21X1 _19238_ (
    .A(\datapath.registers.838[30] [22]),
    .B(\datapath.idinstr_22_bF$buf4 ),
    .C(\datapath.idinstr_20_bF$buf43 ),
    .Y(_8546_)
);

OAI21X1 _19239_ (
    .A(_8545_),
    .B(\datapath.idinstr_22_bF$buf3 ),
    .C(_8546_),
    .Y(_8547_)
);

NAND3X1 _19240_ (
    .A(\datapath.idinstr_21_bF$buf48 ),
    .B(_8547_),
    .C(_8544_),
    .Y(_8548_)
);

INVX1 _19241_ (
    .A(\datapath.registers.838[25] [22]),
    .Y(_8549_)
);

AOI21X1 _19242_ (
    .A(\datapath.registers.838[29] [22]),
    .B(\datapath.idinstr_22_bF$buf2 ),
    .C(_7425__bF$buf0),
    .Y(_8550_)
);

OAI21X1 _19243_ (
    .A(_8549_),
    .B(\datapath.idinstr_22_bF$buf1 ),
    .C(_8550_),
    .Y(_8551_)
);

INVX1 _19244_ (
    .A(\datapath.registers.838[24] [22]),
    .Y(_8552_)
);

AOI21X1 _19245_ (
    .A(\datapath.registers.838[28] [22]),
    .B(\datapath.idinstr_22_bF$buf0 ),
    .C(\datapath.idinstr_20_bF$buf42 ),
    .Y(_8553_)
);

OAI21X1 _19246_ (
    .A(_8552_),
    .B(\datapath.idinstr_22_bF$buf41 ),
    .C(_8553_),
    .Y(_8554_)
);

NAND3X1 _19247_ (
    .A(_7419__bF$buf4),
    .B(_8554_),
    .C(_8551_),
    .Y(_8555_)
);

AOI21X1 _19248_ (
    .A(_8548_),
    .B(_8555_),
    .C(_7423__bF$buf1),
    .Y(_8556_)
);

MUX2X1 _19249_ (
    .A(\datapath.registers.838[18] [22]),
    .B(\datapath.registers.838[16] [22]),
    .S(\datapath.idinstr_21_bF$buf47 ),
    .Y(_8557_)
);

NAND2X1 _19250_ (
    .A(_7425__bF$buf47),
    .B(_8557_),
    .Y(_8558_)
);

MUX2X1 _19251_ (
    .A(\datapath.registers.838[19] [22]),
    .B(\datapath.registers.838[17] [22]),
    .S(\datapath.idinstr_21_bF$buf46 ),
    .Y(_8559_)
);

NAND2X1 _19252_ (
    .A(\datapath.idinstr_20_bF$buf41 ),
    .B(_8559_),
    .Y(_8560_)
);

NAND3X1 _19253_ (
    .A(_7420__bF$buf10),
    .B(_8558_),
    .C(_8560_),
    .Y(_8561_)
);

MUX2X1 _19254_ (
    .A(\datapath.registers.838[22] [22]),
    .B(\datapath.registers.838[20] [22]),
    .S(\datapath.idinstr_21_bF$buf45 ),
    .Y(_8562_)
);

NAND2X1 _19255_ (
    .A(_7425__bF$buf46),
    .B(_8562_),
    .Y(_8563_)
);

MUX2X1 _19256_ (
    .A(\datapath.registers.838[23] [22]),
    .B(\datapath.registers.838[21] [22]),
    .S(\datapath.idinstr_21_bF$buf44 ),
    .Y(_8564_)
);

NAND2X1 _19257_ (
    .A(\datapath.idinstr_20_bF$buf40 ),
    .B(_8564_),
    .Y(_8565_)
);

NAND3X1 _19258_ (
    .A(\datapath.idinstr_22_bF$buf40 ),
    .B(_8563_),
    .C(_8565_),
    .Y(_8566_)
);

AOI21X1 _19259_ (
    .A(_8561_),
    .B(_8566_),
    .C(\datapath.idinstr_23_bF$buf5 ),
    .Y(_8567_)
);

OAI21X1 _19260_ (
    .A(_8556_),
    .B(_8567_),
    .C(\datapath.idinstr_24_bF$buf1 ),
    .Y(_8568_)
);

AOI22X1 _19261_ (
    .A(_7418__bF$buf2),
    .B(_7422__bF$buf2),
    .C(_8568_),
    .D(_8541_),
    .Y(\datapath.registers.regb_data [22])
);

NAND2X1 _19262_ (
    .A(\datapath.registers.838[11] [23]),
    .B(\datapath.idinstr_21_bF$buf43 ),
    .Y(_8569_)
);

NAND2X1 _19263_ (
    .A(\datapath.registers.838[9] [23]),
    .B(_7419__bF$buf3),
    .Y(_8570_)
);

NAND3X1 _19264_ (
    .A(\datapath.idinstr_20_bF$buf39 ),
    .B(_8569_),
    .C(_8570_),
    .Y(_8571_)
);

NAND2X1 _19265_ (
    .A(\datapath.registers.838[10] [23]),
    .B(\datapath.idinstr_21_bF$buf42 ),
    .Y(_8572_)
);

AOI21X1 _19266_ (
    .A(_7419__bF$buf2),
    .B(\datapath.registers.838[8] [23]),
    .C(\datapath.idinstr_20_bF$buf38 ),
    .Y(_8573_)
);

NAND2X1 _19267_ (
    .A(_8572_),
    .B(_8573_),
    .Y(_8574_)
);

NAND3X1 _19268_ (
    .A(_7420__bF$buf9),
    .B(_8571_),
    .C(_8574_),
    .Y(_8575_)
);

NAND2X1 _19269_ (
    .A(\datapath.registers.838[15] [23]),
    .B(\datapath.idinstr_21_bF$buf41 ),
    .Y(_8576_)
);

NAND2X1 _19270_ (
    .A(\datapath.registers.838[13] [23]),
    .B(_7419__bF$buf1),
    .Y(_8577_)
);

NAND3X1 _19271_ (
    .A(\datapath.idinstr_20_bF$buf37 ),
    .B(_8576_),
    .C(_8577_),
    .Y(_8578_)
);

NAND2X1 _19272_ (
    .A(\datapath.registers.838[14] [23]),
    .B(\datapath.idinstr_21_bF$buf40 ),
    .Y(_8579_)
);

AOI21X1 _19273_ (
    .A(_7419__bF$buf0),
    .B(\datapath.registers.838[12] [23]),
    .C(\datapath.idinstr_20_bF$buf36 ),
    .Y(_8580_)
);

NAND2X1 _19274_ (
    .A(_8579_),
    .B(_8580_),
    .Y(_8581_)
);

NAND3X1 _19275_ (
    .A(\datapath.idinstr_22_bF$buf39 ),
    .B(_8578_),
    .C(_8581_),
    .Y(_8582_)
);

AOI21X1 _19276_ (
    .A(_8575_),
    .B(_8582_),
    .C(_7423__bF$buf0),
    .Y(_8583_)
);

INVX1 _19277_ (
    .A(\datapath.registers.838[1] [23]),
    .Y(_8584_)
);

AOI21X1 _19278_ (
    .A(\datapath.registers.838[5] [23]),
    .B(\datapath.idinstr_22_bF$buf38 ),
    .C(_7425__bF$buf45),
    .Y(_8585_)
);

OAI21X1 _19279_ (
    .A(_8584_),
    .B(\datapath.idinstr_22_bF$buf37 ),
    .C(_8585_),
    .Y(_8586_)
);

INVX1 _19280_ (
    .A(\datapath.registers.838[0] [23]),
    .Y(_8587_)
);

AOI21X1 _19281_ (
    .A(\datapath.registers.838[4] [23]),
    .B(\datapath.idinstr_22_bF$buf36 ),
    .C(\datapath.idinstr_20_bF$buf35 ),
    .Y(_8588_)
);

OAI21X1 _19282_ (
    .A(_8587_),
    .B(\datapath.idinstr_22_bF$buf35 ),
    .C(_8588_),
    .Y(_8589_)
);

NAND3X1 _19283_ (
    .A(_7419__bF$buf9),
    .B(_8589_),
    .C(_8586_),
    .Y(_8590_)
);

AOI21X1 _19284_ (
    .A(\datapath.registers.838[7] [23]),
    .B(\datapath.idinstr_22_bF$buf34 ),
    .C(_7425__bF$buf44),
    .Y(_8591_)
);

OAI21X1 _19285_ (
    .A(_5539_),
    .B(\datapath.idinstr_22_bF$buf33 ),
    .C(_8591_),
    .Y(_8592_)
);

INVX1 _19286_ (
    .A(\datapath.registers.838[2] [23]),
    .Y(_8593_)
);

AOI21X1 _19287_ (
    .A(\datapath.registers.838[6] [23]),
    .B(\datapath.idinstr_22_bF$buf32 ),
    .C(\datapath.idinstr_20_bF$buf34 ),
    .Y(_8594_)
);

OAI21X1 _19288_ (
    .A(_8593_),
    .B(\datapath.idinstr_22_bF$buf31 ),
    .C(_8594_),
    .Y(_8595_)
);

NAND3X1 _19289_ (
    .A(\datapath.idinstr_21_bF$buf39 ),
    .B(_8595_),
    .C(_8592_),
    .Y(_8596_)
);

AOI21X1 _19290_ (
    .A(_8590_),
    .B(_8596_),
    .C(\datapath.idinstr_23_bF$buf4 ),
    .Y(_8597_)
);

OAI21X1 _19291_ (
    .A(_8597_),
    .B(_8583_),
    .C(_7451__bF$buf1),
    .Y(_8598_)
);

INVX1 _19292_ (
    .A(\datapath.registers.838[19] [23]),
    .Y(_8599_)
);

AOI21X1 _19293_ (
    .A(\datapath.registers.838[23] [23]),
    .B(\datapath.idinstr_22_bF$buf30 ),
    .C(_7425__bF$buf43),
    .Y(_8600_)
);

OAI21X1 _19294_ (
    .A(_8599_),
    .B(\datapath.idinstr_22_bF$buf29 ),
    .C(_8600_),
    .Y(_8601_)
);

NAND2X1 _19295_ (
    .A(\datapath.registers.838[18] [23]),
    .B(_7420__bF$buf8),
    .Y(_8602_)
);

AOI21X1 _19296_ (
    .A(\datapath.registers.838[22] [23]),
    .B(\datapath.idinstr_22_bF$buf28 ),
    .C(\datapath.idinstr_20_bF$buf33 ),
    .Y(_8603_)
);

AOI21X1 _19297_ (
    .A(_8602_),
    .B(_8603_),
    .C(_7419__bF$buf8),
    .Y(_8604_)
);

AOI21X1 _19298_ (
    .A(\datapath.registers.838[21] [23]),
    .B(\datapath.idinstr_22_bF$buf27 ),
    .C(_7425__bF$buf42),
    .Y(_8605_)
);

OAI21X1 _19299_ (
    .A(_5002_),
    .B(\datapath.idinstr_22_bF$buf26 ),
    .C(_8605_),
    .Y(_8606_)
);

NAND2X1 _19300_ (
    .A(\datapath.registers.838[16] [23]),
    .B(_7420__bF$buf7),
    .Y(_8607_)
);

AOI21X1 _19301_ (
    .A(\datapath.registers.838[20] [23]),
    .B(\datapath.idinstr_22_bF$buf25 ),
    .C(\datapath.idinstr_20_bF$buf32 ),
    .Y(_8608_)
);

AOI21X1 _19302_ (
    .A(_8607_),
    .B(_8608_),
    .C(\datapath.idinstr_21_bF$buf38 ),
    .Y(_8609_)
);

AOI22X1 _19303_ (
    .A(_8604_),
    .B(_8601_),
    .C(_8606_),
    .D(_8609_),
    .Y(_8610_)
);

NOR2X1 _19304_ (
    .A(\datapath.registers.838[24] [23]),
    .B(\datapath.idinstr_20_bF$buf31 ),
    .Y(_8611_)
);

OAI21X1 _19305_ (
    .A(\datapath.registers.838[25] [23]),
    .B(_7425__bF$buf41),
    .C(_7419__bF$buf7),
    .Y(_8612_)
);

NOR2X1 _19306_ (
    .A(\datapath.registers.838[27] [23]),
    .B(_7425__bF$buf40),
    .Y(_8613_)
);

OAI21X1 _19307_ (
    .A(\datapath.registers.838[26] [23]),
    .B(\datapath.idinstr_20_bF$buf30 ),
    .C(\datapath.idinstr_21_bF$buf37 ),
    .Y(_8614_)
);

OAI22X1 _19308_ (
    .A(_8613_),
    .B(_8614_),
    .C(_8611_),
    .D(_8612_),
    .Y(_8615_)
);

NOR2X1 _19309_ (
    .A(\datapath.idinstr_22_bF$buf24 ),
    .B(_8615_),
    .Y(_8616_)
);

MUX2X1 _19310_ (
    .A(\datapath.registers.838[29] [23]),
    .B(\datapath.registers.838[28] [23]),
    .S(\datapath.idinstr_20_bF$buf29 ),
    .Y(_8617_)
);

NOR2X1 _19311_ (
    .A(\datapath.registers.838[31] [23]),
    .B(_7425__bF$buf39),
    .Y(_8618_)
);

OAI21X1 _19312_ (
    .A(\datapath.registers.838[30] [23]),
    .B(\datapath.idinstr_20_bF$buf28 ),
    .C(\datapath.idinstr_21_bF$buf36 ),
    .Y(_8619_)
);

OAI22X1 _19313_ (
    .A(_8619_),
    .B(_8618_),
    .C(\datapath.idinstr_21_bF$buf35 ),
    .D(_8617_),
    .Y(_8620_)
);

OAI21X1 _19314_ (
    .A(_7420__bF$buf6),
    .B(_8620_),
    .C(\datapath.idinstr_23_bF$buf3 ),
    .Y(_8621_)
);

OAI22X1 _19315_ (
    .A(\datapath.idinstr_23_bF$buf2 ),
    .B(_8610_),
    .C(_8616_),
    .D(_8621_),
    .Y(_8622_)
);

NAND2X1 _19316_ (
    .A(\datapath.idinstr_24_bF$buf0 ),
    .B(_8622_),
    .Y(_8623_)
);

AOI22X1 _19317_ (
    .A(_7418__bF$buf1),
    .B(_7422__bF$buf1),
    .C(_8598_),
    .D(_8623_),
    .Y(\datapath.registers.regb_data [23])
);

NAND2X1 _19318_ (
    .A(\datapath.registers.838[27] [24]),
    .B(\datapath.idinstr_20_bF$buf27 ),
    .Y(_8624_)
);

NAND2X1 _19319_ (
    .A(\datapath.registers.838[26] [24]),
    .B(_7425__bF$buf38),
    .Y(_8625_)
);

NAND3X1 _19320_ (
    .A(\datapath.idinstr_21_bF$buf34 ),
    .B(_8624_),
    .C(_8625_),
    .Y(_8626_)
);

NAND2X1 _19321_ (
    .A(\datapath.registers.838[25] [24]),
    .B(\datapath.idinstr_20_bF$buf26 ),
    .Y(_8627_)
);

AOI21X1 _19322_ (
    .A(_7425__bF$buf37),
    .B(\datapath.registers.838[24] [24]),
    .C(\datapath.idinstr_21_bF$buf33 ),
    .Y(_8628_)
);

NAND2X1 _19323_ (
    .A(_8627_),
    .B(_8628_),
    .Y(_8629_)
);

NAND3X1 _19324_ (
    .A(_7420__bF$buf5),
    .B(_8626_),
    .C(_8629_),
    .Y(_8630_)
);

NAND2X1 _19325_ (
    .A(\datapath.registers.838[31] [24]),
    .B(\datapath.idinstr_20_bF$buf25 ),
    .Y(_8631_)
);

AOI21X1 _19326_ (
    .A(_7425__bF$buf36),
    .B(\datapath.registers.838[30] [24]),
    .C(_7419__bF$buf6),
    .Y(_8632_)
);

NAND2X1 _19327_ (
    .A(_8631_),
    .B(_8632_),
    .Y(_8633_)
);

INVX1 _19328_ (
    .A(\datapath.registers.838[28] [24]),
    .Y(_8634_)
);

AOI21X1 _19329_ (
    .A(\datapath.registers.838[29] [24]),
    .B(\datapath.idinstr_20_bF$buf24 ),
    .C(\datapath.idinstr_21_bF$buf32 ),
    .Y(_8635_)
);

OAI21X1 _19330_ (
    .A(_8634_),
    .B(\datapath.idinstr_20_bF$buf23 ),
    .C(_8635_),
    .Y(_8636_)
);

NAND3X1 _19331_ (
    .A(\datapath.idinstr_22_bF$buf23 ),
    .B(_8636_),
    .C(_8633_),
    .Y(_8637_)
);

AOI21X1 _19332_ (
    .A(_8630_),
    .B(_8637_),
    .C(_7423__bF$buf7),
    .Y(_8638_)
);

MUX2X1 _19333_ (
    .A(\datapath.registers.838[17] [24]),
    .B(\datapath.registers.838[16] [24]),
    .S(\datapath.idinstr_20_bF$buf22 ),
    .Y(_8639_)
);

NOR2X1 _19334_ (
    .A(\datapath.registers.838[19] [24]),
    .B(_7425__bF$buf35),
    .Y(_8640_)
);

OAI21X1 _19335_ (
    .A(\datapath.registers.838[18] [24]),
    .B(\datapath.idinstr_20_bF$buf21 ),
    .C(\datapath.idinstr_21_bF$buf31 ),
    .Y(_8641_)
);

OAI22X1 _19336_ (
    .A(_8641_),
    .B(_8640_),
    .C(\datapath.idinstr_21_bF$buf30 ),
    .D(_8639_),
    .Y(_8642_)
);

NAND2X1 _19337_ (
    .A(_7420__bF$buf4),
    .B(_8642_),
    .Y(_8643_)
);

MUX2X1 _19338_ (
    .A(\datapath.registers.838[21] [24]),
    .B(\datapath.registers.838[20] [24]),
    .S(\datapath.idinstr_20_bF$buf20 ),
    .Y(_8644_)
);

NOR2X1 _19339_ (
    .A(\datapath.registers.838[23] [24]),
    .B(_7425__bF$buf34),
    .Y(_8645_)
);

OAI21X1 _19340_ (
    .A(\datapath.registers.838[22] [24]),
    .B(\datapath.idinstr_20_bF$buf19 ),
    .C(\datapath.idinstr_21_bF$buf29 ),
    .Y(_8646_)
);

OAI22X1 _19341_ (
    .A(_8646_),
    .B(_8645_),
    .C(\datapath.idinstr_21_bF$buf28 ),
    .D(_8644_),
    .Y(_8647_)
);

NAND2X1 _19342_ (
    .A(\datapath.idinstr_22_bF$buf22 ),
    .B(_8647_),
    .Y(_8648_)
);

AOI21X1 _19343_ (
    .A(_8643_),
    .B(_8648_),
    .C(\datapath.idinstr_23_bF$buf1 ),
    .Y(_8649_)
);

OAI21X1 _19344_ (
    .A(_8638_),
    .B(_8649_),
    .C(\datapath.idinstr_24_bF$buf5 ),
    .Y(_8650_)
);

NAND2X1 _19345_ (
    .A(\datapath.registers.838[11] [24]),
    .B(\datapath.idinstr_21_bF$buf27 ),
    .Y(_8651_)
);

NAND2X1 _19346_ (
    .A(\datapath.registers.838[9] [24]),
    .B(_7419__bF$buf5),
    .Y(_8652_)
);

NAND3X1 _19347_ (
    .A(\datapath.idinstr_20_bF$buf18 ),
    .B(_8651_),
    .C(_8652_),
    .Y(_8653_)
);

NAND2X1 _19348_ (
    .A(\datapath.registers.838[10] [24]),
    .B(\datapath.idinstr_21_bF$buf26 ),
    .Y(_8654_)
);

AOI21X1 _19349_ (
    .A(_7419__bF$buf4),
    .B(\datapath.registers.838[8] [24]),
    .C(\datapath.idinstr_20_bF$buf17 ),
    .Y(_8655_)
);

NAND2X1 _19350_ (
    .A(_8654_),
    .B(_8655_),
    .Y(_8656_)
);

NAND3X1 _19351_ (
    .A(_7420__bF$buf3),
    .B(_8653_),
    .C(_8656_),
    .Y(_8657_)
);

NAND2X1 _19352_ (
    .A(\datapath.registers.838[15] [24]),
    .B(\datapath.idinstr_21_bF$buf25 ),
    .Y(_8658_)
);

NAND2X1 _19353_ (
    .A(\datapath.registers.838[13] [24]),
    .B(_7419__bF$buf3),
    .Y(_8659_)
);

NAND3X1 _19354_ (
    .A(\datapath.idinstr_20_bF$buf16 ),
    .B(_8658_),
    .C(_8659_),
    .Y(_8660_)
);

NAND2X1 _19355_ (
    .A(\datapath.registers.838[14] [24]),
    .B(\datapath.idinstr_21_bF$buf24 ),
    .Y(_8661_)
);

AOI21X1 _19356_ (
    .A(_7419__bF$buf2),
    .B(\datapath.registers.838[12] [24]),
    .C(\datapath.idinstr_20_bF$buf15 ),
    .Y(_8662_)
);

NAND2X1 _19357_ (
    .A(_8661_),
    .B(_8662_),
    .Y(_8663_)
);

NAND3X1 _19358_ (
    .A(\datapath.idinstr_22_bF$buf21 ),
    .B(_8660_),
    .C(_8663_),
    .Y(_8664_)
);

AOI21X1 _19359_ (
    .A(_8657_),
    .B(_8664_),
    .C(_7423__bF$buf6),
    .Y(_8665_)
);

INVX1 _19360_ (
    .A(\datapath.registers.838[1] [24]),
    .Y(_8666_)
);

AOI21X1 _19361_ (
    .A(\datapath.registers.838[5] [24]),
    .B(\datapath.idinstr_22_bF$buf20 ),
    .C(_7425__bF$buf33),
    .Y(_8667_)
);

OAI21X1 _19362_ (
    .A(_8666_),
    .B(\datapath.idinstr_22_bF$buf19 ),
    .C(_8667_),
    .Y(_8668_)
);

INVX1 _19363_ (
    .A(\datapath.registers.838[0] [24]),
    .Y(_8669_)
);

AOI21X1 _19364_ (
    .A(\datapath.registers.838[4] [24]),
    .B(\datapath.idinstr_22_bF$buf18 ),
    .C(\datapath.idinstr_20_bF$buf14 ),
    .Y(_8670_)
);

OAI21X1 _19365_ (
    .A(_8669_),
    .B(\datapath.idinstr_22_bF$buf17 ),
    .C(_8670_),
    .Y(_8671_)
);

NAND3X1 _19366_ (
    .A(_7419__bF$buf1),
    .B(_8671_),
    .C(_8668_),
    .Y(_8672_)
);

AOI21X1 _19367_ (
    .A(\datapath.registers.838[7] [24]),
    .B(\datapath.idinstr_22_bF$buf16 ),
    .C(_7425__bF$buf32),
    .Y(_8673_)
);

OAI21X1 _19368_ (
    .A(_5541_),
    .B(\datapath.idinstr_22_bF$buf15 ),
    .C(_8673_),
    .Y(_8674_)
);

INVX1 _19369_ (
    .A(\datapath.registers.838[2] [24]),
    .Y(_8675_)
);

AOI21X1 _19370_ (
    .A(\datapath.registers.838[6] [24]),
    .B(\datapath.idinstr_22_bF$buf14 ),
    .C(\datapath.idinstr_20_bF$buf13 ),
    .Y(_8676_)
);

OAI21X1 _19371_ (
    .A(_8675_),
    .B(\datapath.idinstr_22_bF$buf13 ),
    .C(_8676_),
    .Y(_8677_)
);

NAND3X1 _19372_ (
    .A(\datapath.idinstr_21_bF$buf23 ),
    .B(_8677_),
    .C(_8674_),
    .Y(_8678_)
);

AOI21X1 _19373_ (
    .A(_8672_),
    .B(_8678_),
    .C(\datapath.idinstr_23_bF$buf0 ),
    .Y(_8679_)
);

OAI21X1 _19374_ (
    .A(_8679_),
    .B(_8665_),
    .C(_7451__bF$buf0),
    .Y(_8680_)
);

AOI22X1 _19375_ (
    .A(_7418__bF$buf0),
    .B(_7422__bF$buf0),
    .C(_8680_),
    .D(_8650_),
    .Y(\datapath.registers.regb_data [24])
);

MUX2X1 _19376_ (
    .A(\datapath.registers.838[9] [25]),
    .B(\datapath.registers.838[8] [25]),
    .S(\datapath.idinstr_20_bF$buf12 ),
    .Y(_8681_)
);

NOR2X1 _19377_ (
    .A(\datapath.registers.838[11] [25]),
    .B(_7425__bF$buf31),
    .Y(_8682_)
);

OAI21X1 _19378_ (
    .A(\datapath.registers.838[10] [25]),
    .B(\datapath.idinstr_20_bF$buf11 ),
    .C(\datapath.idinstr_21_bF$buf22 ),
    .Y(_8683_)
);

OAI22X1 _19379_ (
    .A(_8683_),
    .B(_8682_),
    .C(\datapath.idinstr_21_bF$buf21 ),
    .D(_8681_),
    .Y(_8684_)
);

INVX1 _19380_ (
    .A(\datapath.registers.838[15] [25]),
    .Y(_8685_)
);

AOI21X1 _19381_ (
    .A(_7425__bF$buf30),
    .B(\datapath.registers.838[14] [25]),
    .C(_7419__bF$buf0),
    .Y(_8686_)
);

OAI21X1 _19382_ (
    .A(_8685_),
    .B(_7425__bF$buf29),
    .C(_8686_),
    .Y(_8687_)
);

NAND2X1 _19383_ (
    .A(\datapath.registers.838[12] [25]),
    .B(_7425__bF$buf28),
    .Y(_8688_)
);

AOI21X1 _19384_ (
    .A(\datapath.registers.838[13] [25]),
    .B(\datapath.idinstr_20_bF$buf10 ),
    .C(\datapath.idinstr_21_bF$buf20 ),
    .Y(_8689_)
);

AOI21X1 _19385_ (
    .A(_8688_),
    .B(_8689_),
    .C(_7420__bF$buf2),
    .Y(_8690_)
);

AOI22X1 _19386_ (
    .A(_8687_),
    .B(_8690_),
    .C(_7420__bF$buf1),
    .D(_8684_),
    .Y(_8691_)
);

NOR2X1 _19387_ (
    .A(\datapath.registers.838[0] [25]),
    .B(\datapath.idinstr_20_bF$buf9 ),
    .Y(_8692_)
);

OAI21X1 _19388_ (
    .A(\datapath.registers.838[1] [25]),
    .B(_7425__bF$buf27),
    .C(_7419__bF$buf9),
    .Y(_8693_)
);

NOR2X1 _19389_ (
    .A(\datapath.registers.838[3] [25]),
    .B(_7425__bF$buf26),
    .Y(_8694_)
);

OAI21X1 _19390_ (
    .A(\datapath.registers.838[2] [25]),
    .B(\datapath.idinstr_20_bF$buf8 ),
    .C(\datapath.idinstr_21_bF$buf19 ),
    .Y(_8695_)
);

OAI22X1 _19391_ (
    .A(_8694_),
    .B(_8695_),
    .C(_8692_),
    .D(_8693_),
    .Y(_8696_)
);

NOR2X1 _19392_ (
    .A(\datapath.idinstr_22_bF$buf12 ),
    .B(_8696_),
    .Y(_8697_)
);

MUX2X1 _19393_ (
    .A(\datapath.registers.838[5] [25]),
    .B(\datapath.registers.838[4] [25]),
    .S(\datapath.idinstr_20_bF$buf7 ),
    .Y(_8698_)
);

NOR2X1 _19394_ (
    .A(\datapath.registers.838[7] [25]),
    .B(_7425__bF$buf25),
    .Y(_8699_)
);

OAI21X1 _19395_ (
    .A(\datapath.registers.838[6] [25]),
    .B(\datapath.idinstr_20_bF$buf6 ),
    .C(\datapath.idinstr_21_bF$buf18 ),
    .Y(_8700_)
);

OAI22X1 _19396_ (
    .A(_8700_),
    .B(_8699_),
    .C(\datapath.idinstr_21_bF$buf17 ),
    .D(_8698_),
    .Y(_8701_)
);

OAI21X1 _19397_ (
    .A(_7420__bF$buf0),
    .B(_8701_),
    .C(_7423__bF$buf5),
    .Y(_8702_)
);

OAI22X1 _19398_ (
    .A(_7423__bF$buf4),
    .B(_8691_),
    .C(_8697_),
    .D(_8702_),
    .Y(_8703_)
);

NAND2X1 _19399_ (
    .A(_7451__bF$buf4),
    .B(_8703_),
    .Y(_8704_)
);

INVX1 _19400_ (
    .A(\datapath.registers.838[19] [25]),
    .Y(_8705_)
);

AOI21X1 _19401_ (
    .A(\datapath.registers.838[23] [25]),
    .B(\datapath.idinstr_22_bF$buf11 ),
    .C(_7425__bF$buf24),
    .Y(_8706_)
);

OAI21X1 _19402_ (
    .A(_8705_),
    .B(\datapath.idinstr_22_bF$buf10 ),
    .C(_8706_),
    .Y(_8707_)
);

NAND2X1 _19403_ (
    .A(\datapath.registers.838[18] [25]),
    .B(_7420__bF$buf10),
    .Y(_8708_)
);

AOI21X1 _19404_ (
    .A(\datapath.registers.838[22] [25]),
    .B(\datapath.idinstr_22_bF$buf9 ),
    .C(\datapath.idinstr_20_bF$buf5 ),
    .Y(_8709_)
);

AOI21X1 _19405_ (
    .A(_8708_),
    .B(_8709_),
    .C(_7419__bF$buf8),
    .Y(_8710_)
);

AOI21X1 _19406_ (
    .A(\datapath.registers.838[21] [25]),
    .B(\datapath.idinstr_22_bF$buf8 ),
    .C(_7425__bF$buf23),
    .Y(_8711_)
);

OAI21X1 _19407_ (
    .A(_5006_),
    .B(\datapath.idinstr_22_bF$buf7 ),
    .C(_8711_),
    .Y(_8712_)
);

NAND2X1 _19408_ (
    .A(\datapath.registers.838[16] [25]),
    .B(_7420__bF$buf9),
    .Y(_8713_)
);

AOI21X1 _19409_ (
    .A(\datapath.registers.838[20] [25]),
    .B(\datapath.idinstr_22_bF$buf6 ),
    .C(\datapath.idinstr_20_bF$buf4 ),
    .Y(_8714_)
);

AOI21X1 _19410_ (
    .A(_8713_),
    .B(_8714_),
    .C(\datapath.idinstr_21_bF$buf16 ),
    .Y(_8715_)
);

AOI22X1 _19411_ (
    .A(_8710_),
    .B(_8707_),
    .C(_8712_),
    .D(_8715_),
    .Y(_8716_)
);

NOR2X1 _19412_ (
    .A(\datapath.registers.838[24] [25]),
    .B(\datapath.idinstr_20_bF$buf3 ),
    .Y(_8717_)
);

OAI21X1 _19413_ (
    .A(\datapath.registers.838[25] [25]),
    .B(_7425__bF$buf22),
    .C(_7419__bF$buf7),
    .Y(_8718_)
);

NOR2X1 _19414_ (
    .A(\datapath.registers.838[27] [25]),
    .B(_7425__bF$buf21),
    .Y(_8719_)
);

OAI21X1 _19415_ (
    .A(\datapath.registers.838[26] [25]),
    .B(\datapath.idinstr_20_bF$buf2 ),
    .C(\datapath.idinstr_21_bF$buf15 ),
    .Y(_8720_)
);

OAI22X1 _19416_ (
    .A(_8719_),
    .B(_8720_),
    .C(_8717_),
    .D(_8718_),
    .Y(_8721_)
);

NOR2X1 _19417_ (
    .A(\datapath.idinstr_22_bF$buf5 ),
    .B(_8721_),
    .Y(_8722_)
);

MUX2X1 _19418_ (
    .A(\datapath.registers.838[29] [25]),
    .B(\datapath.registers.838[28] [25]),
    .S(\datapath.idinstr_20_bF$buf1 ),
    .Y(_8723_)
);

NOR2X1 _19419_ (
    .A(\datapath.registers.838[31] [25]),
    .B(_7425__bF$buf20),
    .Y(_8724_)
);

OAI21X1 _19420_ (
    .A(\datapath.registers.838[30] [25]),
    .B(\datapath.idinstr_20_bF$buf0 ),
    .C(\datapath.idinstr_21_bF$buf14 ),
    .Y(_8725_)
);

OAI22X1 _19421_ (
    .A(_8725_),
    .B(_8724_),
    .C(\datapath.idinstr_21_bF$buf13 ),
    .D(_8723_),
    .Y(_8726_)
);

OAI21X1 _19422_ (
    .A(_7420__bF$buf8),
    .B(_8726_),
    .C(\datapath.idinstr_23_bF$buf6 ),
    .Y(_8727_)
);

OAI22X1 _19423_ (
    .A(\datapath.idinstr_23_bF$buf5 ),
    .B(_8716_),
    .C(_8722_),
    .D(_8727_),
    .Y(_8728_)
);

NAND2X1 _19424_ (
    .A(\datapath.idinstr_24_bF$buf4 ),
    .B(_8728_),
    .Y(_8729_)
);

AOI22X1 _19425_ (
    .A(_7418__bF$buf4),
    .B(_7422__bF$buf4),
    .C(_8729_),
    .D(_8704_),
    .Y(\datapath.registers.regb_data [25])
);

NAND2X1 _19426_ (
    .A(\datapath.registers.838[27] [26]),
    .B(\datapath.idinstr_20_bF$buf55 ),
    .Y(_8730_)
);

NAND2X1 _19427_ (
    .A(\datapath.registers.838[26] [26]),
    .B(_7425__bF$buf19),
    .Y(_8731_)
);

NAND3X1 _19428_ (
    .A(\datapath.idinstr_21_bF$buf12 ),
    .B(_8730_),
    .C(_8731_),
    .Y(_8732_)
);

NAND2X1 _19429_ (
    .A(\datapath.registers.838[25] [26]),
    .B(\datapath.idinstr_20_bF$buf54 ),
    .Y(_8733_)
);

AOI21X1 _19430_ (
    .A(_7425__bF$buf18),
    .B(\datapath.registers.838[24] [26]),
    .C(\datapath.idinstr_21_bF$buf11 ),
    .Y(_8734_)
);

NAND2X1 _19431_ (
    .A(_8733_),
    .B(_8734_),
    .Y(_8735_)
);

NAND3X1 _19432_ (
    .A(_7420__bF$buf7),
    .B(_8732_),
    .C(_8735_),
    .Y(_8736_)
);

NAND2X1 _19433_ (
    .A(\datapath.registers.838[31] [26]),
    .B(\datapath.idinstr_20_bF$buf53 ),
    .Y(_8737_)
);

AOI21X1 _19434_ (
    .A(_7425__bF$buf17),
    .B(\datapath.registers.838[30] [26]),
    .C(_7419__bF$buf6),
    .Y(_8738_)
);

NAND2X1 _19435_ (
    .A(_8737_),
    .B(_8738_),
    .Y(_8739_)
);

AOI21X1 _19436_ (
    .A(\datapath.registers.838[29] [26]),
    .B(\datapath.idinstr_20_bF$buf52 ),
    .C(\datapath.idinstr_21_bF$buf10 ),
    .Y(_8740_)
);

OAI21X1 _19437_ (
    .A(_7124_),
    .B(\datapath.idinstr_20_bF$buf51 ),
    .C(_8740_),
    .Y(_8741_)
);

NAND3X1 _19438_ (
    .A(\datapath.idinstr_22_bF$buf4 ),
    .B(_8741_),
    .C(_8739_),
    .Y(_8742_)
);

AOI21X1 _19439_ (
    .A(_8736_),
    .B(_8742_),
    .C(_7423__bF$buf3),
    .Y(_8743_)
);

MUX2X1 _19440_ (
    .A(\datapath.registers.838[18] [26]),
    .B(\datapath.registers.838[16] [26]),
    .S(\datapath.idinstr_21_bF$buf9 ),
    .Y(_8744_)
);

NAND2X1 _19441_ (
    .A(_7425__bF$buf16),
    .B(_8744_),
    .Y(_8745_)
);

MUX2X1 _19442_ (
    .A(\datapath.registers.838[19] [26]),
    .B(\datapath.registers.838[17] [26]),
    .S(\datapath.idinstr_21_bF$buf8 ),
    .Y(_8746_)
);

NAND2X1 _19443_ (
    .A(\datapath.idinstr_20_bF$buf50 ),
    .B(_8746_),
    .Y(_8747_)
);

NAND3X1 _19444_ (
    .A(_7420__bF$buf6),
    .B(_8745_),
    .C(_8747_),
    .Y(_8748_)
);

MUX2X1 _19445_ (
    .A(\datapath.registers.838[22] [26]),
    .B(\datapath.registers.838[20] [26]),
    .S(\datapath.idinstr_21_bF$buf7 ),
    .Y(_8749_)
);

NAND2X1 _19446_ (
    .A(_7425__bF$buf15),
    .B(_8749_),
    .Y(_8750_)
);

MUX2X1 _19447_ (
    .A(\datapath.registers.838[23] [26]),
    .B(\datapath.registers.838[21] [26]),
    .S(\datapath.idinstr_21_bF$buf6 ),
    .Y(_8751_)
);

NAND2X1 _19448_ (
    .A(\datapath.idinstr_20_bF$buf49 ),
    .B(_8751_),
    .Y(_8752_)
);

NAND3X1 _19449_ (
    .A(\datapath.idinstr_22_bF$buf3 ),
    .B(_8750_),
    .C(_8752_),
    .Y(_8753_)
);

AOI21X1 _19450_ (
    .A(_8748_),
    .B(_8753_),
    .C(\datapath.idinstr_23_bF$buf4 ),
    .Y(_8754_)
);

OAI21X1 _19451_ (
    .A(_8754_),
    .B(_8743_),
    .C(\datapath.idinstr_24_bF$buf3 ),
    .Y(_8755_)
);

MUX2X1 _19452_ (
    .A(\datapath.registers.838[9] [26]),
    .B(\datapath.registers.838[8] [26]),
    .S(\datapath.idinstr_20_bF$buf48 ),
    .Y(_8756_)
);

NOR2X1 _19453_ (
    .A(\datapath.registers.838[11] [26]),
    .B(_7425__bF$buf14),
    .Y(_8757_)
);

OAI21X1 _19454_ (
    .A(\datapath.registers.838[10] [26]),
    .B(\datapath.idinstr_20_bF$buf47 ),
    .C(\datapath.idinstr_21_bF$buf5 ),
    .Y(_8758_)
);

OAI22X1 _19455_ (
    .A(_8758_),
    .B(_8757_),
    .C(\datapath.idinstr_21_bF$buf4 ),
    .D(_8756_),
    .Y(_8759_)
);

AOI21X1 _19456_ (
    .A(_7425__bF$buf13),
    .B(\datapath.registers.838[14] [26]),
    .C(_7419__bF$buf5),
    .Y(_8760_)
);

OAI21X1 _19457_ (
    .A(_7145_),
    .B(_7425__bF$buf12),
    .C(_8760_),
    .Y(_8761_)
);

NAND2X1 _19458_ (
    .A(\datapath.registers.838[12] [26]),
    .B(_7425__bF$buf11),
    .Y(_8762_)
);

AOI21X1 _19459_ (
    .A(\datapath.registers.838[13] [26]),
    .B(\datapath.idinstr_20_bF$buf46 ),
    .C(\datapath.idinstr_21_bF$buf3 ),
    .Y(_8763_)
);

AOI21X1 _19460_ (
    .A(_8762_),
    .B(_8763_),
    .C(_7420__bF$buf5),
    .Y(_8764_)
);

AOI22X1 _19461_ (
    .A(_8761_),
    .B(_8764_),
    .C(_7420__bF$buf4),
    .D(_8759_),
    .Y(_8765_)
);

NOR2X1 _19462_ (
    .A(\datapath.registers.838[0] [26]),
    .B(\datapath.idinstr_20_bF$buf45 ),
    .Y(_8766_)
);

OAI21X1 _19463_ (
    .A(\datapath.registers.838[1] [26]),
    .B(_7425__bF$buf10),
    .C(_7419__bF$buf4),
    .Y(_8767_)
);

NOR2X1 _19464_ (
    .A(\datapath.registers.838[3] [26]),
    .B(_7425__bF$buf9),
    .Y(_8768_)
);

OAI21X1 _19465_ (
    .A(\datapath.registers.838[2] [26]),
    .B(\datapath.idinstr_20_bF$buf44 ),
    .C(\datapath.idinstr_21_bF$buf2 ),
    .Y(_8769_)
);

OAI22X1 _19466_ (
    .A(_8768_),
    .B(_8769_),
    .C(_8766_),
    .D(_8767_),
    .Y(_8770_)
);

NOR2X1 _19467_ (
    .A(\datapath.idinstr_22_bF$buf2 ),
    .B(_8770_),
    .Y(_8771_)
);

MUX2X1 _19468_ (
    .A(\datapath.registers.838[5] [26]),
    .B(\datapath.registers.838[4] [26]),
    .S(\datapath.idinstr_20_bF$buf43 ),
    .Y(_8772_)
);

NOR2X1 _19469_ (
    .A(\datapath.registers.838[7] [26]),
    .B(_7425__bF$buf8),
    .Y(_8773_)
);

OAI21X1 _19470_ (
    .A(\datapath.registers.838[6] [26]),
    .B(\datapath.idinstr_20_bF$buf42 ),
    .C(\datapath.idinstr_21_bF$buf1 ),
    .Y(_8774_)
);

OAI22X1 _19471_ (
    .A(_8774_),
    .B(_8773_),
    .C(\datapath.idinstr_21_bF$buf0 ),
    .D(_8772_),
    .Y(_8775_)
);

OAI21X1 _19472_ (
    .A(_7420__bF$buf3),
    .B(_8775_),
    .C(_7423__bF$buf2),
    .Y(_8776_)
);

OAI22X1 _19473_ (
    .A(_7423__bF$buf1),
    .B(_8765_),
    .C(_8771_),
    .D(_8776_),
    .Y(_8777_)
);

NAND2X1 _19474_ (
    .A(_7451__bF$buf3),
    .B(_8777_),
    .Y(_8778_)
);

AOI22X1 _19475_ (
    .A(_7418__bF$buf3),
    .B(_7422__bF$buf3),
    .C(_8755_),
    .D(_8778_),
    .Y(\datapath.registers.regb_data [26])
);

MUX2X1 _19476_ (
    .A(\datapath.registers.838[9] [27]),
    .B(\datapath.registers.838[8] [27]),
    .S(\datapath.idinstr_20_bF$buf41 ),
    .Y(_8779_)
);

NOR2X1 _19477_ (
    .A(\datapath.registers.838[11] [27]),
    .B(_7425__bF$buf7),
    .Y(_8780_)
);

OAI21X1 _19478_ (
    .A(\datapath.registers.838[10] [27]),
    .B(\datapath.idinstr_20_bF$buf40 ),
    .C(\datapath.idinstr_21_bF$buf51 ),
    .Y(_8781_)
);

OAI22X1 _19479_ (
    .A(_8781_),
    .B(_8780_),
    .C(\datapath.idinstr_21_bF$buf50 ),
    .D(_8779_),
    .Y(_8782_)
);

AOI21X1 _19480_ (
    .A(_7425__bF$buf6),
    .B(\datapath.registers.838[14] [27]),
    .C(_7419__bF$buf3),
    .Y(_8783_)
);

OAI21X1 _19481_ (
    .A(_7169_),
    .B(_7425__bF$buf5),
    .C(_8783_),
    .Y(_8784_)
);

NAND2X1 _19482_ (
    .A(\datapath.registers.838[12] [27]),
    .B(_7425__bF$buf4),
    .Y(_8785_)
);

AOI21X1 _19483_ (
    .A(\datapath.registers.838[13] [27]),
    .B(\datapath.idinstr_20_bF$buf39 ),
    .C(\datapath.idinstr_21_bF$buf49 ),
    .Y(_8786_)
);

AOI21X1 _19484_ (
    .A(_8785_),
    .B(_8786_),
    .C(_7420__bF$buf2),
    .Y(_8787_)
);

AOI22X1 _19485_ (
    .A(_8784_),
    .B(_8787_),
    .C(_7420__bF$buf1),
    .D(_8782_),
    .Y(_8788_)
);

NOR2X1 _19486_ (
    .A(\datapath.registers.838[0] [27]),
    .B(\datapath.idinstr_20_bF$buf38 ),
    .Y(_8789_)
);

OAI21X1 _19487_ (
    .A(\datapath.registers.838[1] [27]),
    .B(_7425__bF$buf3),
    .C(_7419__bF$buf2),
    .Y(_8790_)
);

NOR2X1 _19488_ (
    .A(\datapath.registers.838[3] [27]),
    .B(_7425__bF$buf2),
    .Y(_8791_)
);

OAI21X1 _19489_ (
    .A(\datapath.registers.838[2] [27]),
    .B(\datapath.idinstr_20_bF$buf37 ),
    .C(\datapath.idinstr_21_bF$buf48 ),
    .Y(_8792_)
);

OAI22X1 _19490_ (
    .A(_8791_),
    .B(_8792_),
    .C(_8789_),
    .D(_8790_),
    .Y(_8793_)
);

NOR2X1 _19491_ (
    .A(\datapath.idinstr_22_bF$buf1 ),
    .B(_8793_),
    .Y(_8794_)
);

MUX2X1 _19492_ (
    .A(\datapath.registers.838[5] [27]),
    .B(\datapath.registers.838[4] [27]),
    .S(\datapath.idinstr_20_bF$buf36 ),
    .Y(_8795_)
);

NOR2X1 _19493_ (
    .A(\datapath.registers.838[7] [27]),
    .B(_7425__bF$buf1),
    .Y(_8796_)
);

OAI21X1 _19494_ (
    .A(\datapath.registers.838[6] [27]),
    .B(\datapath.idinstr_20_bF$buf35 ),
    .C(\datapath.idinstr_21_bF$buf47 ),
    .Y(_8797_)
);

OAI22X1 _19495_ (
    .A(_8797_),
    .B(_8796_),
    .C(\datapath.idinstr_21_bF$buf46 ),
    .D(_8795_),
    .Y(_8798_)
);

OAI21X1 _19496_ (
    .A(_7420__bF$buf0),
    .B(_8798_),
    .C(_7423__bF$buf0),
    .Y(_8799_)
);

OAI22X1 _19497_ (
    .A(_7423__bF$buf7),
    .B(_8788_),
    .C(_8794_),
    .D(_8799_),
    .Y(_8800_)
);

NAND2X1 _19498_ (
    .A(_7451__bF$buf2),
    .B(_8800_),
    .Y(_8801_)
);

AOI21X1 _19499_ (
    .A(\datapath.registers.838[23] [27]),
    .B(\datapath.idinstr_22_bF$buf0 ),
    .C(_7425__bF$buf0),
    .Y(_8802_)
);

OAI21X1 _19500_ (
    .A(_7189_),
    .B(\datapath.idinstr_22_bF$buf41 ),
    .C(_8802_),
    .Y(_8803_)
);

NAND2X1 _19501_ (
    .A(\datapath.registers.838[18] [27]),
    .B(_7420__bF$buf10),
    .Y(_8804_)
);

AOI21X1 _19502_ (
    .A(\datapath.registers.838[22] [27]),
    .B(\datapath.idinstr_22_bF$buf40 ),
    .C(\datapath.idinstr_20_bF$buf34 ),
    .Y(_8805_)
);

AOI21X1 _19503_ (
    .A(_8804_),
    .B(_8805_),
    .C(_7419__bF$buf1),
    .Y(_8806_)
);

AOI21X1 _19504_ (
    .A(\datapath.registers.838[21] [27]),
    .B(\datapath.idinstr_22_bF$buf39 ),
    .C(_7425__bF$buf47),
    .Y(_8807_)
);

OAI21X1 _19505_ (
    .A(_5009_),
    .B(\datapath.idinstr_22_bF$buf38 ),
    .C(_8807_),
    .Y(_8808_)
);

NAND2X1 _19506_ (
    .A(\datapath.registers.838[16] [27]),
    .B(_7420__bF$buf9),
    .Y(_8809_)
);

AOI21X1 _19507_ (
    .A(\datapath.registers.838[20] [27]),
    .B(\datapath.idinstr_22_bF$buf37 ),
    .C(\datapath.idinstr_20_bF$buf33 ),
    .Y(_8810_)
);

AOI21X1 _19508_ (
    .A(_8809_),
    .B(_8810_),
    .C(\datapath.idinstr_21_bF$buf45 ),
    .Y(_8811_)
);

AOI22X1 _19509_ (
    .A(_8806_),
    .B(_8803_),
    .C(_8808_),
    .D(_8811_),
    .Y(_8812_)
);

NOR2X1 _19510_ (
    .A(\datapath.registers.838[24] [27]),
    .B(\datapath.idinstr_20_bF$buf32 ),
    .Y(_8813_)
);

OAI21X1 _19511_ (
    .A(\datapath.registers.838[25] [27]),
    .B(_7425__bF$buf46),
    .C(_7419__bF$buf0),
    .Y(_8814_)
);

NOR2X1 _19512_ (
    .A(\datapath.registers.838[27] [27]),
    .B(_7425__bF$buf45),
    .Y(_8815_)
);

OAI21X1 _19513_ (
    .A(\datapath.registers.838[26] [27]),
    .B(\datapath.idinstr_20_bF$buf31 ),
    .C(\datapath.idinstr_21_bF$buf44 ),
    .Y(_8816_)
);

OAI22X1 _19514_ (
    .A(_8815_),
    .B(_8816_),
    .C(_8813_),
    .D(_8814_),
    .Y(_8817_)
);

NOR2X1 _19515_ (
    .A(\datapath.idinstr_22_bF$buf36 ),
    .B(_8817_),
    .Y(_8818_)
);

MUX2X1 _19516_ (
    .A(\datapath.registers.838[29] [27]),
    .B(\datapath.registers.838[28] [27]),
    .S(\datapath.idinstr_20_bF$buf30 ),
    .Y(_8819_)
);

NOR2X1 _19517_ (
    .A(\datapath.registers.838[31] [27]),
    .B(_7425__bF$buf44),
    .Y(_8820_)
);

OAI21X1 _19518_ (
    .A(\datapath.registers.838[30] [27]),
    .B(\datapath.idinstr_20_bF$buf29 ),
    .C(\datapath.idinstr_21_bF$buf43 ),
    .Y(_8821_)
);

OAI22X1 _19519_ (
    .A(_8821_),
    .B(_8820_),
    .C(\datapath.idinstr_21_bF$buf42 ),
    .D(_8819_),
    .Y(_8822_)
);

OAI21X1 _19520_ (
    .A(_7420__bF$buf8),
    .B(_8822_),
    .C(\datapath.idinstr_23_bF$buf3 ),
    .Y(_8823_)
);

OAI22X1 _19521_ (
    .A(\datapath.idinstr_23_bF$buf2 ),
    .B(_8812_),
    .C(_8818_),
    .D(_8823_),
    .Y(_8824_)
);

NAND2X1 _19522_ (
    .A(\datapath.idinstr_24_bF$buf2 ),
    .B(_8824_),
    .Y(_8825_)
);

AOI22X1 _19523_ (
    .A(_7418__bF$buf2),
    .B(_7422__bF$buf2),
    .C(_8825_),
    .D(_8801_),
    .Y(\datapath.registers.regb_data [27])
);

NAND2X1 _19524_ (
    .A(\datapath.registers.838[27] [28]),
    .B(\datapath.idinstr_20_bF$buf28 ),
    .Y(_8826_)
);

NAND2X1 _19525_ (
    .A(\datapath.registers.838[26] [28]),
    .B(_7425__bF$buf43),
    .Y(_8827_)
);

NAND3X1 _19526_ (
    .A(\datapath.idinstr_21_bF$buf41 ),
    .B(_8826_),
    .C(_8827_),
    .Y(_8828_)
);

NAND2X1 _19527_ (
    .A(\datapath.registers.838[25] [28]),
    .B(\datapath.idinstr_20_bF$buf27 ),
    .Y(_8829_)
);

AOI21X1 _19528_ (
    .A(_7425__bF$buf42),
    .B(\datapath.registers.838[24] [28]),
    .C(\datapath.idinstr_21_bF$buf40 ),
    .Y(_8830_)
);

NAND2X1 _19529_ (
    .A(_8829_),
    .B(_8830_),
    .Y(_8831_)
);

NAND3X1 _19530_ (
    .A(_7420__bF$buf7),
    .B(_8828_),
    .C(_8831_),
    .Y(_8832_)
);

NAND2X1 _19531_ (
    .A(\datapath.registers.838[31] [28]),
    .B(\datapath.idinstr_20_bF$buf26 ),
    .Y(_8833_)
);

AOI21X1 _19532_ (
    .A(_7425__bF$buf41),
    .B(\datapath.registers.838[30] [28]),
    .C(_7419__bF$buf9),
    .Y(_8834_)
);

NAND2X1 _19533_ (
    .A(_8833_),
    .B(_8834_),
    .Y(_8835_)
);

INVX1 _19534_ (
    .A(\datapath.registers.838[28] [28]),
    .Y(_8836_)
);

AOI21X1 _19535_ (
    .A(\datapath.registers.838[29] [28]),
    .B(\datapath.idinstr_20_bF$buf25 ),
    .C(\datapath.idinstr_21_bF$buf39 ),
    .Y(_8837_)
);

OAI21X1 _19536_ (
    .A(_8836_),
    .B(\datapath.idinstr_20_bF$buf24 ),
    .C(_8837_),
    .Y(_8838_)
);

NAND3X1 _19537_ (
    .A(\datapath.idinstr_22_bF$buf35 ),
    .B(_8838_),
    .C(_8835_),
    .Y(_8839_)
);

AOI21X1 _19538_ (
    .A(_8832_),
    .B(_8839_),
    .C(_7423__bF$buf6),
    .Y(_8840_)
);

MUX2X1 _19539_ (
    .A(\datapath.registers.838[18] [28]),
    .B(\datapath.registers.838[16] [28]),
    .S(\datapath.idinstr_21_bF$buf38 ),
    .Y(_8841_)
);

NAND2X1 _19540_ (
    .A(_7425__bF$buf40),
    .B(_8841_),
    .Y(_8842_)
);

MUX2X1 _19541_ (
    .A(\datapath.registers.838[19] [28]),
    .B(\datapath.registers.838[17] [28]),
    .S(\datapath.idinstr_21_bF$buf37 ),
    .Y(_8843_)
);

NAND2X1 _19542_ (
    .A(\datapath.idinstr_20_bF$buf23 ),
    .B(_8843_),
    .Y(_8844_)
);

NAND3X1 _19543_ (
    .A(_7420__bF$buf6),
    .B(_8842_),
    .C(_8844_),
    .Y(_8845_)
);

MUX2X1 _19544_ (
    .A(\datapath.registers.838[22] [28]),
    .B(\datapath.registers.838[20] [28]),
    .S(\datapath.idinstr_21_bF$buf36 ),
    .Y(_8846_)
);

NAND2X1 _19545_ (
    .A(_7425__bF$buf39),
    .B(_8846_),
    .Y(_8847_)
);

MUX2X1 _19546_ (
    .A(\datapath.registers.838[23] [28]),
    .B(\datapath.registers.838[21] [28]),
    .S(\datapath.idinstr_21_bF$buf35 ),
    .Y(_8848_)
);

NAND2X1 _19547_ (
    .A(\datapath.idinstr_20_bF$buf22 ),
    .B(_8848_),
    .Y(_8849_)
);

NAND3X1 _19548_ (
    .A(\datapath.idinstr_22_bF$buf34 ),
    .B(_8847_),
    .C(_8849_),
    .Y(_8850_)
);

AOI21X1 _19549_ (
    .A(_8845_),
    .B(_8850_),
    .C(\datapath.idinstr_23_bF$buf1 ),
    .Y(_8851_)
);

OAI21X1 _19550_ (
    .A(_8851_),
    .B(_8840_),
    .C(\datapath.idinstr_24_bF$buf1 ),
    .Y(_8852_)
);

MUX2X1 _19551_ (
    .A(\datapath.registers.838[9] [28]),
    .B(\datapath.registers.838[8] [28]),
    .S(\datapath.idinstr_20_bF$buf21 ),
    .Y(_8853_)
);

NOR2X1 _19552_ (
    .A(\datapath.registers.838[11] [28]),
    .B(_7425__bF$buf38),
    .Y(_8854_)
);

OAI21X1 _19553_ (
    .A(\datapath.registers.838[10] [28]),
    .B(\datapath.idinstr_20_bF$buf20 ),
    .C(\datapath.idinstr_21_bF$buf34 ),
    .Y(_8855_)
);

OAI22X1 _19554_ (
    .A(_8855_),
    .B(_8854_),
    .C(\datapath.idinstr_21_bF$buf33 ),
    .D(_8853_),
    .Y(_8856_)
);

AOI21X1 _19555_ (
    .A(_7425__bF$buf37),
    .B(\datapath.registers.838[14] [28]),
    .C(_7419__bF$buf8),
    .Y(_8857_)
);

OAI21X1 _19556_ (
    .A(_7218_),
    .B(_7425__bF$buf36),
    .C(_8857_),
    .Y(_8858_)
);

NAND2X1 _19557_ (
    .A(\datapath.registers.838[12] [28]),
    .B(_7425__bF$buf35),
    .Y(_8859_)
);

AOI21X1 _19558_ (
    .A(\datapath.registers.838[13] [28]),
    .B(\datapath.idinstr_20_bF$buf19 ),
    .C(\datapath.idinstr_21_bF$buf32 ),
    .Y(_8860_)
);

AOI21X1 _19559_ (
    .A(_8859_),
    .B(_8860_),
    .C(_7420__bF$buf5),
    .Y(_8861_)
);

AOI22X1 _19560_ (
    .A(_8858_),
    .B(_8861_),
    .C(_7420__bF$buf4),
    .D(_8856_),
    .Y(_8862_)
);

NOR2X1 _19561_ (
    .A(\datapath.registers.838[0] [28]),
    .B(\datapath.idinstr_20_bF$buf18 ),
    .Y(_8863_)
);

OAI21X1 _19562_ (
    .A(\datapath.registers.838[1] [28]),
    .B(_7425__bF$buf34),
    .C(_7419__bF$buf7),
    .Y(_8864_)
);

NOR2X1 _19563_ (
    .A(\datapath.registers.838[3] [28]),
    .B(_7425__bF$buf33),
    .Y(_8865_)
);

OAI21X1 _19564_ (
    .A(\datapath.registers.838[2] [28]),
    .B(\datapath.idinstr_20_bF$buf17 ),
    .C(\datapath.idinstr_21_bF$buf31 ),
    .Y(_8866_)
);

OAI22X1 _19565_ (
    .A(_8865_),
    .B(_8866_),
    .C(_8863_),
    .D(_8864_),
    .Y(_8867_)
);

NOR2X1 _19566_ (
    .A(\datapath.idinstr_22_bF$buf33 ),
    .B(_8867_),
    .Y(_8868_)
);

MUX2X1 _19567_ (
    .A(\datapath.registers.838[5] [28]),
    .B(\datapath.registers.838[4] [28]),
    .S(\datapath.idinstr_20_bF$buf16 ),
    .Y(_8869_)
);

NOR2X1 _19568_ (
    .A(\datapath.registers.838[7] [28]),
    .B(_7425__bF$buf32),
    .Y(_8870_)
);

OAI21X1 _19569_ (
    .A(\datapath.registers.838[6] [28]),
    .B(\datapath.idinstr_20_bF$buf15 ),
    .C(\datapath.idinstr_21_bF$buf30 ),
    .Y(_8871_)
);

OAI22X1 _19570_ (
    .A(_8871_),
    .B(_8870_),
    .C(\datapath.idinstr_21_bF$buf29 ),
    .D(_8869_),
    .Y(_8872_)
);

OAI21X1 _19571_ (
    .A(_7420__bF$buf3),
    .B(_8872_),
    .C(_7423__bF$buf5),
    .Y(_8873_)
);

OAI22X1 _19572_ (
    .A(_7423__bF$buf4),
    .B(_8862_),
    .C(_8868_),
    .D(_8873_),
    .Y(_8874_)
);

NAND2X1 _19573_ (
    .A(_7451__bF$buf1),
    .B(_8874_),
    .Y(_8875_)
);

AOI22X1 _19574_ (
    .A(_7418__bF$buf1),
    .B(_7422__bF$buf1),
    .C(_8852_),
    .D(_8875_),
    .Y(\datapath.registers.regb_data [28])
);

NAND2X1 _19575_ (
    .A(\datapath.registers.838[27] [29]),
    .B(\datapath.idinstr_20_bF$buf14 ),
    .Y(_8876_)
);

NAND2X1 _19576_ (
    .A(\datapath.registers.838[26] [29]),
    .B(_7425__bF$buf31),
    .Y(_8877_)
);

NAND3X1 _19577_ (
    .A(\datapath.idinstr_21_bF$buf28 ),
    .B(_8876_),
    .C(_8877_),
    .Y(_8878_)
);

NAND2X1 _19578_ (
    .A(\datapath.registers.838[25] [29]),
    .B(\datapath.idinstr_20_bF$buf13 ),
    .Y(_8879_)
);

AOI21X1 _19579_ (
    .A(_7425__bF$buf30),
    .B(\datapath.registers.838[24] [29]),
    .C(\datapath.idinstr_21_bF$buf27 ),
    .Y(_8880_)
);

NAND2X1 _19580_ (
    .A(_8879_),
    .B(_8880_),
    .Y(_8881_)
);

NAND3X1 _19581_ (
    .A(_7420__bF$buf2),
    .B(_8878_),
    .C(_8881_),
    .Y(_8882_)
);

NAND2X1 _19582_ (
    .A(\datapath.registers.838[31] [29]),
    .B(\datapath.idinstr_20_bF$buf12 ),
    .Y(_8883_)
);

AOI21X1 _19583_ (
    .A(_7425__bF$buf29),
    .B(\datapath.registers.838[30] [29]),
    .C(_7419__bF$buf6),
    .Y(_8884_)
);

NAND2X1 _19584_ (
    .A(_8883_),
    .B(_8884_),
    .Y(_8885_)
);

AOI21X1 _19585_ (
    .A(\datapath.registers.838[29] [29]),
    .B(\datapath.idinstr_20_bF$buf11 ),
    .C(\datapath.idinstr_21_bF$buf26 ),
    .Y(_8886_)
);

OAI21X1 _19586_ (
    .A(_7275_),
    .B(\datapath.idinstr_20_bF$buf10 ),
    .C(_8886_),
    .Y(_8887_)
);

NAND3X1 _19587_ (
    .A(\datapath.idinstr_22_bF$buf32 ),
    .B(_8887_),
    .C(_8885_),
    .Y(_8888_)
);

AOI21X1 _19588_ (
    .A(_8882_),
    .B(_8888_),
    .C(_7423__bF$buf3),
    .Y(_8889_)
);

MUX2X1 _19589_ (
    .A(\datapath.registers.838[18] [29]),
    .B(\datapath.registers.838[16] [29]),
    .S(\datapath.idinstr_21_bF$buf25 ),
    .Y(_8890_)
);

NAND2X1 _19590_ (
    .A(_7425__bF$buf28),
    .B(_8890_),
    .Y(_8891_)
);

MUX2X1 _19591_ (
    .A(\datapath.registers.838[19] [29]),
    .B(\datapath.registers.838[17] [29]),
    .S(\datapath.idinstr_21_bF$buf24 ),
    .Y(_8892_)
);

NAND2X1 _19592_ (
    .A(\datapath.idinstr_20_bF$buf9 ),
    .B(_8892_),
    .Y(_8893_)
);

NAND3X1 _19593_ (
    .A(_7420__bF$buf1),
    .B(_8891_),
    .C(_8893_),
    .Y(_8894_)
);

MUX2X1 _19594_ (
    .A(\datapath.registers.838[22] [29]),
    .B(\datapath.registers.838[20] [29]),
    .S(\datapath.idinstr_21_bF$buf23 ),
    .Y(_8895_)
);

NAND2X1 _19595_ (
    .A(_7425__bF$buf27),
    .B(_8895_),
    .Y(_8896_)
);

MUX2X1 _19596_ (
    .A(\datapath.registers.838[23] [29]),
    .B(\datapath.registers.838[21] [29]),
    .S(\datapath.idinstr_21_bF$buf22 ),
    .Y(_8897_)
);

NAND2X1 _19597_ (
    .A(\datapath.idinstr_20_bF$buf8 ),
    .B(_8897_),
    .Y(_8898_)
);

NAND3X1 _19598_ (
    .A(\datapath.idinstr_22_bF$buf31 ),
    .B(_8896_),
    .C(_8898_),
    .Y(_8899_)
);

AOI21X1 _19599_ (
    .A(_8894_),
    .B(_8899_),
    .C(\datapath.idinstr_23_bF$buf0 ),
    .Y(_8900_)
);

OAI21X1 _19600_ (
    .A(_8900_),
    .B(_8889_),
    .C(\datapath.idinstr_24_bF$buf0 ),
    .Y(_8901_)
);

MUX2X1 _19601_ (
    .A(\datapath.registers.838[9] [29]),
    .B(\datapath.registers.838[8] [29]),
    .S(\datapath.idinstr_20_bF$buf7 ),
    .Y(_8902_)
);

NOR2X1 _19602_ (
    .A(\datapath.registers.838[11] [29]),
    .B(_7425__bF$buf26),
    .Y(_8903_)
);

OAI21X1 _19603_ (
    .A(\datapath.registers.838[10] [29]),
    .B(\datapath.idinstr_20_bF$buf6 ),
    .C(\datapath.idinstr_21_bF$buf21 ),
    .Y(_8904_)
);

OAI22X1 _19604_ (
    .A(_8904_),
    .B(_8903_),
    .C(\datapath.idinstr_21_bF$buf20 ),
    .D(_8902_),
    .Y(_8905_)
);

AOI21X1 _19605_ (
    .A(_7425__bF$buf25),
    .B(\datapath.registers.838[14] [29]),
    .C(_7419__bF$buf5),
    .Y(_8906_)
);

OAI21X1 _19606_ (
    .A(_7296_),
    .B(_7425__bF$buf24),
    .C(_8906_),
    .Y(_8907_)
);

NAND2X1 _19607_ (
    .A(\datapath.registers.838[12] [29]),
    .B(_7425__bF$buf23),
    .Y(_8908_)
);

AOI21X1 _19608_ (
    .A(\datapath.registers.838[13] [29]),
    .B(\datapath.idinstr_20_bF$buf5 ),
    .C(\datapath.idinstr_21_bF$buf19 ),
    .Y(_8909_)
);

AOI21X1 _19609_ (
    .A(_8908_),
    .B(_8909_),
    .C(_7420__bF$buf0),
    .Y(_8910_)
);

AOI22X1 _19610_ (
    .A(_8907_),
    .B(_8910_),
    .C(_7420__bF$buf10),
    .D(_8905_),
    .Y(_8911_)
);

NOR2X1 _19611_ (
    .A(\datapath.registers.838[0] [29]),
    .B(\datapath.idinstr_20_bF$buf4 ),
    .Y(_8912_)
);

OAI21X1 _19612_ (
    .A(\datapath.registers.838[1] [29]),
    .B(_7425__bF$buf22),
    .C(_7419__bF$buf4),
    .Y(_8913_)
);

NOR2X1 _19613_ (
    .A(\datapath.registers.838[3] [29]),
    .B(_7425__bF$buf21),
    .Y(_8914_)
);

OAI21X1 _19614_ (
    .A(\datapath.registers.838[2] [29]),
    .B(\datapath.idinstr_20_bF$buf3 ),
    .C(\datapath.idinstr_21_bF$buf18 ),
    .Y(_8915_)
);

OAI22X1 _19615_ (
    .A(_8914_),
    .B(_8915_),
    .C(_8912_),
    .D(_8913_),
    .Y(_8916_)
);

NOR2X1 _19616_ (
    .A(\datapath.idinstr_22_bF$buf30 ),
    .B(_8916_),
    .Y(_8917_)
);

MUX2X1 _19617_ (
    .A(\datapath.registers.838[5] [29]),
    .B(\datapath.registers.838[4] [29]),
    .S(\datapath.idinstr_20_bF$buf2 ),
    .Y(_8918_)
);

NOR2X1 _19618_ (
    .A(\datapath.registers.838[7] [29]),
    .B(_7425__bF$buf20),
    .Y(_8919_)
);

OAI21X1 _19619_ (
    .A(\datapath.registers.838[6] [29]),
    .B(\datapath.idinstr_20_bF$buf1 ),
    .C(\datapath.idinstr_21_bF$buf17 ),
    .Y(_8920_)
);

OAI22X1 _19620_ (
    .A(_8920_),
    .B(_8919_),
    .C(\datapath.idinstr_21_bF$buf16 ),
    .D(_8918_),
    .Y(_8921_)
);

OAI21X1 _19621_ (
    .A(_7420__bF$buf9),
    .B(_8921_),
    .C(_7423__bF$buf2),
    .Y(_8922_)
);

OAI22X1 _19622_ (
    .A(_7423__bF$buf1),
    .B(_8911_),
    .C(_8917_),
    .D(_8922_),
    .Y(_8923_)
);

NAND2X1 _19623_ (
    .A(_7451__bF$buf0),
    .B(_8923_),
    .Y(_8924_)
);

AOI22X1 _19624_ (
    .A(_7418__bF$buf0),
    .B(_7422__bF$buf0),
    .C(_8901_),
    .D(_8924_),
    .Y(\datapath.registers.regb_data [29])
);

NAND2X1 _19625_ (
    .A(\datapath.registers.838[27] [30]),
    .B(\datapath.idinstr_20_bF$buf0 ),
    .Y(_8925_)
);

NAND2X1 _19626_ (
    .A(\datapath.registers.838[26] [30]),
    .B(_7425__bF$buf19),
    .Y(_8926_)
);

NAND3X1 _19627_ (
    .A(\datapath.idinstr_21_bF$buf15 ),
    .B(_8925_),
    .C(_8926_),
    .Y(_8927_)
);

NAND2X1 _19628_ (
    .A(\datapath.registers.838[25] [30]),
    .B(\datapath.idinstr_20_bF$buf55 ),
    .Y(_8928_)
);

AOI21X1 _19629_ (
    .A(_7425__bF$buf18),
    .B(\datapath.registers.838[24] [30]),
    .C(\datapath.idinstr_21_bF$buf14 ),
    .Y(_8929_)
);

NAND2X1 _19630_ (
    .A(_8928_),
    .B(_8929_),
    .Y(_8930_)
);

NAND3X1 _19631_ (
    .A(_7420__bF$buf8),
    .B(_8927_),
    .C(_8930_),
    .Y(_8931_)
);

NAND2X1 _19632_ (
    .A(\datapath.registers.838[31] [30]),
    .B(\datapath.idinstr_20_bF$buf54 ),
    .Y(_8932_)
);

AOI21X1 _19633_ (
    .A(_7425__bF$buf17),
    .B(\datapath.registers.838[30] [30]),
    .C(_7419__bF$buf3),
    .Y(_8933_)
);

NAND2X1 _19634_ (
    .A(_8932_),
    .B(_8933_),
    .Y(_8934_)
);

AOI21X1 _19635_ (
    .A(\datapath.registers.838[29] [30]),
    .B(\datapath.idinstr_20_bF$buf53 ),
    .C(\datapath.idinstr_21_bF$buf13 ),
    .Y(_8935_)
);

OAI21X1 _19636_ (
    .A(_7326_),
    .B(\datapath.idinstr_20_bF$buf52 ),
    .C(_8935_),
    .Y(_8936_)
);

NAND3X1 _19637_ (
    .A(\datapath.idinstr_22_bF$buf29 ),
    .B(_8936_),
    .C(_8934_),
    .Y(_8937_)
);

AOI21X1 _19638_ (
    .A(_8931_),
    .B(_8937_),
    .C(_7423__bF$buf0),
    .Y(_8938_)
);

MUX2X1 _19639_ (
    .A(\datapath.registers.838[18] [30]),
    .B(\datapath.registers.838[16] [30]),
    .S(\datapath.idinstr_21_bF$buf12 ),
    .Y(_8939_)
);

NAND2X1 _19640_ (
    .A(_7425__bF$buf16),
    .B(_8939_),
    .Y(_8940_)
);

MUX2X1 _19641_ (
    .A(\datapath.registers.838[19] [30]),
    .B(\datapath.registers.838[17] [30]),
    .S(\datapath.idinstr_21_bF$buf11 ),
    .Y(_8941_)
);

NAND2X1 _19642_ (
    .A(\datapath.idinstr_20_bF$buf51 ),
    .B(_8941_),
    .Y(_8942_)
);

NAND3X1 _19643_ (
    .A(_7420__bF$buf7),
    .B(_8940_),
    .C(_8942_),
    .Y(_8943_)
);

MUX2X1 _19644_ (
    .A(\datapath.registers.838[22] [30]),
    .B(\datapath.registers.838[20] [30]),
    .S(\datapath.idinstr_21_bF$buf10 ),
    .Y(_8944_)
);

NAND2X1 _19645_ (
    .A(_7425__bF$buf15),
    .B(_8944_),
    .Y(_8945_)
);

MUX2X1 _19646_ (
    .A(\datapath.registers.838[23] [30]),
    .B(\datapath.registers.838[21] [30]),
    .S(\datapath.idinstr_21_bF$buf9 ),
    .Y(_8946_)
);

NAND2X1 _19647_ (
    .A(\datapath.idinstr_20_bF$buf50 ),
    .B(_8946_),
    .Y(_8947_)
);

NAND3X1 _19648_ (
    .A(\datapath.idinstr_22_bF$buf28 ),
    .B(_8945_),
    .C(_8947_),
    .Y(_8948_)
);

AOI21X1 _19649_ (
    .A(_8943_),
    .B(_8948_),
    .C(\datapath.idinstr_23_bF$buf6 ),
    .Y(_8949_)
);

OAI21X1 _19650_ (
    .A(_8949_),
    .B(_8938_),
    .C(\datapath.idinstr_24_bF$buf5 ),
    .Y(_8950_)
);

AOI21X1 _19651_ (
    .A(\datapath.registers.838[13] [30]),
    .B(\datapath.idinstr_22_bF$buf27 ),
    .C(_7425__bF$buf14),
    .Y(_8951_)
);

OAI21X1 _19652_ (
    .A(_5304_),
    .B(\datapath.idinstr_22_bF$buf26 ),
    .C(_8951_),
    .Y(_8952_)
);

INVX1 _19653_ (
    .A(\datapath.registers.838[8] [30]),
    .Y(_8953_)
);

AOI21X1 _19654_ (
    .A(\datapath.registers.838[12] [30]),
    .B(\datapath.idinstr_22_bF$buf25 ),
    .C(\datapath.idinstr_20_bF$buf49 ),
    .Y(_8954_)
);

OAI21X1 _19655_ (
    .A(_8953_),
    .B(\datapath.idinstr_22_bF$buf24 ),
    .C(_8954_),
    .Y(_8955_)
);

NAND3X1 _19656_ (
    .A(_7419__bF$buf2),
    .B(_8955_),
    .C(_8952_),
    .Y(_8956_)
);

INVX1 _19657_ (
    .A(\datapath.registers.838[11] [30]),
    .Y(_8957_)
);

AOI21X1 _19658_ (
    .A(\datapath.registers.838[15] [30]),
    .B(\datapath.idinstr_22_bF$buf23 ),
    .C(_7425__bF$buf13),
    .Y(_8958_)
);

OAI21X1 _19659_ (
    .A(_8957_),
    .B(\datapath.idinstr_22_bF$buf22 ),
    .C(_8958_),
    .Y(_8959_)
);

AOI21X1 _19660_ (
    .A(\datapath.registers.838[14] [30]),
    .B(\datapath.idinstr_22_bF$buf21 ),
    .C(\datapath.idinstr_20_bF$buf48 ),
    .Y(_8960_)
);

OAI21X1 _19661_ (
    .A(_5260_),
    .B(\datapath.idinstr_22_bF$buf20 ),
    .C(_8960_),
    .Y(_8961_)
);

NAND3X1 _19662_ (
    .A(\datapath.idinstr_21_bF$buf8 ),
    .B(_8961_),
    .C(_8959_),
    .Y(_8962_)
);

AOI21X1 _19663_ (
    .A(_8956_),
    .B(_8962_),
    .C(_7423__bF$buf7),
    .Y(_8963_)
);

MUX2X1 _19664_ (
    .A(\datapath.registers.838[1] [30]),
    .B(\datapath.registers.838[0] [30]),
    .S(\datapath.idinstr_20_bF$buf47 ),
    .Y(_8964_)
);

NOR2X1 _19665_ (
    .A(\datapath.registers.838[3] [30]),
    .B(_7425__bF$buf12),
    .Y(_8965_)
);

OAI21X1 _19666_ (
    .A(\datapath.registers.838[2] [30]),
    .B(\datapath.idinstr_20_bF$buf46 ),
    .C(\datapath.idinstr_21_bF$buf7 ),
    .Y(_8966_)
);

OAI22X1 _19667_ (
    .A(_8966_),
    .B(_8965_),
    .C(\datapath.idinstr_21_bF$buf6 ),
    .D(_8964_),
    .Y(_8967_)
);

NAND2X1 _19668_ (
    .A(_7420__bF$buf6),
    .B(_8967_),
    .Y(_8968_)
);

MUX2X1 _19669_ (
    .A(\datapath.registers.838[5] [30]),
    .B(\datapath.registers.838[4] [30]),
    .S(\datapath.idinstr_20_bF$buf45 ),
    .Y(_8969_)
);

NOR2X1 _19670_ (
    .A(\datapath.registers.838[7] [30]),
    .B(_7425__bF$buf11),
    .Y(_8970_)
);

OAI21X1 _19671_ (
    .A(\datapath.registers.838[6] [30]),
    .B(\datapath.idinstr_20_bF$buf44 ),
    .C(\datapath.idinstr_21_bF$buf5 ),
    .Y(_8971_)
);

OAI22X1 _19672_ (
    .A(_8971_),
    .B(_8970_),
    .C(\datapath.idinstr_21_bF$buf4 ),
    .D(_8969_),
    .Y(_8972_)
);

NAND2X1 _19673_ (
    .A(\datapath.idinstr_22_bF$buf19 ),
    .B(_8972_),
    .Y(_8973_)
);

AOI21X1 _19674_ (
    .A(_8968_),
    .B(_8973_),
    .C(\datapath.idinstr_23_bF$buf5 ),
    .Y(_8974_)
);

OAI21X1 _19675_ (
    .A(_8963_),
    .B(_8974_),
    .C(_7451__bF$buf4),
    .Y(_8975_)
);

AOI22X1 _19676_ (
    .A(_7418__bF$buf4),
    .B(_7422__bF$buf4),
    .C(_8950_),
    .D(_8975_),
    .Y(\datapath.registers.regb_data [30])
);

NAND2X1 _19677_ (
    .A(\datapath.registers.838[27] [31]),
    .B(\datapath.idinstr_20_bF$buf43 ),
    .Y(_8976_)
);

NAND2X1 _19678_ (
    .A(\datapath.registers.838[26] [31]),
    .B(_7425__bF$buf10),
    .Y(_8977_)
);

NAND3X1 _19679_ (
    .A(\datapath.idinstr_21_bF$buf3 ),
    .B(_8976_),
    .C(_8977_),
    .Y(_8978_)
);

NAND2X1 _19680_ (
    .A(\datapath.registers.838[25] [31]),
    .B(\datapath.idinstr_20_bF$buf42 ),
    .Y(_8979_)
);

AOI21X1 _19681_ (
    .A(_7425__bF$buf9),
    .B(\datapath.registers.838[24] [31]),
    .C(\datapath.idinstr_21_bF$buf2 ),
    .Y(_8980_)
);

NAND2X1 _19682_ (
    .A(_8979_),
    .B(_8980_),
    .Y(_8981_)
);

NAND3X1 _19683_ (
    .A(_7420__bF$buf5),
    .B(_8978_),
    .C(_8981_),
    .Y(_8982_)
);

NAND2X1 _19684_ (
    .A(\datapath.registers.838[31] [31]),
    .B(\datapath.idinstr_20_bF$buf41 ),
    .Y(_8983_)
);

AOI21X1 _19685_ (
    .A(_7425__bF$buf8),
    .B(\datapath.registers.838[30] [31]),
    .C(_7419__bF$buf1),
    .Y(_8984_)
);

NAND2X1 _19686_ (
    .A(_8983_),
    .B(_8984_),
    .Y(_8985_)
);

AOI21X1 _19687_ (
    .A(\datapath.registers.838[29] [31]),
    .B(\datapath.idinstr_20_bF$buf40 ),
    .C(\datapath.idinstr_21_bF$buf1 ),
    .Y(_8986_)
);

OAI21X1 _19688_ (
    .A(_7377_),
    .B(\datapath.idinstr_20_bF$buf39 ),
    .C(_8986_),
    .Y(_8987_)
);

NAND3X1 _19689_ (
    .A(\datapath.idinstr_22_bF$buf18 ),
    .B(_8987_),
    .C(_8985_),
    .Y(_8988_)
);

AOI21X1 _19690_ (
    .A(_8982_),
    .B(_8988_),
    .C(_7423__bF$buf6),
    .Y(_8989_)
);

MUX2X1 _19691_ (
    .A(\datapath.registers.838[18] [31]),
    .B(\datapath.registers.838[16] [31]),
    .S(\datapath.idinstr_21_bF$buf0 ),
    .Y(_8990_)
);

NAND2X1 _19692_ (
    .A(_7425__bF$buf7),
    .B(_8990_),
    .Y(_8991_)
);

MUX2X1 _19693_ (
    .A(\datapath.registers.838[19] [31]),
    .B(\datapath.registers.838[17] [31]),
    .S(\datapath.idinstr_21_bF$buf51 ),
    .Y(_8992_)
);

NAND2X1 _19694_ (
    .A(\datapath.idinstr_20_bF$buf38 ),
    .B(_8992_),
    .Y(_8993_)
);

NAND3X1 _19695_ (
    .A(_7420__bF$buf4),
    .B(_8991_),
    .C(_8993_),
    .Y(_8994_)
);

MUX2X1 _19696_ (
    .A(\datapath.registers.838[22] [31]),
    .B(\datapath.registers.838[20] [31]),
    .S(\datapath.idinstr_21_bF$buf50 ),
    .Y(_8995_)
);

NAND2X1 _19697_ (
    .A(_7425__bF$buf6),
    .B(_8995_),
    .Y(_8996_)
);

MUX2X1 _19698_ (
    .A(\datapath.registers.838[23] [31]),
    .B(\datapath.registers.838[21] [31]),
    .S(\datapath.idinstr_21_bF$buf49 ),
    .Y(_8997_)
);

NAND2X1 _19699_ (
    .A(\datapath.idinstr_20_bF$buf37 ),
    .B(_8997_),
    .Y(_8998_)
);

NAND3X1 _19700_ (
    .A(\datapath.idinstr_22_bF$buf17 ),
    .B(_8996_),
    .C(_8998_),
    .Y(_8999_)
);

AOI21X1 _19701_ (
    .A(_8994_),
    .B(_8999_),
    .C(\datapath.idinstr_23_bF$buf4 ),
    .Y(_9000_)
);

OAI21X1 _19702_ (
    .A(_9000_),
    .B(_8989_),
    .C(\datapath.idinstr_24_bF$buf4 ),
    .Y(_9001_)
);

MUX2X1 _19703_ (
    .A(\datapath.registers.838[9] [31]),
    .B(\datapath.registers.838[8] [31]),
    .S(\datapath.idinstr_20_bF$buf36 ),
    .Y(_9002_)
);

NOR2X1 _19704_ (
    .A(\datapath.registers.838[11] [31]),
    .B(_7425__bF$buf5),
    .Y(_9003_)
);

OAI21X1 _19705_ (
    .A(\datapath.registers.838[10] [31]),
    .B(\datapath.idinstr_20_bF$buf35 ),
    .C(\datapath.idinstr_21_bF$buf48 ),
    .Y(_9004_)
);

OAI22X1 _19706_ (
    .A(_9004_),
    .B(_9003_),
    .C(\datapath.idinstr_21_bF$buf47 ),
    .D(_9002_),
    .Y(_9005_)
);

AOI21X1 _19707_ (
    .A(_7425__bF$buf4),
    .B(\datapath.registers.838[14] [31]),
    .C(_7419__bF$buf0),
    .Y(_9006_)
);

OAI21X1 _19708_ (
    .A(_7398_),
    .B(_7425__bF$buf3),
    .C(_9006_),
    .Y(_9007_)
);

NAND2X1 _19709_ (
    .A(\datapath.registers.838[12] [31]),
    .B(_7425__bF$buf2),
    .Y(_9008_)
);

AOI21X1 _19710_ (
    .A(\datapath.registers.838[13] [31]),
    .B(\datapath.idinstr_20_bF$buf34 ),
    .C(\datapath.idinstr_21_bF$buf46 ),
    .Y(_9009_)
);

AOI21X1 _19711_ (
    .A(_9008_),
    .B(_9009_),
    .C(_7420__bF$buf3),
    .Y(_9010_)
);

AOI22X1 _19712_ (
    .A(_9007_),
    .B(_9010_),
    .C(_7420__bF$buf2),
    .D(_9005_),
    .Y(_9011_)
);

NOR2X1 _19713_ (
    .A(\datapath.registers.838[0] [31]),
    .B(\datapath.idinstr_20_bF$buf33 ),
    .Y(_9012_)
);

OAI21X1 _19714_ (
    .A(\datapath.registers.838[1] [31]),
    .B(_7425__bF$buf1),
    .C(_7419__bF$buf9),
    .Y(_9013_)
);

NOR2X1 _19715_ (
    .A(\datapath.registers.838[3] [31]),
    .B(_7425__bF$buf0),
    .Y(_9014_)
);

OAI21X1 _19716_ (
    .A(\datapath.registers.838[2] [31]),
    .B(\datapath.idinstr_20_bF$buf32 ),
    .C(\datapath.idinstr_21_bF$buf45 ),
    .Y(_9015_)
);

OAI22X1 _19717_ (
    .A(_9014_),
    .B(_9015_),
    .C(_9012_),
    .D(_9013_),
    .Y(_9016_)
);

NOR2X1 _19718_ (
    .A(\datapath.idinstr_22_bF$buf16 ),
    .B(_9016_),
    .Y(_9017_)
);

MUX2X1 _19719_ (
    .A(\datapath.registers.838[5] [31]),
    .B(\datapath.registers.838[4] [31]),
    .S(\datapath.idinstr_20_bF$buf31 ),
    .Y(_9018_)
);

NOR2X1 _19720_ (
    .A(\datapath.registers.838[7] [31]),
    .B(_7425__bF$buf47),
    .Y(_9019_)
);

OAI21X1 _19721_ (
    .A(\datapath.registers.838[6] [31]),
    .B(\datapath.idinstr_20_bF$buf30 ),
    .C(\datapath.idinstr_21_bF$buf44 ),
    .Y(_9020_)
);

OAI22X1 _19722_ (
    .A(_9020_),
    .B(_9019_),
    .C(\datapath.idinstr_21_bF$buf43 ),
    .D(_9018_),
    .Y(_9021_)
);

OAI21X1 _19723_ (
    .A(_7420__bF$buf1),
    .B(_9021_),
    .C(_7423__bF$buf5),
    .Y(_9022_)
);

OAI22X1 _19724_ (
    .A(_7423__bF$buf4),
    .B(_9011_),
    .C(_9017_),
    .D(_9022_),
    .Y(_9023_)
);

NAND2X1 _19725_ (
    .A(_7451__bF$buf3),
    .B(_9023_),
    .Y(_9024_)
);

AOI22X1 _19726_ (
    .A(_7418__bF$buf3),
    .B(_7422__bF$buf3),
    .C(_9001_),
    .D(_9024_),
    .Y(\datapath.registers.regb_data [31])
);

NAND2X1 _19727_ (
    .A(_5688_),
    .B(_5619_),
    .Y(_9025_)
);

OAI21X1 _19728_ (
    .A(_5687__bF$buf6),
    .B(_4968__bF$buf2),
    .C(\datapath.registers.838[29] [0]),
    .Y(_9026_)
);

OAI21X1 _19729_ (
    .A(_4786__bF$buf0),
    .B(_9025__bF$buf4),
    .C(_9026_),
    .Y(_4434_)
);

OAI21X1 _19730_ (
    .A(_5687__bF$buf5),
    .B(_4968__bF$buf1),
    .C(\datapath.registers.838[29] [1]),
    .Y(_9027_)
);

OAI21X1 _19731_ (
    .A(_4801__bF$buf3),
    .B(_9025__bF$buf3),
    .C(_9027_),
    .Y(_4445_)
);

OAI21X1 _19732_ (
    .A(_5687__bF$buf4),
    .B(_4968__bF$buf0),
    .C(\datapath.registers.838[29] [2]),
    .Y(_9028_)
);

OAI21X1 _19733_ (
    .A(_4803__bF$buf0),
    .B(_9025__bF$buf2),
    .C(_9028_),
    .Y(_4456_)
);

OAI21X1 _19734_ (
    .A(_5687__bF$buf3),
    .B(_4968__bF$buf9),
    .C(\datapath.registers.838[29] [3]),
    .Y(_9029_)
);

OAI21X1 _19735_ (
    .A(_4805__bF$buf1),
    .B(_9025__bF$buf1),
    .C(_9029_),
    .Y(_4459_)
);

OAI21X1 _19736_ (
    .A(_5687__bF$buf2),
    .B(_4968__bF$buf8),
    .C(\datapath.registers.838[29] [4]),
    .Y(_9030_)
);

OAI21X1 _19737_ (
    .A(_4807__bF$buf4),
    .B(_9025__bF$buf0),
    .C(_9030_),
    .Y(_4460_)
);

OAI21X1 _19738_ (
    .A(_5687__bF$buf1),
    .B(_4968__bF$buf7),
    .C(\datapath.registers.838[29] [5]),
    .Y(_9031_)
);

OAI21X1 _19739_ (
    .A(_4809__bF$buf4),
    .B(_9025__bF$buf4),
    .C(_9031_),
    .Y(_4461_)
);

OAI21X1 _19740_ (
    .A(_5687__bF$buf0),
    .B(_4968__bF$buf6),
    .C(\datapath.registers.838[29] [6]),
    .Y(_9032_)
);

OAI21X1 _19741_ (
    .A(_4811__bF$buf1),
    .B(_9025__bF$buf3),
    .C(_9032_),
    .Y(_4462_)
);

OAI21X1 _19742_ (
    .A(_5687__bF$buf8),
    .B(_4968__bF$buf5),
    .C(\datapath.registers.838[29] [7]),
    .Y(_9033_)
);

OAI21X1 _19743_ (
    .A(_4813__bF$buf3),
    .B(_9025__bF$buf2),
    .C(_9033_),
    .Y(_4463_)
);

OAI21X1 _19744_ (
    .A(_5687__bF$buf7),
    .B(_4968__bF$buf4),
    .C(\datapath.registers.838[29] [8]),
    .Y(_9034_)
);

OAI21X1 _19745_ (
    .A(_4815__bF$buf4),
    .B(_9025__bF$buf1),
    .C(_9034_),
    .Y(_4464_)
);

OAI21X1 _19746_ (
    .A(_5687__bF$buf6),
    .B(_4968__bF$buf3),
    .C(\datapath.registers.838[29] [9]),
    .Y(_9035_)
);

OAI21X1 _19747_ (
    .A(_4817__bF$buf2),
    .B(_9025__bF$buf0),
    .C(_9035_),
    .Y(_4465_)
);

OAI21X1 _19748_ (
    .A(_5687__bF$buf5),
    .B(_4968__bF$buf2),
    .C(\datapath.registers.838[29] [10]),
    .Y(_9036_)
);

OAI21X1 _19749_ (
    .A(_4819__bF$buf0),
    .B(_9025__bF$buf4),
    .C(_9036_),
    .Y(_4435_)
);

OAI21X1 _19750_ (
    .A(_5687__bF$buf4),
    .B(_4968__bF$buf1),
    .C(\datapath.registers.838[29] [11]),
    .Y(_9037_)
);

OAI21X1 _19751_ (
    .A(_4821__bF$buf3),
    .B(_9025__bF$buf3),
    .C(_9037_),
    .Y(_4436_)
);

OAI21X1 _19752_ (
    .A(_5687__bF$buf3),
    .B(_4968__bF$buf0),
    .C(\datapath.registers.838[29] [12]),
    .Y(_9038_)
);

OAI21X1 _19753_ (
    .A(_4823__bF$buf1),
    .B(_9025__bF$buf2),
    .C(_9038_),
    .Y(_4437_)
);

OAI21X1 _19754_ (
    .A(_5687__bF$buf2),
    .B(_4968__bF$buf9),
    .C(\datapath.registers.838[29] [13]),
    .Y(_9039_)
);

OAI21X1 _19755_ (
    .A(_4825__bF$buf3),
    .B(_9025__bF$buf1),
    .C(_9039_),
    .Y(_4438_)
);

OAI21X1 _19756_ (
    .A(_5687__bF$buf1),
    .B(_4968__bF$buf8),
    .C(\datapath.registers.838[29] [14]),
    .Y(_9040_)
);

OAI21X1 _19757_ (
    .A(_4827__bF$buf3),
    .B(_9025__bF$buf0),
    .C(_9040_),
    .Y(_4439_)
);

OAI21X1 _19758_ (
    .A(_5687__bF$buf0),
    .B(_4968__bF$buf7),
    .C(\datapath.registers.838[29] [15]),
    .Y(_9041_)
);

OAI21X1 _19759_ (
    .A(_4829__bF$buf3),
    .B(_9025__bF$buf4),
    .C(_9041_),
    .Y(_4440_)
);

OAI21X1 _19760_ (
    .A(_5687__bF$buf8),
    .B(_4968__bF$buf6),
    .C(\datapath.registers.838[29] [16]),
    .Y(_9042_)
);

OAI21X1 _19761_ (
    .A(_4831__bF$buf3),
    .B(_9025__bF$buf3),
    .C(_9042_),
    .Y(_4441_)
);

OAI21X1 _19762_ (
    .A(_5687__bF$buf7),
    .B(_4968__bF$buf5),
    .C(\datapath.registers.838[29] [17]),
    .Y(_9043_)
);

OAI21X1 _19763_ (
    .A(_4833__bF$buf0),
    .B(_9025__bF$buf2),
    .C(_9043_),
    .Y(_4442_)
);

OAI21X1 _19764_ (
    .A(_5687__bF$buf6),
    .B(_4968__bF$buf4),
    .C(\datapath.registers.838[29] [18]),
    .Y(_9044_)
);

OAI21X1 _19765_ (
    .A(_4835__bF$buf0),
    .B(_9025__bF$buf1),
    .C(_9044_),
    .Y(_4443_)
);

OAI21X1 _19766_ (
    .A(_5687__bF$buf5),
    .B(_4968__bF$buf3),
    .C(\datapath.registers.838[29] [19]),
    .Y(_9045_)
);

OAI21X1 _19767_ (
    .A(_4837__bF$buf1),
    .B(_9025__bF$buf0),
    .C(_9045_),
    .Y(_4444_)
);

OAI21X1 _19768_ (
    .A(_5687__bF$buf4),
    .B(_4968__bF$buf2),
    .C(\datapath.registers.838[29] [20]),
    .Y(_9046_)
);

OAI21X1 _19769_ (
    .A(_4839__bF$buf3),
    .B(_9025__bF$buf4),
    .C(_9046_),
    .Y(_4446_)
);

OAI21X1 _19770_ (
    .A(_5687__bF$buf3),
    .B(_4968__bF$buf1),
    .C(\datapath.registers.838[29] [21]),
    .Y(_9047_)
);

OAI21X1 _19771_ (
    .A(_4841__bF$buf0),
    .B(_9025__bF$buf3),
    .C(_9047_),
    .Y(_4447_)
);

OAI21X1 _19772_ (
    .A(_5687__bF$buf2),
    .B(_4968__bF$buf0),
    .C(\datapath.registers.838[29] [22]),
    .Y(_9048_)
);

OAI21X1 _19773_ (
    .A(_4843__bF$buf4),
    .B(_9025__bF$buf2),
    .C(_9048_),
    .Y(_4448_)
);

OAI21X1 _19774_ (
    .A(_5687__bF$buf1),
    .B(_4968__bF$buf9),
    .C(\datapath.registers.838[29] [23]),
    .Y(_9049_)
);

OAI21X1 _19775_ (
    .A(_4845__bF$buf0),
    .B(_9025__bF$buf1),
    .C(_9049_),
    .Y(_4449_)
);

OAI21X1 _19776_ (
    .A(_5687__bF$buf0),
    .B(_4968__bF$buf8),
    .C(\datapath.registers.838[29] [24]),
    .Y(_9050_)
);

OAI21X1 _19777_ (
    .A(_4847__bF$buf2),
    .B(_9025__bF$buf0),
    .C(_9050_),
    .Y(_4450_)
);

OAI21X1 _19778_ (
    .A(_5687__bF$buf8),
    .B(_4968__bF$buf7),
    .C(\datapath.registers.838[29] [25]),
    .Y(_9051_)
);

OAI21X1 _19779_ (
    .A(_4849__bF$buf0),
    .B(_9025__bF$buf4),
    .C(_9051_),
    .Y(_4451_)
);

OAI21X1 _19780_ (
    .A(_5687__bF$buf7),
    .B(_4968__bF$buf6),
    .C(\datapath.registers.838[29] [26]),
    .Y(_9052_)
);

OAI21X1 _19781_ (
    .A(_4851__bF$buf3),
    .B(_9025__bF$buf3),
    .C(_9052_),
    .Y(_4452_)
);

OAI21X1 _19782_ (
    .A(_5687__bF$buf6),
    .B(_4968__bF$buf5),
    .C(\datapath.registers.838[29] [27]),
    .Y(_9053_)
);

OAI21X1 _19783_ (
    .A(_4853__bF$buf4),
    .B(_9025__bF$buf2),
    .C(_9053_),
    .Y(_4453_)
);

OAI21X1 _19784_ (
    .A(_5687__bF$buf5),
    .B(_4968__bF$buf4),
    .C(\datapath.registers.838[29] [28]),
    .Y(_9054_)
);

OAI21X1 _19785_ (
    .A(_4855__bF$buf3),
    .B(_9025__bF$buf1),
    .C(_9054_),
    .Y(_4454_)
);

OAI21X1 _19786_ (
    .A(_5687__bF$buf4),
    .B(_4968__bF$buf3),
    .C(\datapath.registers.838[29] [29]),
    .Y(_9055_)
);

OAI21X1 _19787_ (
    .A(_4857__bF$buf3),
    .B(_9025__bF$buf0),
    .C(_9055_),
    .Y(_4455_)
);

OAI21X1 _19788_ (
    .A(_5687__bF$buf3),
    .B(_4968__bF$buf2),
    .C(\datapath.registers.838[29] [30]),
    .Y(_9056_)
);

OAI21X1 _19789_ (
    .A(_4859__bF$buf0),
    .B(_9025__bF$buf4),
    .C(_9056_),
    .Y(_4457_)
);

OAI21X1 _19790_ (
    .A(_5687__bF$buf2),
    .B(_4968__bF$buf1),
    .C(\datapath.registers.838[29] [31]),
    .Y(_9057_)
);

OAI21X1 _19791_ (
    .A(_4861__bF$buf3),
    .B(_9025__bF$buf3),
    .C(_9057_),
    .Y(_4458_)
);

NAND3X1 _19792_ (
    .A(_4789_),
    .B(_5688_),
    .C(_5015_),
    .Y(_9058_)
);

NAND2X1 _19793_ (
    .A(\datapath.registers.838[28] [0]),
    .B(_9058__bF$buf7),
    .Y(_9059_)
);

OAI21X1 _19794_ (
    .A(_4786__bF$buf4),
    .B(_9058__bF$buf6),
    .C(_9059_),
    .Y(_4402_)
);

NAND2X1 _19795_ (
    .A(\datapath.registers.838[28] [1]),
    .B(_9058__bF$buf5),
    .Y(_9060_)
);

OAI21X1 _19796_ (
    .A(_4801__bF$buf2),
    .B(_9058__bF$buf4),
    .C(_9060_),
    .Y(_4413_)
);

NAND2X1 _19797_ (
    .A(\datapath.registers.838[28] [2]),
    .B(_9058__bF$buf3),
    .Y(_9061_)
);

OAI21X1 _19798_ (
    .A(_4803__bF$buf4),
    .B(_9058__bF$buf2),
    .C(_9061_),
    .Y(_4424_)
);

NAND2X1 _19799_ (
    .A(\datapath.registers.838[28] [3]),
    .B(_9058__bF$buf1),
    .Y(_9062_)
);

OAI21X1 _19800_ (
    .A(_4805__bF$buf0),
    .B(_9058__bF$buf0),
    .C(_9062_),
    .Y(_4427_)
);

NAND2X1 _19801_ (
    .A(\datapath.registers.838[28] [4]),
    .B(_9058__bF$buf7),
    .Y(_9063_)
);

OAI21X1 _19802_ (
    .A(_4807__bF$buf3),
    .B(_9058__bF$buf6),
    .C(_9063_),
    .Y(_4428_)
);

NAND2X1 _19803_ (
    .A(\datapath.registers.838[28] [5]),
    .B(_9058__bF$buf5),
    .Y(_9064_)
);

OAI21X1 _19804_ (
    .A(_4809__bF$buf3),
    .B(_9058__bF$buf4),
    .C(_9064_),
    .Y(_4429_)
);

NAND2X1 _19805_ (
    .A(\datapath.registers.838[28] [6]),
    .B(_9058__bF$buf3),
    .Y(_9065_)
);

OAI21X1 _19806_ (
    .A(_4811__bF$buf0),
    .B(_9058__bF$buf2),
    .C(_9065_),
    .Y(_4430_)
);

NAND2X1 _19807_ (
    .A(\datapath.registers.838[28] [7]),
    .B(_9058__bF$buf1),
    .Y(_9066_)
);

OAI21X1 _19808_ (
    .A(_4813__bF$buf2),
    .B(_9058__bF$buf0),
    .C(_9066_),
    .Y(_4431_)
);

NAND2X1 _19809_ (
    .A(\datapath.registers.838[28] [8]),
    .B(_9058__bF$buf7),
    .Y(_9067_)
);

OAI21X1 _19810_ (
    .A(_4815__bF$buf3),
    .B(_9058__bF$buf6),
    .C(_9067_),
    .Y(_4432_)
);

NAND2X1 _19811_ (
    .A(\datapath.registers.838[28] [9]),
    .B(_9058__bF$buf5),
    .Y(_9068_)
);

OAI21X1 _19812_ (
    .A(_4817__bF$buf1),
    .B(_9058__bF$buf4),
    .C(_9068_),
    .Y(_4433_)
);

NAND2X1 _19813_ (
    .A(\datapath.registers.838[28] [10]),
    .B(_9058__bF$buf3),
    .Y(_9069_)
);

OAI21X1 _19814_ (
    .A(_4819__bF$buf4),
    .B(_9058__bF$buf2),
    .C(_9069_),
    .Y(_4403_)
);

NAND2X1 _19815_ (
    .A(\datapath.registers.838[28] [11]),
    .B(_9058__bF$buf1),
    .Y(_9070_)
);

OAI21X1 _19816_ (
    .A(_4821__bF$buf2),
    .B(_9058__bF$buf0),
    .C(_9070_),
    .Y(_4404_)
);

NAND2X1 _19817_ (
    .A(\datapath.registers.838[28] [12]),
    .B(_9058__bF$buf7),
    .Y(_9071_)
);

OAI21X1 _19818_ (
    .A(_4823__bF$buf0),
    .B(_9058__bF$buf6),
    .C(_9071_),
    .Y(_4405_)
);

NAND2X1 _19819_ (
    .A(\datapath.registers.838[28] [13]),
    .B(_9058__bF$buf5),
    .Y(_9072_)
);

OAI21X1 _19820_ (
    .A(_4825__bF$buf2),
    .B(_9058__bF$buf4),
    .C(_9072_),
    .Y(_4406_)
);

NAND2X1 _19821_ (
    .A(\datapath.registers.838[28] [14]),
    .B(_9058__bF$buf3),
    .Y(_9073_)
);

OAI21X1 _19822_ (
    .A(_4827__bF$buf2),
    .B(_9058__bF$buf2),
    .C(_9073_),
    .Y(_4407_)
);

NAND2X1 _19823_ (
    .A(\datapath.registers.838[28] [15]),
    .B(_9058__bF$buf1),
    .Y(_9074_)
);

OAI21X1 _19824_ (
    .A(_4829__bF$buf2),
    .B(_9058__bF$buf0),
    .C(_9074_),
    .Y(_4408_)
);

NAND2X1 _19825_ (
    .A(\datapath.registers.838[28] [16]),
    .B(_9058__bF$buf7),
    .Y(_9075_)
);

OAI21X1 _19826_ (
    .A(_4831__bF$buf2),
    .B(_9058__bF$buf6),
    .C(_9075_),
    .Y(_4409_)
);

NAND2X1 _19827_ (
    .A(\datapath.registers.838[28] [17]),
    .B(_9058__bF$buf5),
    .Y(_9076_)
);

OAI21X1 _19828_ (
    .A(_4833__bF$buf4),
    .B(_9058__bF$buf4),
    .C(_9076_),
    .Y(_4410_)
);

NAND2X1 _19829_ (
    .A(\datapath.registers.838[28] [18]),
    .B(_9058__bF$buf3),
    .Y(_9077_)
);

OAI21X1 _19830_ (
    .A(_4835__bF$buf4),
    .B(_9058__bF$buf2),
    .C(_9077_),
    .Y(_4411_)
);

NAND2X1 _19831_ (
    .A(\datapath.registers.838[28] [19]),
    .B(_9058__bF$buf1),
    .Y(_9078_)
);

OAI21X1 _19832_ (
    .A(_4837__bF$buf0),
    .B(_9058__bF$buf0),
    .C(_9078_),
    .Y(_4412_)
);

NAND2X1 _19833_ (
    .A(\datapath.registers.838[28] [20]),
    .B(_9058__bF$buf7),
    .Y(_9079_)
);

OAI21X1 _19834_ (
    .A(_4839__bF$buf2),
    .B(_9058__bF$buf6),
    .C(_9079_),
    .Y(_4414_)
);

NAND2X1 _19835_ (
    .A(\datapath.registers.838[28] [21]),
    .B(_9058__bF$buf5),
    .Y(_9080_)
);

OAI21X1 _19836_ (
    .A(_4841__bF$buf4),
    .B(_9058__bF$buf4),
    .C(_9080_),
    .Y(_4415_)
);

NAND2X1 _19837_ (
    .A(\datapath.registers.838[28] [22]),
    .B(_9058__bF$buf3),
    .Y(_9081_)
);

OAI21X1 _19838_ (
    .A(_4843__bF$buf3),
    .B(_9058__bF$buf2),
    .C(_9081_),
    .Y(_4416_)
);

NAND2X1 _19839_ (
    .A(\datapath.registers.838[28] [23]),
    .B(_9058__bF$buf1),
    .Y(_9082_)
);

OAI21X1 _19840_ (
    .A(_4845__bF$buf4),
    .B(_9058__bF$buf0),
    .C(_9082_),
    .Y(_4417_)
);

NAND2X1 _19841_ (
    .A(\datapath.registers.838[28] [24]),
    .B(_9058__bF$buf7),
    .Y(_9083_)
);

OAI21X1 _19842_ (
    .A(_4847__bF$buf1),
    .B(_9058__bF$buf6),
    .C(_9083_),
    .Y(_4418_)
);

NAND2X1 _19843_ (
    .A(\datapath.registers.838[28] [25]),
    .B(_9058__bF$buf5),
    .Y(_9084_)
);

OAI21X1 _19844_ (
    .A(_4849__bF$buf4),
    .B(_9058__bF$buf4),
    .C(_9084_),
    .Y(_4419_)
);

NAND2X1 _19845_ (
    .A(\datapath.registers.838[28] [26]),
    .B(_9058__bF$buf3),
    .Y(_9085_)
);

OAI21X1 _19846_ (
    .A(_4851__bF$buf2),
    .B(_9058__bF$buf2),
    .C(_9085_),
    .Y(_4420_)
);

NAND2X1 _19847_ (
    .A(\datapath.registers.838[28] [27]),
    .B(_9058__bF$buf1),
    .Y(_9086_)
);

OAI21X1 _19848_ (
    .A(_4853__bF$buf3),
    .B(_9058__bF$buf0),
    .C(_9086_),
    .Y(_4421_)
);

NAND2X1 _19849_ (
    .A(\datapath.registers.838[28] [28]),
    .B(_9058__bF$buf7),
    .Y(_9087_)
);

OAI21X1 _19850_ (
    .A(_4855__bF$buf2),
    .B(_9058__bF$buf6),
    .C(_9087_),
    .Y(_4422_)
);

NAND2X1 _19851_ (
    .A(\datapath.registers.838[28] [29]),
    .B(_9058__bF$buf5),
    .Y(_9088_)
);

OAI21X1 _19852_ (
    .A(_4857__bF$buf2),
    .B(_9058__bF$buf4),
    .C(_9088_),
    .Y(_4423_)
);

NAND2X1 _19853_ (
    .A(\datapath.registers.838[28] [30]),
    .B(_9058__bF$buf3),
    .Y(_9089_)
);

OAI21X1 _19854_ (
    .A(_4859__bF$buf4),
    .B(_9058__bF$buf2),
    .C(_9089_),
    .Y(_4425_)
);

NAND2X1 _19855_ (
    .A(\datapath.registers.838[28] [31]),
    .B(_9058__bF$buf1),
    .Y(_9090_)
);

OAI21X1 _19856_ (
    .A(_4861__bF$buf2),
    .B(_9058__bF$buf0),
    .C(_9090_),
    .Y(_4426_)
);

NAND2X1 _19857_ (
    .A(_5476_),
    .B(_5686_),
    .Y(_9091_)
);

INVX8 _19858_ (
    .A(_5476_),
    .Y(_9092_)
);

OAI21X1 _19859_ (
    .A(_9092__bF$buf8),
    .B(_4899__bF$buf1),
    .C(\datapath.registers.838[27] [0]),
    .Y(_9093_)
);

OAI21X1 _19860_ (
    .A(_4786__bF$buf3),
    .B(_9091__bF$buf4),
    .C(_9093_),
    .Y(_4370_)
);

OAI21X1 _19861_ (
    .A(_9092__bF$buf7),
    .B(_4899__bF$buf0),
    .C(\datapath.registers.838[27] [1]),
    .Y(_9094_)
);

OAI21X1 _19862_ (
    .A(_4801__bF$buf1),
    .B(_9091__bF$buf3),
    .C(_9094_),
    .Y(_4381_)
);

OAI21X1 _19863_ (
    .A(_9092__bF$buf6),
    .B(_4899__bF$buf13),
    .C(\datapath.registers.838[27] [2]),
    .Y(_9095_)
);

OAI21X1 _19864_ (
    .A(_4803__bF$buf3),
    .B(_9091__bF$buf2),
    .C(_9095_),
    .Y(_4392_)
);

OAI21X1 _19865_ (
    .A(_9092__bF$buf5),
    .B(_4899__bF$buf12),
    .C(\datapath.registers.838[27] [3]),
    .Y(_9096_)
);

OAI21X1 _19866_ (
    .A(_4805__bF$buf4),
    .B(_9091__bF$buf1),
    .C(_9096_),
    .Y(_4395_)
);

OAI21X1 _19867_ (
    .A(_9092__bF$buf4),
    .B(_4899__bF$buf11),
    .C(\datapath.registers.838[27] [4]),
    .Y(_9097_)
);

OAI21X1 _19868_ (
    .A(_4807__bF$buf2),
    .B(_9091__bF$buf0),
    .C(_9097_),
    .Y(_4396_)
);

OAI21X1 _19869_ (
    .A(_9092__bF$buf3),
    .B(_4899__bF$buf10),
    .C(\datapath.registers.838[27] [5]),
    .Y(_9098_)
);

OAI21X1 _19870_ (
    .A(_4809__bF$buf2),
    .B(_9091__bF$buf4),
    .C(_9098_),
    .Y(_4397_)
);

OAI21X1 _19871_ (
    .A(_9092__bF$buf2),
    .B(_4899__bF$buf9),
    .C(\datapath.registers.838[27] [6]),
    .Y(_9099_)
);

OAI21X1 _19872_ (
    .A(_4811__bF$buf4),
    .B(_9091__bF$buf3),
    .C(_9099_),
    .Y(_4398_)
);

OAI21X1 _19873_ (
    .A(_9092__bF$buf1),
    .B(_4899__bF$buf8),
    .C(\datapath.registers.838[27] [7]),
    .Y(_9100_)
);

OAI21X1 _19874_ (
    .A(_4813__bF$buf1),
    .B(_9091__bF$buf2),
    .C(_9100_),
    .Y(_4399_)
);

OAI21X1 _19875_ (
    .A(_9092__bF$buf0),
    .B(_4899__bF$buf7),
    .C(\datapath.registers.838[27] [8]),
    .Y(_9101_)
);

OAI21X1 _19876_ (
    .A(_4815__bF$buf2),
    .B(_9091__bF$buf1),
    .C(_9101_),
    .Y(_4400_)
);

OAI21X1 _19877_ (
    .A(_9092__bF$buf8),
    .B(_4899__bF$buf6),
    .C(\datapath.registers.838[27] [9]),
    .Y(_9102_)
);

OAI21X1 _19878_ (
    .A(_4817__bF$buf0),
    .B(_9091__bF$buf0),
    .C(_9102_),
    .Y(_4401_)
);

OAI21X1 _19879_ (
    .A(_9092__bF$buf7),
    .B(_4899__bF$buf5),
    .C(\datapath.registers.838[27] [10]),
    .Y(_9103_)
);

OAI21X1 _19880_ (
    .A(_4819__bF$buf3),
    .B(_9091__bF$buf4),
    .C(_9103_),
    .Y(_4371_)
);

OAI21X1 _19881_ (
    .A(_9092__bF$buf6),
    .B(_4899__bF$buf4),
    .C(\datapath.registers.838[27] [11]),
    .Y(_9104_)
);

OAI21X1 _19882_ (
    .A(_4821__bF$buf1),
    .B(_9091__bF$buf3),
    .C(_9104_),
    .Y(_4372_)
);

OAI21X1 _19883_ (
    .A(_9092__bF$buf5),
    .B(_4899__bF$buf3),
    .C(\datapath.registers.838[27] [12]),
    .Y(_9105_)
);

OAI21X1 _19884_ (
    .A(_4823__bF$buf4),
    .B(_9091__bF$buf2),
    .C(_9105_),
    .Y(_4373_)
);

OAI21X1 _19885_ (
    .A(_9092__bF$buf4),
    .B(_4899__bF$buf2),
    .C(\datapath.registers.838[27] [13]),
    .Y(_9106_)
);

OAI21X1 _19886_ (
    .A(_4825__bF$buf1),
    .B(_9091__bF$buf1),
    .C(_9106_),
    .Y(_4374_)
);

OAI21X1 _19887_ (
    .A(_9092__bF$buf3),
    .B(_4899__bF$buf1),
    .C(\datapath.registers.838[27] [14]),
    .Y(_9107_)
);

OAI21X1 _19888_ (
    .A(_4827__bF$buf1),
    .B(_9091__bF$buf0),
    .C(_9107_),
    .Y(_4375_)
);

OAI21X1 _19889_ (
    .A(_9092__bF$buf2),
    .B(_4899__bF$buf0),
    .C(\datapath.registers.838[27] [15]),
    .Y(_9108_)
);

OAI21X1 _19890_ (
    .A(_4829__bF$buf1),
    .B(_9091__bF$buf4),
    .C(_9108_),
    .Y(_4376_)
);

OAI21X1 _19891_ (
    .A(_9092__bF$buf1),
    .B(_4899__bF$buf13),
    .C(\datapath.registers.838[27] [16]),
    .Y(_9109_)
);

OAI21X1 _19892_ (
    .A(_4831__bF$buf1),
    .B(_9091__bF$buf3),
    .C(_9109_),
    .Y(_4377_)
);

OAI21X1 _19893_ (
    .A(_9092__bF$buf0),
    .B(_4899__bF$buf12),
    .C(\datapath.registers.838[27] [17]),
    .Y(_9110_)
);

OAI21X1 _19894_ (
    .A(_4833__bF$buf3),
    .B(_9091__bF$buf2),
    .C(_9110_),
    .Y(_4378_)
);

OAI21X1 _19895_ (
    .A(_9092__bF$buf8),
    .B(_4899__bF$buf11),
    .C(\datapath.registers.838[27] [18]),
    .Y(_9111_)
);

OAI21X1 _19896_ (
    .A(_4835__bF$buf3),
    .B(_9091__bF$buf1),
    .C(_9111_),
    .Y(_4379_)
);

OAI21X1 _19897_ (
    .A(_9092__bF$buf7),
    .B(_4899__bF$buf10),
    .C(\datapath.registers.838[27] [19]),
    .Y(_9112_)
);

OAI21X1 _19898_ (
    .A(_4837__bF$buf4),
    .B(_9091__bF$buf0),
    .C(_9112_),
    .Y(_4380_)
);

OAI21X1 _19899_ (
    .A(_9092__bF$buf6),
    .B(_4899__bF$buf9),
    .C(\datapath.registers.838[27] [20]),
    .Y(_9113_)
);

OAI21X1 _19900_ (
    .A(_4839__bF$buf1),
    .B(_9091__bF$buf4),
    .C(_9113_),
    .Y(_4382_)
);

OAI21X1 _19901_ (
    .A(_9092__bF$buf5),
    .B(_4899__bF$buf8),
    .C(\datapath.registers.838[27] [21]),
    .Y(_9114_)
);

OAI21X1 _19902_ (
    .A(_4841__bF$buf3),
    .B(_9091__bF$buf3),
    .C(_9114_),
    .Y(_4383_)
);

OAI21X1 _19903_ (
    .A(_9092__bF$buf4),
    .B(_4899__bF$buf7),
    .C(\datapath.registers.838[27] [22]),
    .Y(_9115_)
);

OAI21X1 _19904_ (
    .A(_4843__bF$buf2),
    .B(_9091__bF$buf2),
    .C(_9115_),
    .Y(_4384_)
);

OAI21X1 _19905_ (
    .A(_9092__bF$buf3),
    .B(_4899__bF$buf6),
    .C(\datapath.registers.838[27] [23]),
    .Y(_9116_)
);

OAI21X1 _19906_ (
    .A(_4845__bF$buf3),
    .B(_9091__bF$buf1),
    .C(_9116_),
    .Y(_4385_)
);

OAI21X1 _19907_ (
    .A(_9092__bF$buf2),
    .B(_4899__bF$buf5),
    .C(\datapath.registers.838[27] [24]),
    .Y(_9117_)
);

OAI21X1 _19908_ (
    .A(_4847__bF$buf0),
    .B(_9091__bF$buf0),
    .C(_9117_),
    .Y(_4386_)
);

OAI21X1 _19909_ (
    .A(_9092__bF$buf1),
    .B(_4899__bF$buf4),
    .C(\datapath.registers.838[27] [25]),
    .Y(_9118_)
);

OAI21X1 _19910_ (
    .A(_4849__bF$buf3),
    .B(_9091__bF$buf4),
    .C(_9118_),
    .Y(_4387_)
);

OAI21X1 _19911_ (
    .A(_9092__bF$buf0),
    .B(_4899__bF$buf3),
    .C(\datapath.registers.838[27] [26]),
    .Y(_9119_)
);

OAI21X1 _19912_ (
    .A(_4851__bF$buf1),
    .B(_9091__bF$buf3),
    .C(_9119_),
    .Y(_4388_)
);

OAI21X1 _19913_ (
    .A(_9092__bF$buf8),
    .B(_4899__bF$buf2),
    .C(\datapath.registers.838[27] [27]),
    .Y(_9120_)
);

OAI21X1 _19914_ (
    .A(_4853__bF$buf2),
    .B(_9091__bF$buf2),
    .C(_9120_),
    .Y(_4389_)
);

OAI21X1 _19915_ (
    .A(_9092__bF$buf7),
    .B(_4899__bF$buf1),
    .C(\datapath.registers.838[27] [28]),
    .Y(_9121_)
);

OAI21X1 _19916_ (
    .A(_4855__bF$buf1),
    .B(_9091__bF$buf1),
    .C(_9121_),
    .Y(_4390_)
);

OAI21X1 _19917_ (
    .A(_9092__bF$buf6),
    .B(_4899__bF$buf0),
    .C(\datapath.registers.838[27] [29]),
    .Y(_9122_)
);

OAI21X1 _19918_ (
    .A(_4857__bF$buf1),
    .B(_9091__bF$buf0),
    .C(_9122_),
    .Y(_4391_)
);

OAI21X1 _19919_ (
    .A(_9092__bF$buf5),
    .B(_4899__bF$buf13),
    .C(\datapath.registers.838[27] [30]),
    .Y(_9123_)
);

OAI21X1 _19920_ (
    .A(_4859__bF$buf3),
    .B(_9091__bF$buf4),
    .C(_9123_),
    .Y(_4393_)
);

OAI21X1 _19921_ (
    .A(_9092__bF$buf4),
    .B(_4899__bF$buf12),
    .C(\datapath.registers.838[27] [31]),
    .Y(_9124_)
);

OAI21X1 _19922_ (
    .A(_4861__bF$buf1),
    .B(_9091__bF$buf3),
    .C(_9124_),
    .Y(_4394_)
);

NAND2X1 _19923_ (
    .A(_5476_),
    .B(_5585_),
    .Y(_9125_)
);

OAI21X1 _19924_ (
    .A(_4934__bF$buf0),
    .B(_9092__bF$buf3),
    .C(\datapath.registers.838[26] [0]),
    .Y(_9126_)
);

OAI21X1 _19925_ (
    .A(_4786__bF$buf2),
    .B(_9125__bF$buf4),
    .C(_9126_),
    .Y(_4338_)
);

OAI21X1 _19926_ (
    .A(_4934__bF$buf9),
    .B(_9092__bF$buf2),
    .C(\datapath.registers.838[26] [1]),
    .Y(_9127_)
);

OAI21X1 _19927_ (
    .A(_4801__bF$buf0),
    .B(_9125__bF$buf3),
    .C(_9127_),
    .Y(_4349_)
);

OAI21X1 _19928_ (
    .A(_4934__bF$buf8),
    .B(_9092__bF$buf1),
    .C(\datapath.registers.838[26] [2]),
    .Y(_9128_)
);

OAI21X1 _19929_ (
    .A(_4803__bF$buf2),
    .B(_9125__bF$buf2),
    .C(_9128_),
    .Y(_4360_)
);

OAI21X1 _19930_ (
    .A(_4934__bF$buf7),
    .B(_9092__bF$buf0),
    .C(\datapath.registers.838[26] [3]),
    .Y(_9129_)
);

OAI21X1 _19931_ (
    .A(_4805__bF$buf3),
    .B(_9125__bF$buf1),
    .C(_9129_),
    .Y(_4363_)
);

OAI21X1 _19932_ (
    .A(_4934__bF$buf6),
    .B(_9092__bF$buf8),
    .C(\datapath.registers.838[26] [4]),
    .Y(_9130_)
);

OAI21X1 _19933_ (
    .A(_4807__bF$buf1),
    .B(_9125__bF$buf0),
    .C(_9130_),
    .Y(_4364_)
);

OAI21X1 _19934_ (
    .A(_4934__bF$buf5),
    .B(_9092__bF$buf7),
    .C(\datapath.registers.838[26] [5]),
    .Y(_9131_)
);

OAI21X1 _19935_ (
    .A(_4809__bF$buf1),
    .B(_9125__bF$buf4),
    .C(_9131_),
    .Y(_4365_)
);

OAI21X1 _19936_ (
    .A(_4934__bF$buf4),
    .B(_9092__bF$buf6),
    .C(\datapath.registers.838[26] [6]),
    .Y(_9132_)
);

OAI21X1 _19937_ (
    .A(_4811__bF$buf3),
    .B(_9125__bF$buf3),
    .C(_9132_),
    .Y(_4366_)
);

OAI21X1 _19938_ (
    .A(_4934__bF$buf3),
    .B(_9092__bF$buf5),
    .C(\datapath.registers.838[26] [7]),
    .Y(_9133_)
);

OAI21X1 _19939_ (
    .A(_4813__bF$buf0),
    .B(_9125__bF$buf2),
    .C(_9133_),
    .Y(_4367_)
);

OAI21X1 _19940_ (
    .A(_4934__bF$buf2),
    .B(_9092__bF$buf4),
    .C(\datapath.registers.838[26] [8]),
    .Y(_9134_)
);

OAI21X1 _19941_ (
    .A(_4815__bF$buf1),
    .B(_9125__bF$buf1),
    .C(_9134_),
    .Y(_4368_)
);

OAI21X1 _19942_ (
    .A(_4934__bF$buf1),
    .B(_9092__bF$buf3),
    .C(\datapath.registers.838[26] [9]),
    .Y(_9135_)
);

OAI21X1 _19943_ (
    .A(_4817__bF$buf4),
    .B(_9125__bF$buf0),
    .C(_9135_),
    .Y(_4369_)
);

OAI21X1 _19944_ (
    .A(_4934__bF$buf0),
    .B(_9092__bF$buf2),
    .C(\datapath.registers.838[26] [10]),
    .Y(_9136_)
);

OAI21X1 _19945_ (
    .A(_4819__bF$buf2),
    .B(_9125__bF$buf4),
    .C(_9136_),
    .Y(_4339_)
);

OAI21X1 _19946_ (
    .A(_4934__bF$buf9),
    .B(_9092__bF$buf1),
    .C(\datapath.registers.838[26] [11]),
    .Y(_9137_)
);

OAI21X1 _19947_ (
    .A(_4821__bF$buf0),
    .B(_9125__bF$buf3),
    .C(_9137_),
    .Y(_4340_)
);

OAI21X1 _19948_ (
    .A(_4934__bF$buf8),
    .B(_9092__bF$buf0),
    .C(\datapath.registers.838[26] [12]),
    .Y(_9138_)
);

OAI21X1 _19949_ (
    .A(_4823__bF$buf3),
    .B(_9125__bF$buf2),
    .C(_9138_),
    .Y(_4341_)
);

OAI21X1 _19950_ (
    .A(_4934__bF$buf7),
    .B(_9092__bF$buf8),
    .C(\datapath.registers.838[26] [13]),
    .Y(_9139_)
);

OAI21X1 _19951_ (
    .A(_4825__bF$buf0),
    .B(_9125__bF$buf1),
    .C(_9139_),
    .Y(_4342_)
);

OAI21X1 _19952_ (
    .A(_4934__bF$buf6),
    .B(_9092__bF$buf7),
    .C(\datapath.registers.838[26] [14]),
    .Y(_9140_)
);

OAI21X1 _19953_ (
    .A(_4827__bF$buf0),
    .B(_9125__bF$buf0),
    .C(_9140_),
    .Y(_4343_)
);

OAI21X1 _19954_ (
    .A(_4934__bF$buf5),
    .B(_9092__bF$buf6),
    .C(\datapath.registers.838[26] [15]),
    .Y(_9141_)
);

OAI21X1 _19955_ (
    .A(_4829__bF$buf0),
    .B(_9125__bF$buf4),
    .C(_9141_),
    .Y(_4344_)
);

OAI21X1 _19956_ (
    .A(_4934__bF$buf4),
    .B(_9092__bF$buf5),
    .C(\datapath.registers.838[26] [16]),
    .Y(_9142_)
);

OAI21X1 _19957_ (
    .A(_4831__bF$buf0),
    .B(_9125__bF$buf3),
    .C(_9142_),
    .Y(_4345_)
);

OAI21X1 _19958_ (
    .A(_4934__bF$buf3),
    .B(_9092__bF$buf4),
    .C(\datapath.registers.838[26] [17]),
    .Y(_9143_)
);

OAI21X1 _19959_ (
    .A(_4833__bF$buf2),
    .B(_9125__bF$buf2),
    .C(_9143_),
    .Y(_4346_)
);

OAI21X1 _19960_ (
    .A(_4934__bF$buf2),
    .B(_9092__bF$buf3),
    .C(\datapath.registers.838[26] [18]),
    .Y(_9144_)
);

OAI21X1 _19961_ (
    .A(_4835__bF$buf2),
    .B(_9125__bF$buf1),
    .C(_9144_),
    .Y(_4347_)
);

OAI21X1 _19962_ (
    .A(_4934__bF$buf1),
    .B(_9092__bF$buf2),
    .C(\datapath.registers.838[26] [19]),
    .Y(_9145_)
);

OAI21X1 _19963_ (
    .A(_4837__bF$buf3),
    .B(_9125__bF$buf0),
    .C(_9145_),
    .Y(_4348_)
);

OAI21X1 _19964_ (
    .A(_4934__bF$buf0),
    .B(_9092__bF$buf1),
    .C(\datapath.registers.838[26] [20]),
    .Y(_9146_)
);

OAI21X1 _19965_ (
    .A(_4839__bF$buf0),
    .B(_9125__bF$buf4),
    .C(_9146_),
    .Y(_4350_)
);

OAI21X1 _19966_ (
    .A(_4934__bF$buf9),
    .B(_9092__bF$buf0),
    .C(\datapath.registers.838[26] [21]),
    .Y(_9147_)
);

OAI21X1 _19967_ (
    .A(_4841__bF$buf2),
    .B(_9125__bF$buf3),
    .C(_9147_),
    .Y(_4351_)
);

OAI21X1 _19968_ (
    .A(_4934__bF$buf8),
    .B(_9092__bF$buf8),
    .C(\datapath.registers.838[26] [22]),
    .Y(_9148_)
);

OAI21X1 _19969_ (
    .A(_4843__bF$buf1),
    .B(_9125__bF$buf2),
    .C(_9148_),
    .Y(_4352_)
);

OAI21X1 _19970_ (
    .A(_4934__bF$buf7),
    .B(_9092__bF$buf7),
    .C(\datapath.registers.838[26] [23]),
    .Y(_9149_)
);

OAI21X1 _19971_ (
    .A(_4845__bF$buf2),
    .B(_9125__bF$buf1),
    .C(_9149_),
    .Y(_4353_)
);

OAI21X1 _19972_ (
    .A(_4934__bF$buf6),
    .B(_9092__bF$buf6),
    .C(\datapath.registers.838[26] [24]),
    .Y(_9150_)
);

OAI21X1 _19973_ (
    .A(_4847__bF$buf4),
    .B(_9125__bF$buf0),
    .C(_9150_),
    .Y(_4354_)
);

OAI21X1 _19974_ (
    .A(_4934__bF$buf5),
    .B(_9092__bF$buf5),
    .C(\datapath.registers.838[26] [25]),
    .Y(_9151_)
);

OAI21X1 _19975_ (
    .A(_4849__bF$buf2),
    .B(_9125__bF$buf4),
    .C(_9151_),
    .Y(_4355_)
);

OAI21X1 _19976_ (
    .A(_4934__bF$buf4),
    .B(_9092__bF$buf4),
    .C(\datapath.registers.838[26] [26]),
    .Y(_9152_)
);

OAI21X1 _19977_ (
    .A(_4851__bF$buf0),
    .B(_9125__bF$buf3),
    .C(_9152_),
    .Y(_4356_)
);

OAI21X1 _19978_ (
    .A(_4934__bF$buf3),
    .B(_9092__bF$buf3),
    .C(\datapath.registers.838[26] [27]),
    .Y(_9153_)
);

OAI21X1 _19979_ (
    .A(_4853__bF$buf1),
    .B(_9125__bF$buf2),
    .C(_9153_),
    .Y(_4357_)
);

OAI21X1 _19980_ (
    .A(_4934__bF$buf2),
    .B(_9092__bF$buf2),
    .C(\datapath.registers.838[26] [28]),
    .Y(_9154_)
);

OAI21X1 _19981_ (
    .A(_4855__bF$buf0),
    .B(_9125__bF$buf1),
    .C(_9154_),
    .Y(_4358_)
);

OAI21X1 _19982_ (
    .A(_4934__bF$buf1),
    .B(_9092__bF$buf1),
    .C(\datapath.registers.838[26] [29]),
    .Y(_9155_)
);

OAI21X1 _19983_ (
    .A(_4857__bF$buf0),
    .B(_9125__bF$buf0),
    .C(_9155_),
    .Y(_4359_)
);

OAI21X1 _19984_ (
    .A(_4934__bF$buf0),
    .B(_9092__bF$buf0),
    .C(\datapath.registers.838[26] [30]),
    .Y(_9156_)
);

OAI21X1 _19985_ (
    .A(_4859__bF$buf2),
    .B(_9125__bF$buf4),
    .C(_9156_),
    .Y(_4361_)
);

OAI21X1 _19986_ (
    .A(_4934__bF$buf9),
    .B(_9092__bF$buf8),
    .C(\datapath.registers.838[26] [31]),
    .Y(_9157_)
);

OAI21X1 _19987_ (
    .A(_4861__bF$buf0),
    .B(_9125__bF$buf3),
    .C(_9157_),
    .Y(_4362_)
);

NAND2X1 _19988_ (
    .A(_5476_),
    .B(_5619_),
    .Y(_9158_)
);

OAI21X1 _19989_ (
    .A(_4968__bF$buf0),
    .B(_9092__bF$buf7),
    .C(\datapath.registers.838[25] [0]),
    .Y(_9159_)
);

OAI21X1 _19990_ (
    .A(_4786__bF$buf1),
    .B(_9158__bF$buf4),
    .C(_9159_),
    .Y(_4306_)
);

OAI21X1 _19991_ (
    .A(_4968__bF$buf9),
    .B(_9092__bF$buf6),
    .C(\datapath.registers.838[25] [1]),
    .Y(_9160_)
);

OAI21X1 _19992_ (
    .A(_4801__bF$buf4),
    .B(_9158__bF$buf3),
    .C(_9160_),
    .Y(_4317_)
);

OAI21X1 _19993_ (
    .A(_4968__bF$buf8),
    .B(_9092__bF$buf5),
    .C(\datapath.registers.838[25] [2]),
    .Y(_9161_)
);

OAI21X1 _19994_ (
    .A(_4803__bF$buf1),
    .B(_9158__bF$buf2),
    .C(_9161_),
    .Y(_4328_)
);

OAI21X1 _19995_ (
    .A(_4968__bF$buf7),
    .B(_9092__bF$buf4),
    .C(\datapath.registers.838[25] [3]),
    .Y(_9162_)
);

OAI21X1 _19996_ (
    .A(_4805__bF$buf2),
    .B(_9158__bF$buf1),
    .C(_9162_),
    .Y(_4331_)
);

OAI21X1 _19997_ (
    .A(_4968__bF$buf6),
    .B(_9092__bF$buf3),
    .C(\datapath.registers.838[25] [4]),
    .Y(_9163_)
);

OAI21X1 _19998_ (
    .A(_4807__bF$buf0),
    .B(_9158__bF$buf0),
    .C(_9163_),
    .Y(_4332_)
);

OAI21X1 _19999_ (
    .A(_4968__bF$buf5),
    .B(_9092__bF$buf2),
    .C(\datapath.registers.838[25] [5]),
    .Y(_9164_)
);

OAI21X1 _20000_ (
    .A(_4809__bF$buf0),
    .B(_9158__bF$buf4),
    .C(_9164_),
    .Y(_4333_)
);

OAI21X1 _20001_ (
    .A(_4968__bF$buf4),
    .B(_9092__bF$buf1),
    .C(\datapath.registers.838[25] [6]),
    .Y(_9165_)
);

OAI21X1 _20002_ (
    .A(_4811__bF$buf2),
    .B(_9158__bF$buf3),
    .C(_9165_),
    .Y(_4334_)
);

OAI21X1 _20003_ (
    .A(_4968__bF$buf3),
    .B(_9092__bF$buf0),
    .C(\datapath.registers.838[25] [7]),
    .Y(_9166_)
);

OAI21X1 _20004_ (
    .A(_4813__bF$buf4),
    .B(_9158__bF$buf2),
    .C(_9166_),
    .Y(_4335_)
);

OAI21X1 _20005_ (
    .A(_4968__bF$buf2),
    .B(_9092__bF$buf8),
    .C(\datapath.registers.838[25] [8]),
    .Y(_9167_)
);

OAI21X1 _20006_ (
    .A(_4815__bF$buf0),
    .B(_9158__bF$buf1),
    .C(_9167_),
    .Y(_4336_)
);

OAI21X1 _20007_ (
    .A(_4968__bF$buf1),
    .B(_9092__bF$buf7),
    .C(\datapath.registers.838[25] [9]),
    .Y(_9168_)
);

OAI21X1 _20008_ (
    .A(_4817__bF$buf3),
    .B(_9158__bF$buf0),
    .C(_9168_),
    .Y(_4337_)
);

OAI21X1 _20009_ (
    .A(_4968__bF$buf0),
    .B(_9092__bF$buf6),
    .C(\datapath.registers.838[25] [10]),
    .Y(_9169_)
);

OAI21X1 _20010_ (
    .A(_4819__bF$buf1),
    .B(_9158__bF$buf4),
    .C(_9169_),
    .Y(_4307_)
);

OAI21X1 _20011_ (
    .A(_4968__bF$buf9),
    .B(_9092__bF$buf5),
    .C(\datapath.registers.838[25] [11]),
    .Y(_9170_)
);

OAI21X1 _20012_ (
    .A(_4821__bF$buf4),
    .B(_9158__bF$buf3),
    .C(_9170_),
    .Y(_4308_)
);

OAI21X1 _20013_ (
    .A(_4968__bF$buf8),
    .B(_9092__bF$buf4),
    .C(\datapath.registers.838[25] [12]),
    .Y(_9171_)
);

OAI21X1 _20014_ (
    .A(_4823__bF$buf2),
    .B(_9158__bF$buf2),
    .C(_9171_),
    .Y(_4309_)
);

OAI21X1 _20015_ (
    .A(_4968__bF$buf7),
    .B(_9092__bF$buf3),
    .C(\datapath.registers.838[25] [13]),
    .Y(_9172_)
);

OAI21X1 _20016_ (
    .A(_4825__bF$buf4),
    .B(_9158__bF$buf1),
    .C(_9172_),
    .Y(_4310_)
);

OAI21X1 _20017_ (
    .A(_4968__bF$buf6),
    .B(_9092__bF$buf2),
    .C(\datapath.registers.838[25] [14]),
    .Y(_9173_)
);

OAI21X1 _20018_ (
    .A(_4827__bF$buf4),
    .B(_9158__bF$buf0),
    .C(_9173_),
    .Y(_4311_)
);

OAI21X1 _20019_ (
    .A(_4968__bF$buf5),
    .B(_9092__bF$buf1),
    .C(\datapath.registers.838[25] [15]),
    .Y(_9174_)
);

OAI21X1 _20020_ (
    .A(_4829__bF$buf4),
    .B(_9158__bF$buf4),
    .C(_9174_),
    .Y(_4312_)
);

OAI21X1 _20021_ (
    .A(_4968__bF$buf4),
    .B(_9092__bF$buf0),
    .C(\datapath.registers.838[25] [16]),
    .Y(_9175_)
);

OAI21X1 _20022_ (
    .A(_4831__bF$buf4),
    .B(_9158__bF$buf3),
    .C(_9175_),
    .Y(_4313_)
);

OAI21X1 _20023_ (
    .A(_4968__bF$buf3),
    .B(_9092__bF$buf8),
    .C(\datapath.registers.838[25] [17]),
    .Y(_9176_)
);

OAI21X1 _20024_ (
    .A(_4833__bF$buf1),
    .B(_9158__bF$buf2),
    .C(_9176_),
    .Y(_4314_)
);

OAI21X1 _20025_ (
    .A(_4968__bF$buf2),
    .B(_9092__bF$buf7),
    .C(\datapath.registers.838[25] [18]),
    .Y(_9177_)
);

OAI21X1 _20026_ (
    .A(_4835__bF$buf1),
    .B(_9158__bF$buf1),
    .C(_9177_),
    .Y(_4315_)
);

OAI21X1 _20027_ (
    .A(_4968__bF$buf1),
    .B(_9092__bF$buf6),
    .C(\datapath.registers.838[25] [19]),
    .Y(_9178_)
);

OAI21X1 _20028_ (
    .A(_4837__bF$buf2),
    .B(_9158__bF$buf0),
    .C(_9178_),
    .Y(_4316_)
);

OAI21X1 _20029_ (
    .A(_4968__bF$buf0),
    .B(_9092__bF$buf5),
    .C(\datapath.registers.838[25] [20]),
    .Y(_9179_)
);

OAI21X1 _20030_ (
    .A(_4839__bF$buf4),
    .B(_9158__bF$buf4),
    .C(_9179_),
    .Y(_4318_)
);

OAI21X1 _20031_ (
    .A(_4968__bF$buf9),
    .B(_9092__bF$buf4),
    .C(\datapath.registers.838[25] [21]),
    .Y(_9180_)
);

OAI21X1 _20032_ (
    .A(_4841__bF$buf1),
    .B(_9158__bF$buf3),
    .C(_9180_),
    .Y(_4319_)
);

OAI21X1 _20033_ (
    .A(_4968__bF$buf8),
    .B(_9092__bF$buf3),
    .C(\datapath.registers.838[25] [22]),
    .Y(_9181_)
);

OAI21X1 _20034_ (
    .A(_4843__bF$buf0),
    .B(_9158__bF$buf2),
    .C(_9181_),
    .Y(_4320_)
);

OAI21X1 _20035_ (
    .A(_4968__bF$buf7),
    .B(_9092__bF$buf2),
    .C(\datapath.registers.838[25] [23]),
    .Y(_9182_)
);

OAI21X1 _20036_ (
    .A(_4845__bF$buf1),
    .B(_9158__bF$buf1),
    .C(_9182_),
    .Y(_4321_)
);

OAI21X1 _20037_ (
    .A(_4968__bF$buf6),
    .B(_9092__bF$buf1),
    .C(\datapath.registers.838[25] [24]),
    .Y(_9183_)
);

OAI21X1 _20038_ (
    .A(_4847__bF$buf3),
    .B(_9158__bF$buf0),
    .C(_9183_),
    .Y(_4322_)
);

OAI21X1 _20039_ (
    .A(_4968__bF$buf5),
    .B(_9092__bF$buf0),
    .C(\datapath.registers.838[25] [25]),
    .Y(_9184_)
);

OAI21X1 _20040_ (
    .A(_4849__bF$buf1),
    .B(_9158__bF$buf4),
    .C(_9184_),
    .Y(_4323_)
);

OAI21X1 _20041_ (
    .A(_4968__bF$buf4),
    .B(_9092__bF$buf8),
    .C(\datapath.registers.838[25] [26]),
    .Y(_9185_)
);

OAI21X1 _20042_ (
    .A(_4851__bF$buf4),
    .B(_9158__bF$buf3),
    .C(_9185_),
    .Y(_4324_)
);

OAI21X1 _20043_ (
    .A(_4968__bF$buf3),
    .B(_9092__bF$buf7),
    .C(\datapath.registers.838[25] [27]),
    .Y(_9186_)
);

OAI21X1 _20044_ (
    .A(_4853__bF$buf0),
    .B(_9158__bF$buf2),
    .C(_9186_),
    .Y(_4325_)
);

OAI21X1 _20045_ (
    .A(_4968__bF$buf2),
    .B(_9092__bF$buf6),
    .C(\datapath.registers.838[25] [28]),
    .Y(_9187_)
);

OAI21X1 _20046_ (
    .A(_4855__bF$buf4),
    .B(_9158__bF$buf1),
    .C(_9187_),
    .Y(_4326_)
);

OAI21X1 _20047_ (
    .A(_4968__bF$buf1),
    .B(_9092__bF$buf5),
    .C(\datapath.registers.838[25] [29]),
    .Y(_9188_)
);

OAI21X1 _20048_ (
    .A(_4857__bF$buf4),
    .B(_9158__bF$buf0),
    .C(_9188_),
    .Y(_4327_)
);

OAI21X1 _20049_ (
    .A(_4968__bF$buf0),
    .B(_9092__bF$buf4),
    .C(\datapath.registers.838[25] [30]),
    .Y(_9189_)
);

OAI21X1 _20050_ (
    .A(_4859__bF$buf1),
    .B(_9158__bF$buf4),
    .C(_9189_),
    .Y(_4329_)
);

OAI21X1 _20051_ (
    .A(_4968__bF$buf9),
    .B(_9092__bF$buf3),
    .C(\datapath.registers.838[25] [31]),
    .Y(_9190_)
);

OAI21X1 _20052_ (
    .A(_4861__bF$buf4),
    .B(_9158__bF$buf3),
    .C(_9190_),
    .Y(_4330_)
);

BUFX2 _20053_ (
    .A(\datapath.registers.838[0] [0]),
    .Y(_3762_)
);

BUFX2 _20054_ (
    .A(\datapath.registers.838[0] [1]),
    .Y(_3773_)
);

BUFX2 _20055_ (
    .A(\datapath.registers.838[0] [2]),
    .Y(_3784_)
);

BUFX2 _20056_ (
    .A(\datapath.registers.838[0] [3]),
    .Y(_3787_)
);

BUFX2 _20057_ (
    .A(\datapath.registers.838[0] [4]),
    .Y(_3788_)
);

BUFX2 _20058_ (
    .A(\datapath.registers.838[0] [5]),
    .Y(_3789_)
);

BUFX2 _20059_ (
    .A(\datapath.registers.838[0] [6]),
    .Y(_3790_)
);

BUFX2 _20060_ (
    .A(\datapath.registers.838[0] [7]),
    .Y(_3791_)
);

BUFX2 _20061_ (
    .A(\datapath.registers.838[0] [8]),
    .Y(_3792_)
);

BUFX2 _20062_ (
    .A(\datapath.registers.838[0] [9]),
    .Y(_3793_)
);

BUFX2 _20063_ (
    .A(\datapath.registers.838[0] [10]),
    .Y(_3763_)
);

BUFX2 _20064_ (
    .A(\datapath.registers.838[0] [11]),
    .Y(_3764_)
);

BUFX2 _20065_ (
    .A(\datapath.registers.838[0] [12]),
    .Y(_3765_)
);

BUFX2 _20066_ (
    .A(\datapath.registers.838[0] [13]),
    .Y(_3766_)
);

BUFX2 _20067_ (
    .A(\datapath.registers.838[0] [14]),
    .Y(_3767_)
);

BUFX2 _20068_ (
    .A(\datapath.registers.838[0] [15]),
    .Y(_3768_)
);

BUFX2 _20069_ (
    .A(\datapath.registers.838[0] [16]),
    .Y(_3769_)
);

BUFX2 _20070_ (
    .A(\datapath.registers.838[0] [17]),
    .Y(_3770_)
);

BUFX2 _20071_ (
    .A(\datapath.registers.838[0] [18]),
    .Y(_3771_)
);

BUFX2 _20072_ (
    .A(\datapath.registers.838[0] [19]),
    .Y(_3772_)
);

BUFX2 _20073_ (
    .A(\datapath.registers.838[0] [20]),
    .Y(_3774_)
);

BUFX2 _20074_ (
    .A(\datapath.registers.838[0] [21]),
    .Y(_3775_)
);

BUFX2 _20075_ (
    .A(\datapath.registers.838[0] [22]),
    .Y(_3776_)
);

BUFX2 _20076_ (
    .A(\datapath.registers.838[0] [23]),
    .Y(_3777_)
);

BUFX2 _20077_ (
    .A(\datapath.registers.838[0] [24]),
    .Y(_3778_)
);

BUFX2 _20078_ (
    .A(\datapath.registers.838[0] [25]),
    .Y(_3779_)
);

BUFX2 _20079_ (
    .A(\datapath.registers.838[0] [26]),
    .Y(_3780_)
);

BUFX2 _20080_ (
    .A(\datapath.registers.838[0] [27]),
    .Y(_3781_)
);

BUFX2 _20081_ (
    .A(\datapath.registers.838[0] [28]),
    .Y(_3782_)
);

BUFX2 _20082_ (
    .A(\datapath.registers.838[0] [29]),
    .Y(_3783_)
);

BUFX2 _20083_ (
    .A(\datapath.registers.838[0] [30]),
    .Y(_3785_)
);

BUFX2 _20084_ (
    .A(\datapath.registers.838[0] [31]),
    .Y(_3786_)
);

DFFPOSX1 _20085_ (
    .CLK(CLK_bF$buf47),
    .D(_4370_),
    .Q(\datapath.registers.838[27] [0])
);

DFFPOSX1 _20086_ (
    .CLK(CLK_bF$buf46),
    .D(_4381_),
    .Q(\datapath.registers.838[27] [1])
);

DFFPOSX1 _20087_ (
    .CLK(CLK_bF$buf45),
    .D(_4392_),
    .Q(\datapath.registers.838[27] [2])
);

DFFPOSX1 _20088_ (
    .CLK(CLK_bF$buf44),
    .D(_4395_),
    .Q(\datapath.registers.838[27] [3])
);

DFFPOSX1 _20089_ (
    .CLK(CLK_bF$buf43),
    .D(_4396_),
    .Q(\datapath.registers.838[27] [4])
);

DFFPOSX1 _20090_ (
    .CLK(CLK_bF$buf42),
    .D(_4397_),
    .Q(\datapath.registers.838[27] [5])
);

DFFPOSX1 _20091_ (
    .CLK(CLK_bF$buf41),
    .D(_4398_),
    .Q(\datapath.registers.838[27] [6])
);

DFFPOSX1 _20092_ (
    .CLK(CLK_bF$buf40),
    .D(_4399_),
    .Q(\datapath.registers.838[27] [7])
);

DFFPOSX1 _20093_ (
    .CLK(CLK_bF$buf39),
    .D(_4400_),
    .Q(\datapath.registers.838[27] [8])
);

DFFPOSX1 _20094_ (
    .CLK(CLK_bF$buf38),
    .D(_4401_),
    .Q(\datapath.registers.838[27] [9])
);

DFFPOSX1 _20095_ (
    .CLK(CLK_bF$buf37),
    .D(_4371_),
    .Q(\datapath.registers.838[27] [10])
);

DFFPOSX1 _20096_ (
    .CLK(CLK_bF$buf36),
    .D(_4372_),
    .Q(\datapath.registers.838[27] [11])
);

DFFPOSX1 _20097_ (
    .CLK(CLK_bF$buf35),
    .D(_4373_),
    .Q(\datapath.registers.838[27] [12])
);

DFFPOSX1 _20098_ (
    .CLK(CLK_bF$buf34),
    .D(_4374_),
    .Q(\datapath.registers.838[27] [13])
);

DFFPOSX1 _20099_ (
    .CLK(CLK_bF$buf33),
    .D(_4375_),
    .Q(\datapath.registers.838[27] [14])
);

DFFPOSX1 _20100_ (
    .CLK(CLK_bF$buf32),
    .D(_4376_),
    .Q(\datapath.registers.838[27] [15])
);

DFFPOSX1 _20101_ (
    .CLK(CLK_bF$buf31),
    .D(_4377_),
    .Q(\datapath.registers.838[27] [16])
);

DFFPOSX1 _20102_ (
    .CLK(CLK_bF$buf30),
    .D(_4378_),
    .Q(\datapath.registers.838[27] [17])
);

DFFPOSX1 _20103_ (
    .CLK(CLK_bF$buf29),
    .D(_4379_),
    .Q(\datapath.registers.838[27] [18])
);

DFFPOSX1 _20104_ (
    .CLK(CLK_bF$buf28),
    .D(_4380_),
    .Q(\datapath.registers.838[27] [19])
);

DFFPOSX1 _20105_ (
    .CLK(CLK_bF$buf27),
    .D(_4382_),
    .Q(\datapath.registers.838[27] [20])
);

DFFPOSX1 _20106_ (
    .CLK(CLK_bF$buf26),
    .D(_4383_),
    .Q(\datapath.registers.838[27] [21])
);

DFFPOSX1 _20107_ (
    .CLK(CLK_bF$buf25),
    .D(_4384_),
    .Q(\datapath.registers.838[27] [22])
);

DFFPOSX1 _20108_ (
    .CLK(CLK_bF$buf24),
    .D(_4385_),
    .Q(\datapath.registers.838[27] [23])
);

DFFPOSX1 _20109_ (
    .CLK(CLK_bF$buf23),
    .D(_4386_),
    .Q(\datapath.registers.838[27] [24])
);

DFFPOSX1 _20110_ (
    .CLK(CLK_bF$buf22),
    .D(_4387_),
    .Q(\datapath.registers.838[27] [25])
);

DFFPOSX1 _20111_ (
    .CLK(CLK_bF$buf21),
    .D(_4388_),
    .Q(\datapath.registers.838[27] [26])
);

DFFPOSX1 _20112_ (
    .CLK(CLK_bF$buf20),
    .D(_4389_),
    .Q(\datapath.registers.838[27] [27])
);

DFFPOSX1 _20113_ (
    .CLK(CLK_bF$buf19),
    .D(_4390_),
    .Q(\datapath.registers.838[27] [28])
);

DFFPOSX1 _20114_ (
    .CLK(CLK_bF$buf18),
    .D(_4391_),
    .Q(\datapath.registers.838[27] [29])
);

DFFPOSX1 _20115_ (
    .CLK(CLK_bF$buf17),
    .D(_4393_),
    .Q(\datapath.registers.838[27] [30])
);

DFFPOSX1 _20116_ (
    .CLK(CLK_bF$buf16),
    .D(_4394_),
    .Q(\datapath.registers.838[27] [31])
);

DFFPOSX1 _20117_ (
    .CLK(CLK_bF$buf15),
    .D(_4338_),
    .Q(\datapath.registers.838[26] [0])
);

DFFPOSX1 _20118_ (
    .CLK(CLK_bF$buf14),
    .D(_4349_),
    .Q(\datapath.registers.838[26] [1])
);

DFFPOSX1 _20119_ (
    .CLK(CLK_bF$buf13),
    .D(_4360_),
    .Q(\datapath.registers.838[26] [2])
);

DFFPOSX1 _20120_ (
    .CLK(CLK_bF$buf12),
    .D(_4363_),
    .Q(\datapath.registers.838[26] [3])
);

DFFPOSX1 _20121_ (
    .CLK(CLK_bF$buf11),
    .D(_4364_),
    .Q(\datapath.registers.838[26] [4])
);

DFFPOSX1 _20122_ (
    .CLK(CLK_bF$buf10),
    .D(_4365_),
    .Q(\datapath.registers.838[26] [5])
);

DFFPOSX1 _20123_ (
    .CLK(CLK_bF$buf9),
    .D(_4366_),
    .Q(\datapath.registers.838[26] [6])
);

DFFPOSX1 _20124_ (
    .CLK(CLK_bF$buf8),
    .D(_4367_),
    .Q(\datapath.registers.838[26] [7])
);

DFFPOSX1 _20125_ (
    .CLK(CLK_bF$buf7),
    .D(_4368_),
    .Q(\datapath.registers.838[26] [8])
);

DFFPOSX1 _20126_ (
    .CLK(CLK_bF$buf6),
    .D(_4369_),
    .Q(\datapath.registers.838[26] [9])
);

DFFPOSX1 _20127_ (
    .CLK(CLK_bF$buf5),
    .D(_4339_),
    .Q(\datapath.registers.838[26] [10])
);

DFFPOSX1 _20128_ (
    .CLK(CLK_bF$buf4),
    .D(_4340_),
    .Q(\datapath.registers.838[26] [11])
);

DFFPOSX1 _20129_ (
    .CLK(CLK_bF$buf3),
    .D(_4341_),
    .Q(\datapath.registers.838[26] [12])
);

DFFPOSX1 _20130_ (
    .CLK(CLK_bF$buf2),
    .D(_4342_),
    .Q(\datapath.registers.838[26] [13])
);

DFFPOSX1 _20131_ (
    .CLK(CLK_bF$buf1),
    .D(_4343_),
    .Q(\datapath.registers.838[26] [14])
);

DFFPOSX1 _20132_ (
    .CLK(CLK_bF$buf0),
    .D(_4344_),
    .Q(\datapath.registers.838[26] [15])
);

DFFPOSX1 _20133_ (
    .CLK(CLK_bF$buf151),
    .D(_4345_),
    .Q(\datapath.registers.838[26] [16])
);

DFFPOSX1 _20134_ (
    .CLK(CLK_bF$buf150),
    .D(_4346_),
    .Q(\datapath.registers.838[26] [17])
);

DFFPOSX1 _20135_ (
    .CLK(CLK_bF$buf149),
    .D(_4347_),
    .Q(\datapath.registers.838[26] [18])
);

DFFPOSX1 _20136_ (
    .CLK(CLK_bF$buf148),
    .D(_4348_),
    .Q(\datapath.registers.838[26] [19])
);

DFFPOSX1 _20137_ (
    .CLK(CLK_bF$buf147),
    .D(_4350_),
    .Q(\datapath.registers.838[26] [20])
);

DFFPOSX1 _20138_ (
    .CLK(CLK_bF$buf146),
    .D(_4351_),
    .Q(\datapath.registers.838[26] [21])
);

DFFPOSX1 _20139_ (
    .CLK(CLK_bF$buf145),
    .D(_4352_),
    .Q(\datapath.registers.838[26] [22])
);

DFFPOSX1 _20140_ (
    .CLK(CLK_bF$buf144),
    .D(_4353_),
    .Q(\datapath.registers.838[26] [23])
);

DFFPOSX1 _20141_ (
    .CLK(CLK_bF$buf143),
    .D(_4354_),
    .Q(\datapath.registers.838[26] [24])
);

DFFPOSX1 _20142_ (
    .CLK(CLK_bF$buf142),
    .D(_4355_),
    .Q(\datapath.registers.838[26] [25])
);

DFFPOSX1 _20143_ (
    .CLK(CLK_bF$buf141),
    .D(_4356_),
    .Q(\datapath.registers.838[26] [26])
);

DFFPOSX1 _20144_ (
    .CLK(CLK_bF$buf140),
    .D(_4357_),
    .Q(\datapath.registers.838[26] [27])
);

DFFPOSX1 _20145_ (
    .CLK(CLK_bF$buf139),
    .D(_4358_),
    .Q(\datapath.registers.838[26] [28])
);

DFFPOSX1 _20146_ (
    .CLK(CLK_bF$buf138),
    .D(_4359_),
    .Q(\datapath.registers.838[26] [29])
);

DFFPOSX1 _20147_ (
    .CLK(CLK_bF$buf137),
    .D(_4361_),
    .Q(\datapath.registers.838[26] [30])
);

DFFPOSX1 _20148_ (
    .CLK(CLK_bF$buf136),
    .D(_4362_),
    .Q(\datapath.registers.838[26] [31])
);

DFFPOSX1 _20149_ (
    .CLK(CLK_bF$buf135),
    .D(_4306_),
    .Q(\datapath.registers.838[25] [0])
);

DFFPOSX1 _20150_ (
    .CLK(CLK_bF$buf134),
    .D(_4317_),
    .Q(\datapath.registers.838[25] [1])
);

DFFPOSX1 _20151_ (
    .CLK(CLK_bF$buf133),
    .D(_4328_),
    .Q(\datapath.registers.838[25] [2])
);

DFFPOSX1 _20152_ (
    .CLK(CLK_bF$buf132),
    .D(_4331_),
    .Q(\datapath.registers.838[25] [3])
);

DFFPOSX1 _20153_ (
    .CLK(CLK_bF$buf131),
    .D(_4332_),
    .Q(\datapath.registers.838[25] [4])
);

DFFPOSX1 _20154_ (
    .CLK(CLK_bF$buf130),
    .D(_4333_),
    .Q(\datapath.registers.838[25] [5])
);

DFFPOSX1 _20155_ (
    .CLK(CLK_bF$buf129),
    .D(_4334_),
    .Q(\datapath.registers.838[25] [6])
);

DFFPOSX1 _20156_ (
    .CLK(CLK_bF$buf128),
    .D(_4335_),
    .Q(\datapath.registers.838[25] [7])
);

DFFPOSX1 _20157_ (
    .CLK(CLK_bF$buf127),
    .D(_4336_),
    .Q(\datapath.registers.838[25] [8])
);

DFFPOSX1 _20158_ (
    .CLK(CLK_bF$buf126),
    .D(_4337_),
    .Q(\datapath.registers.838[25] [9])
);

DFFPOSX1 _20159_ (
    .CLK(CLK_bF$buf125),
    .D(_4307_),
    .Q(\datapath.registers.838[25] [10])
);

DFFPOSX1 _20160_ (
    .CLK(CLK_bF$buf124),
    .D(_4308_),
    .Q(\datapath.registers.838[25] [11])
);

DFFPOSX1 _20161_ (
    .CLK(CLK_bF$buf123),
    .D(_4309_),
    .Q(\datapath.registers.838[25] [12])
);

DFFPOSX1 _20162_ (
    .CLK(CLK_bF$buf122),
    .D(_4310_),
    .Q(\datapath.registers.838[25] [13])
);

DFFPOSX1 _20163_ (
    .CLK(CLK_bF$buf121),
    .D(_4311_),
    .Q(\datapath.registers.838[25] [14])
);

DFFPOSX1 _20164_ (
    .CLK(CLK_bF$buf120),
    .D(_4312_),
    .Q(\datapath.registers.838[25] [15])
);

DFFPOSX1 _20165_ (
    .CLK(CLK_bF$buf119),
    .D(_4313_),
    .Q(\datapath.registers.838[25] [16])
);

DFFPOSX1 _20166_ (
    .CLK(CLK_bF$buf118),
    .D(_4314_),
    .Q(\datapath.registers.838[25] [17])
);

DFFPOSX1 _20167_ (
    .CLK(CLK_bF$buf117),
    .D(_4315_),
    .Q(\datapath.registers.838[25] [18])
);

DFFPOSX1 _20168_ (
    .CLK(CLK_bF$buf116),
    .D(_4316_),
    .Q(\datapath.registers.838[25] [19])
);

DFFPOSX1 _20169_ (
    .CLK(CLK_bF$buf115),
    .D(_4318_),
    .Q(\datapath.registers.838[25] [20])
);

DFFPOSX1 _20170_ (
    .CLK(CLK_bF$buf114),
    .D(_4319_),
    .Q(\datapath.registers.838[25] [21])
);

DFFPOSX1 _20171_ (
    .CLK(CLK_bF$buf113),
    .D(_4320_),
    .Q(\datapath.registers.838[25] [22])
);

DFFPOSX1 _20172_ (
    .CLK(CLK_bF$buf112),
    .D(_4321_),
    .Q(\datapath.registers.838[25] [23])
);

DFFPOSX1 _20173_ (
    .CLK(CLK_bF$buf111),
    .D(_4322_),
    .Q(\datapath.registers.838[25] [24])
);

DFFPOSX1 _20174_ (
    .CLK(CLK_bF$buf110),
    .D(_4323_),
    .Q(\datapath.registers.838[25] [25])
);

DFFPOSX1 _20175_ (
    .CLK(CLK_bF$buf109),
    .D(_4324_),
    .Q(\datapath.registers.838[25] [26])
);

DFFPOSX1 _20176_ (
    .CLK(CLK_bF$buf108),
    .D(_4325_),
    .Q(\datapath.registers.838[25] [27])
);

DFFPOSX1 _20177_ (
    .CLK(CLK_bF$buf107),
    .D(_4326_),
    .Q(\datapath.registers.838[25] [28])
);

DFFPOSX1 _20178_ (
    .CLK(CLK_bF$buf106),
    .D(_4327_),
    .Q(\datapath.registers.838[25] [29])
);

DFFPOSX1 _20179_ (
    .CLK(CLK_bF$buf105),
    .D(_4329_),
    .Q(\datapath.registers.838[25] [30])
);

DFFPOSX1 _20180_ (
    .CLK(CLK_bF$buf104),
    .D(_4330_),
    .Q(\datapath.registers.838[25] [31])
);

DFFPOSX1 _20181_ (
    .CLK(CLK_bF$buf103),
    .D(_3986_),
    .Q(\datapath.registers.838[16] [0])
);

DFFPOSX1 _20182_ (
    .CLK(CLK_bF$buf102),
    .D(_3997_),
    .Q(\datapath.registers.838[16] [1])
);

DFFPOSX1 _20183_ (
    .CLK(CLK_bF$buf101),
    .D(_4008_),
    .Q(\datapath.registers.838[16] [2])
);

DFFPOSX1 _20184_ (
    .CLK(CLK_bF$buf100),
    .D(_4011_),
    .Q(\datapath.registers.838[16] [3])
);

DFFPOSX1 _20185_ (
    .CLK(CLK_bF$buf99),
    .D(_4012_),
    .Q(\datapath.registers.838[16] [4])
);

DFFPOSX1 _20186_ (
    .CLK(CLK_bF$buf98),
    .D(_4013_),
    .Q(\datapath.registers.838[16] [5])
);

DFFPOSX1 _20187_ (
    .CLK(CLK_bF$buf97),
    .D(_4014_),
    .Q(\datapath.registers.838[16] [6])
);

DFFPOSX1 _20188_ (
    .CLK(CLK_bF$buf96),
    .D(_4015_),
    .Q(\datapath.registers.838[16] [7])
);

DFFPOSX1 _20189_ (
    .CLK(CLK_bF$buf95),
    .D(_4016_),
    .Q(\datapath.registers.838[16] [8])
);

DFFPOSX1 _20190_ (
    .CLK(CLK_bF$buf94),
    .D(_4017_),
    .Q(\datapath.registers.838[16] [9])
);

DFFPOSX1 _20191_ (
    .CLK(CLK_bF$buf93),
    .D(_3987_),
    .Q(\datapath.registers.838[16] [10])
);

DFFPOSX1 _20192_ (
    .CLK(CLK_bF$buf92),
    .D(_3988_),
    .Q(\datapath.registers.838[16] [11])
);

DFFPOSX1 _20193_ (
    .CLK(CLK_bF$buf91),
    .D(_3989_),
    .Q(\datapath.registers.838[16] [12])
);

DFFPOSX1 _20194_ (
    .CLK(CLK_bF$buf90),
    .D(_3990_),
    .Q(\datapath.registers.838[16] [13])
);

DFFPOSX1 _20195_ (
    .CLK(CLK_bF$buf89),
    .D(_3991_),
    .Q(\datapath.registers.838[16] [14])
);

DFFPOSX1 _20196_ (
    .CLK(CLK_bF$buf88),
    .D(_3992_),
    .Q(\datapath.registers.838[16] [15])
);

DFFPOSX1 _20197_ (
    .CLK(CLK_bF$buf87),
    .D(_3993_),
    .Q(\datapath.registers.838[16] [16])
);

DFFPOSX1 _20198_ (
    .CLK(CLK_bF$buf86),
    .D(_3994_),
    .Q(\datapath.registers.838[16] [17])
);

DFFPOSX1 _20199_ (
    .CLK(CLK_bF$buf85),
    .D(_3995_),
    .Q(\datapath.registers.838[16] [18])
);

DFFPOSX1 _20200_ (
    .CLK(CLK_bF$buf84),
    .D(_3996_),
    .Q(\datapath.registers.838[16] [19])
);

DFFPOSX1 _20201_ (
    .CLK(CLK_bF$buf83),
    .D(_3998_),
    .Q(\datapath.registers.838[16] [20])
);

DFFPOSX1 _20202_ (
    .CLK(CLK_bF$buf82),
    .D(_3999_),
    .Q(\datapath.registers.838[16] [21])
);

DFFPOSX1 _20203_ (
    .CLK(CLK_bF$buf81),
    .D(_4000_),
    .Q(\datapath.registers.838[16] [22])
);

DFFPOSX1 _20204_ (
    .CLK(CLK_bF$buf80),
    .D(_4001_),
    .Q(\datapath.registers.838[16] [23])
);

DFFPOSX1 _20205_ (
    .CLK(CLK_bF$buf79),
    .D(_4002_),
    .Q(\datapath.registers.838[16] [24])
);

DFFPOSX1 _20206_ (
    .CLK(CLK_bF$buf78),
    .D(_4003_),
    .Q(\datapath.registers.838[16] [25])
);

DFFPOSX1 _20207_ (
    .CLK(CLK_bF$buf77),
    .D(_4004_),
    .Q(\datapath.registers.838[16] [26])
);

DFFPOSX1 _20208_ (
    .CLK(CLK_bF$buf76),
    .D(_4005_),
    .Q(\datapath.registers.838[16] [27])
);

DFFPOSX1 _20209_ (
    .CLK(CLK_bF$buf75),
    .D(_4006_),
    .Q(\datapath.registers.838[16] [28])
);

DFFPOSX1 _20210_ (
    .CLK(CLK_bF$buf74),
    .D(_4007_),
    .Q(\datapath.registers.838[16] [29])
);

DFFPOSX1 _20211_ (
    .CLK(CLK_bF$buf73),
    .D(_4009_),
    .Q(\datapath.registers.838[16] [30])
);

DFFPOSX1 _20212_ (
    .CLK(CLK_bF$buf72),
    .D(_4010_),
    .Q(\datapath.registers.838[16] [31])
);

DFFPOSX1 _20213_ (
    .CLK(CLK_bF$buf71),
    .D(_4466_),
    .Q(\datapath.registers.838[2] [0])
);

DFFPOSX1 _20214_ (
    .CLK(CLK_bF$buf70),
    .D(_4477_),
    .Q(\datapath.registers.838[2] [1])
);

DFFPOSX1 _20215_ (
    .CLK(CLK_bF$buf69),
    .D(_4488_),
    .Q(\datapath.registers.838[2] [2])
);

DFFPOSX1 _20216_ (
    .CLK(CLK_bF$buf68),
    .D(_4491_),
    .Q(\datapath.registers.838[2] [3])
);

DFFPOSX1 _20217_ (
    .CLK(CLK_bF$buf67),
    .D(_4492_),
    .Q(\datapath.registers.838[2] [4])
);

DFFPOSX1 _20218_ (
    .CLK(CLK_bF$buf66),
    .D(_4493_),
    .Q(\datapath.registers.838[2] [5])
);

DFFPOSX1 _20219_ (
    .CLK(CLK_bF$buf65),
    .D(_4494_),
    .Q(\datapath.registers.838[2] [6])
);

DFFPOSX1 _20220_ (
    .CLK(CLK_bF$buf64),
    .D(_4495_),
    .Q(\datapath.registers.838[2] [7])
);

DFFPOSX1 _20221_ (
    .CLK(CLK_bF$buf63),
    .D(_4496_),
    .Q(\datapath.registers.838[2] [8])
);

DFFPOSX1 _20222_ (
    .CLK(CLK_bF$buf62),
    .D(_4497_),
    .Q(\datapath.registers.838[2] [9])
);

DFFPOSX1 _20223_ (
    .CLK(CLK_bF$buf61),
    .D(_4467_),
    .Q(\datapath.registers.838[2] [10])
);

DFFPOSX1 _20224_ (
    .CLK(CLK_bF$buf60),
    .D(_4468_),
    .Q(\datapath.registers.838[2] [11])
);

DFFPOSX1 _20225_ (
    .CLK(CLK_bF$buf59),
    .D(_4469_),
    .Q(\datapath.registers.838[2] [12])
);

DFFPOSX1 _20226_ (
    .CLK(CLK_bF$buf58),
    .D(_4470_),
    .Q(\datapath.registers.838[2] [13])
);

DFFPOSX1 _20227_ (
    .CLK(CLK_bF$buf57),
    .D(_4471_),
    .Q(\datapath.registers.838[2] [14])
);

DFFPOSX1 _20228_ (
    .CLK(CLK_bF$buf56),
    .D(_4472_),
    .Q(\datapath.registers.838[2] [15])
);

DFFPOSX1 _20229_ (
    .CLK(CLK_bF$buf55),
    .D(_4473_),
    .Q(\datapath.registers.838[2] [16])
);

DFFPOSX1 _20230_ (
    .CLK(CLK_bF$buf54),
    .D(_4474_),
    .Q(\datapath.registers.838[2] [17])
);

DFFPOSX1 _20231_ (
    .CLK(CLK_bF$buf53),
    .D(_4475_),
    .Q(\datapath.registers.838[2] [18])
);

DFFPOSX1 _20232_ (
    .CLK(CLK_bF$buf52),
    .D(_4476_),
    .Q(\datapath.registers.838[2] [19])
);

DFFPOSX1 _20233_ (
    .CLK(CLK_bF$buf51),
    .D(_4478_),
    .Q(\datapath.registers.838[2] [20])
);

DFFPOSX1 _20234_ (
    .CLK(CLK_bF$buf50),
    .D(_4479_),
    .Q(\datapath.registers.838[2] [21])
);

DFFPOSX1 _20235_ (
    .CLK(CLK_bF$buf49),
    .D(_4480_),
    .Q(\datapath.registers.838[2] [22])
);

DFFPOSX1 _20236_ (
    .CLK(CLK_bF$buf48),
    .D(_4481_),
    .Q(\datapath.registers.838[2] [23])
);

DFFPOSX1 _20237_ (
    .CLK(CLK_bF$buf47),
    .D(_4482_),
    .Q(\datapath.registers.838[2] [24])
);

DFFPOSX1 _20238_ (
    .CLK(CLK_bF$buf46),
    .D(_4483_),
    .Q(\datapath.registers.838[2] [25])
);

DFFPOSX1 _20239_ (
    .CLK(CLK_bF$buf45),
    .D(_4484_),
    .Q(\datapath.registers.838[2] [26])
);

DFFPOSX1 _20240_ (
    .CLK(CLK_bF$buf44),
    .D(_4485_),
    .Q(\datapath.registers.838[2] [27])
);

DFFPOSX1 _20241_ (
    .CLK(CLK_bF$buf43),
    .D(_4486_),
    .Q(\datapath.registers.838[2] [28])
);

DFFPOSX1 _20242_ (
    .CLK(CLK_bF$buf42),
    .D(_4487_),
    .Q(\datapath.registers.838[2] [29])
);

DFFPOSX1 _20243_ (
    .CLK(CLK_bF$buf41),
    .D(_4489_),
    .Q(\datapath.registers.838[2] [30])
);

DFFPOSX1 _20244_ (
    .CLK(CLK_bF$buf40),
    .D(_4490_),
    .Q(\datapath.registers.838[2] [31])
);

DFFPOSX1 _20245_ (
    .CLK(CLK_bF$buf39),
    .D(_4274_),
    .Q(\datapath.registers.838[24] [0])
);

DFFPOSX1 _20246_ (
    .CLK(CLK_bF$buf38),
    .D(_4285_),
    .Q(\datapath.registers.838[24] [1])
);

DFFPOSX1 _20247_ (
    .CLK(CLK_bF$buf37),
    .D(_4296_),
    .Q(\datapath.registers.838[24] [2])
);

DFFPOSX1 _20248_ (
    .CLK(CLK_bF$buf36),
    .D(_4299_),
    .Q(\datapath.registers.838[24] [3])
);

DFFPOSX1 _20249_ (
    .CLK(CLK_bF$buf35),
    .D(_4300_),
    .Q(\datapath.registers.838[24] [4])
);

DFFPOSX1 _20250_ (
    .CLK(CLK_bF$buf34),
    .D(_4301_),
    .Q(\datapath.registers.838[24] [5])
);

DFFPOSX1 _20251_ (
    .CLK(CLK_bF$buf33),
    .D(_4302_),
    .Q(\datapath.registers.838[24] [6])
);

DFFPOSX1 _20252_ (
    .CLK(CLK_bF$buf32),
    .D(_4303_),
    .Q(\datapath.registers.838[24] [7])
);

DFFPOSX1 _20253_ (
    .CLK(CLK_bF$buf31),
    .D(_4304_),
    .Q(\datapath.registers.838[24] [8])
);

DFFPOSX1 _20254_ (
    .CLK(CLK_bF$buf30),
    .D(_4305_),
    .Q(\datapath.registers.838[24] [9])
);

DFFPOSX1 _20255_ (
    .CLK(CLK_bF$buf29),
    .D(_4275_),
    .Q(\datapath.registers.838[24] [10])
);

DFFPOSX1 _20256_ (
    .CLK(CLK_bF$buf28),
    .D(_4276_),
    .Q(\datapath.registers.838[24] [11])
);

DFFPOSX1 _20257_ (
    .CLK(CLK_bF$buf27),
    .D(_4277_),
    .Q(\datapath.registers.838[24] [12])
);

DFFPOSX1 _20258_ (
    .CLK(CLK_bF$buf26),
    .D(_4278_),
    .Q(\datapath.registers.838[24] [13])
);

DFFPOSX1 _20259_ (
    .CLK(CLK_bF$buf25),
    .D(_4279_),
    .Q(\datapath.registers.838[24] [14])
);

DFFPOSX1 _20260_ (
    .CLK(CLK_bF$buf24),
    .D(_4280_),
    .Q(\datapath.registers.838[24] [15])
);

DFFPOSX1 _20261_ (
    .CLK(CLK_bF$buf23),
    .D(_4281_),
    .Q(\datapath.registers.838[24] [16])
);

DFFPOSX1 _20262_ (
    .CLK(CLK_bF$buf22),
    .D(_4282_),
    .Q(\datapath.registers.838[24] [17])
);

DFFPOSX1 _20263_ (
    .CLK(CLK_bF$buf21),
    .D(_4283_),
    .Q(\datapath.registers.838[24] [18])
);

DFFPOSX1 _20264_ (
    .CLK(CLK_bF$buf20),
    .D(_4284_),
    .Q(\datapath.registers.838[24] [19])
);

DFFPOSX1 _20265_ (
    .CLK(CLK_bF$buf19),
    .D(_4286_),
    .Q(\datapath.registers.838[24] [20])
);

DFFPOSX1 _20266_ (
    .CLK(CLK_bF$buf18),
    .D(_4287_),
    .Q(\datapath.registers.838[24] [21])
);

DFFPOSX1 _20267_ (
    .CLK(CLK_bF$buf17),
    .D(_4288_),
    .Q(\datapath.registers.838[24] [22])
);

DFFPOSX1 _20268_ (
    .CLK(CLK_bF$buf16),
    .D(_4289_),
    .Q(\datapath.registers.838[24] [23])
);

DFFPOSX1 _20269_ (
    .CLK(CLK_bF$buf15),
    .D(_4290_),
    .Q(\datapath.registers.838[24] [24])
);

DFFPOSX1 _20270_ (
    .CLK(CLK_bF$buf14),
    .D(_4291_),
    .Q(\datapath.registers.838[24] [25])
);

DFFPOSX1 _20271_ (
    .CLK(CLK_bF$buf13),
    .D(_4292_),
    .Q(\datapath.registers.838[24] [26])
);

DFFPOSX1 _20272_ (
    .CLK(CLK_bF$buf12),
    .D(_4293_),
    .Q(\datapath.registers.838[24] [27])
);

DFFPOSX1 _20273_ (
    .CLK(CLK_bF$buf11),
    .D(_4294_),
    .Q(\datapath.registers.838[24] [28])
);

DFFPOSX1 _20274_ (
    .CLK(CLK_bF$buf10),
    .D(_4295_),
    .Q(\datapath.registers.838[24] [29])
);

DFFPOSX1 _20275_ (
    .CLK(CLK_bF$buf9),
    .D(_4297_),
    .Q(\datapath.registers.838[24] [30])
);

DFFPOSX1 _20276_ (
    .CLK(CLK_bF$buf8),
    .D(_4298_),
    .Q(\datapath.registers.838[24] [31])
);

DFFPOSX1 _20277_ (
    .CLK(CLK_bF$buf7),
    .D(_4210_),
    .Q(\datapath.registers.838[22] [0])
);

DFFPOSX1 _20278_ (
    .CLK(CLK_bF$buf6),
    .D(_4221_),
    .Q(\datapath.registers.838[22] [1])
);

DFFPOSX1 _20279_ (
    .CLK(CLK_bF$buf5),
    .D(_4232_),
    .Q(\datapath.registers.838[22] [2])
);

DFFPOSX1 _20280_ (
    .CLK(CLK_bF$buf4),
    .D(_4235_),
    .Q(\datapath.registers.838[22] [3])
);

DFFPOSX1 _20281_ (
    .CLK(CLK_bF$buf3),
    .D(_4236_),
    .Q(\datapath.registers.838[22] [4])
);

DFFPOSX1 _20282_ (
    .CLK(CLK_bF$buf2),
    .D(_4237_),
    .Q(\datapath.registers.838[22] [5])
);

DFFPOSX1 _20283_ (
    .CLK(CLK_bF$buf1),
    .D(_4238_),
    .Q(\datapath.registers.838[22] [6])
);

DFFPOSX1 _20284_ (
    .CLK(CLK_bF$buf0),
    .D(_4239_),
    .Q(\datapath.registers.838[22] [7])
);

DFFPOSX1 _20285_ (
    .CLK(CLK_bF$buf151),
    .D(_4240_),
    .Q(\datapath.registers.838[22] [8])
);

DFFPOSX1 _20286_ (
    .CLK(CLK_bF$buf150),
    .D(_4241_),
    .Q(\datapath.registers.838[22] [9])
);

DFFPOSX1 _20287_ (
    .CLK(CLK_bF$buf149),
    .D(_4211_),
    .Q(\datapath.registers.838[22] [10])
);

DFFPOSX1 _20288_ (
    .CLK(CLK_bF$buf148),
    .D(_4212_),
    .Q(\datapath.registers.838[22] [11])
);

DFFPOSX1 _20289_ (
    .CLK(CLK_bF$buf147),
    .D(_4213_),
    .Q(\datapath.registers.838[22] [12])
);

DFFPOSX1 _20290_ (
    .CLK(CLK_bF$buf146),
    .D(_4214_),
    .Q(\datapath.registers.838[22] [13])
);

DFFPOSX1 _20291_ (
    .CLK(CLK_bF$buf145),
    .D(_4215_),
    .Q(\datapath.registers.838[22] [14])
);

DFFPOSX1 _20292_ (
    .CLK(CLK_bF$buf144),
    .D(_4216_),
    .Q(\datapath.registers.838[22] [15])
);

DFFPOSX1 _20293_ (
    .CLK(CLK_bF$buf143),
    .D(_4217_),
    .Q(\datapath.registers.838[22] [16])
);

DFFPOSX1 _20294_ (
    .CLK(CLK_bF$buf142),
    .D(_4218_),
    .Q(\datapath.registers.838[22] [17])
);

DFFPOSX1 _20295_ (
    .CLK(CLK_bF$buf141),
    .D(_4219_),
    .Q(\datapath.registers.838[22] [18])
);

DFFPOSX1 _20296_ (
    .CLK(CLK_bF$buf140),
    .D(_4220_),
    .Q(\datapath.registers.838[22] [19])
);

DFFPOSX1 _20297_ (
    .CLK(CLK_bF$buf139),
    .D(_4222_),
    .Q(\datapath.registers.838[22] [20])
);

DFFPOSX1 _20298_ (
    .CLK(CLK_bF$buf138),
    .D(_4223_),
    .Q(\datapath.registers.838[22] [21])
);

DFFPOSX1 _20299_ (
    .CLK(CLK_bF$buf137),
    .D(_4224_),
    .Q(\datapath.registers.838[22] [22])
);

DFFPOSX1 _20300_ (
    .CLK(CLK_bF$buf136),
    .D(_4225_),
    .Q(\datapath.registers.838[22] [23])
);

DFFPOSX1 _20301_ (
    .CLK(CLK_bF$buf135),
    .D(_4226_),
    .Q(\datapath.registers.838[22] [24])
);

DFFPOSX1 _20302_ (
    .CLK(CLK_bF$buf134),
    .D(_4227_),
    .Q(\datapath.registers.838[22] [25])
);

DFFPOSX1 _20303_ (
    .CLK(CLK_bF$buf133),
    .D(_4228_),
    .Q(\datapath.registers.838[22] [26])
);

DFFPOSX1 _20304_ (
    .CLK(CLK_bF$buf132),
    .D(_4229_),
    .Q(\datapath.registers.838[22] [27])
);

DFFPOSX1 _20305_ (
    .CLK(CLK_bF$buf131),
    .D(_4230_),
    .Q(\datapath.registers.838[22] [28])
);

DFFPOSX1 _20306_ (
    .CLK(CLK_bF$buf130),
    .D(_4231_),
    .Q(\datapath.registers.838[22] [29])
);

DFFPOSX1 _20307_ (
    .CLK(CLK_bF$buf129),
    .D(_4233_),
    .Q(\datapath.registers.838[22] [30])
);

DFFPOSX1 _20308_ (
    .CLK(CLK_bF$buf128),
    .D(_4234_),
    .Q(\datapath.registers.838[22] [31])
);

DFFPOSX1 _20309_ (
    .CLK(CLK_bF$buf127),
    .D(_4594_),
    .Q(\datapath.registers.838[4] [0])
);

DFFPOSX1 _20310_ (
    .CLK(CLK_bF$buf126),
    .D(_4605_),
    .Q(\datapath.registers.838[4] [1])
);

DFFPOSX1 _20311_ (
    .CLK(CLK_bF$buf125),
    .D(_4616_),
    .Q(\datapath.registers.838[4] [2])
);

DFFPOSX1 _20312_ (
    .CLK(CLK_bF$buf124),
    .D(_4619_),
    .Q(\datapath.registers.838[4] [3])
);

DFFPOSX1 _20313_ (
    .CLK(CLK_bF$buf123),
    .D(_4620_),
    .Q(\datapath.registers.838[4] [4])
);

DFFPOSX1 _20314_ (
    .CLK(CLK_bF$buf122),
    .D(_4621_),
    .Q(\datapath.registers.838[4] [5])
);

DFFPOSX1 _20315_ (
    .CLK(CLK_bF$buf121),
    .D(_4622_),
    .Q(\datapath.registers.838[4] [6])
);

DFFPOSX1 _20316_ (
    .CLK(CLK_bF$buf120),
    .D(_4623_),
    .Q(\datapath.registers.838[4] [7])
);

DFFPOSX1 _20317_ (
    .CLK(CLK_bF$buf119),
    .D(_4624_),
    .Q(\datapath.registers.838[4] [8])
);

DFFPOSX1 _20318_ (
    .CLK(CLK_bF$buf118),
    .D(_4625_),
    .Q(\datapath.registers.838[4] [9])
);

DFFPOSX1 _20319_ (
    .CLK(CLK_bF$buf117),
    .D(_4595_),
    .Q(\datapath.registers.838[4] [10])
);

DFFPOSX1 _20320_ (
    .CLK(CLK_bF$buf116),
    .D(_4596_),
    .Q(\datapath.registers.838[4] [11])
);

DFFPOSX1 _20321_ (
    .CLK(CLK_bF$buf115),
    .D(_4597_),
    .Q(\datapath.registers.838[4] [12])
);

DFFPOSX1 _20322_ (
    .CLK(CLK_bF$buf114),
    .D(_4598_),
    .Q(\datapath.registers.838[4] [13])
);

DFFPOSX1 _20323_ (
    .CLK(CLK_bF$buf113),
    .D(_4599_),
    .Q(\datapath.registers.838[4] [14])
);

DFFPOSX1 _20324_ (
    .CLK(CLK_bF$buf112),
    .D(_4600_),
    .Q(\datapath.registers.838[4] [15])
);

DFFPOSX1 _20325_ (
    .CLK(CLK_bF$buf111),
    .D(_4601_),
    .Q(\datapath.registers.838[4] [16])
);

DFFPOSX1 _20326_ (
    .CLK(CLK_bF$buf110),
    .D(_4602_),
    .Q(\datapath.registers.838[4] [17])
);

DFFPOSX1 _20327_ (
    .CLK(CLK_bF$buf109),
    .D(_4603_),
    .Q(\datapath.registers.838[4] [18])
);

DFFPOSX1 _20328_ (
    .CLK(CLK_bF$buf108),
    .D(_4604_),
    .Q(\datapath.registers.838[4] [19])
);

DFFPOSX1 _20329_ (
    .CLK(CLK_bF$buf107),
    .D(_4606_),
    .Q(\datapath.registers.838[4] [20])
);

DFFPOSX1 _20330_ (
    .CLK(CLK_bF$buf106),
    .D(_4607_),
    .Q(\datapath.registers.838[4] [21])
);

DFFPOSX1 _20331_ (
    .CLK(CLK_bF$buf105),
    .D(_4608_),
    .Q(\datapath.registers.838[4] [22])
);

DFFPOSX1 _20332_ (
    .CLK(CLK_bF$buf104),
    .D(_4609_),
    .Q(\datapath.registers.838[4] [23])
);

DFFPOSX1 _20333_ (
    .CLK(CLK_bF$buf103),
    .D(_4610_),
    .Q(\datapath.registers.838[4] [24])
);

DFFPOSX1 _20334_ (
    .CLK(CLK_bF$buf102),
    .D(_4611_),
    .Q(\datapath.registers.838[4] [25])
);

DFFPOSX1 _20335_ (
    .CLK(CLK_bF$buf101),
    .D(_4612_),
    .Q(\datapath.registers.838[4] [26])
);

DFFPOSX1 _20336_ (
    .CLK(CLK_bF$buf100),
    .D(_4613_),
    .Q(\datapath.registers.838[4] [27])
);

DFFPOSX1 _20337_ (
    .CLK(CLK_bF$buf99),
    .D(_4614_),
    .Q(\datapath.registers.838[4] [28])
);

DFFPOSX1 _20338_ (
    .CLK(CLK_bF$buf98),
    .D(_4615_),
    .Q(\datapath.registers.838[4] [29])
);

DFFPOSX1 _20339_ (
    .CLK(CLK_bF$buf97),
    .D(_4617_),
    .Q(\datapath.registers.838[4] [30])
);

DFFPOSX1 _20340_ (
    .CLK(CLK_bF$buf96),
    .D(_4618_),
    .Q(\datapath.registers.838[4] [31])
);

DFFPOSX1 _20341_ (
    .CLK(CLK_bF$buf95),
    .D(_4690_),
    .Q(\datapath.registers.838[7] [0])
);

DFFPOSX1 _20342_ (
    .CLK(CLK_bF$buf94),
    .D(_4701_),
    .Q(\datapath.registers.838[7] [1])
);

DFFPOSX1 _20343_ (
    .CLK(CLK_bF$buf93),
    .D(_4712_),
    .Q(\datapath.registers.838[7] [2])
);

DFFPOSX1 _20344_ (
    .CLK(CLK_bF$buf92),
    .D(_4715_),
    .Q(\datapath.registers.838[7] [3])
);

DFFPOSX1 _20345_ (
    .CLK(CLK_bF$buf91),
    .D(_4716_),
    .Q(\datapath.registers.838[7] [4])
);

DFFPOSX1 _20346_ (
    .CLK(CLK_bF$buf90),
    .D(_4717_),
    .Q(\datapath.registers.838[7] [5])
);

DFFPOSX1 _20347_ (
    .CLK(CLK_bF$buf89),
    .D(_4718_),
    .Q(\datapath.registers.838[7] [6])
);

DFFPOSX1 _20348_ (
    .CLK(CLK_bF$buf88),
    .D(_4719_),
    .Q(\datapath.registers.838[7] [7])
);

DFFPOSX1 _20349_ (
    .CLK(CLK_bF$buf87),
    .D(_4720_),
    .Q(\datapath.registers.838[7] [8])
);

DFFPOSX1 _20350_ (
    .CLK(CLK_bF$buf86),
    .D(_4721_),
    .Q(\datapath.registers.838[7] [9])
);

DFFPOSX1 _20351_ (
    .CLK(CLK_bF$buf85),
    .D(_4691_),
    .Q(\datapath.registers.838[7] [10])
);

DFFPOSX1 _20352_ (
    .CLK(CLK_bF$buf84),
    .D(_4692_),
    .Q(\datapath.registers.838[7] [11])
);

DFFPOSX1 _20353_ (
    .CLK(CLK_bF$buf83),
    .D(_4693_),
    .Q(\datapath.registers.838[7] [12])
);

DFFPOSX1 _20354_ (
    .CLK(CLK_bF$buf82),
    .D(_4694_),
    .Q(\datapath.registers.838[7] [13])
);

DFFPOSX1 _20355_ (
    .CLK(CLK_bF$buf81),
    .D(_4695_),
    .Q(\datapath.registers.838[7] [14])
);

DFFPOSX1 _20356_ (
    .CLK(CLK_bF$buf80),
    .D(_4696_),
    .Q(\datapath.registers.838[7] [15])
);

DFFPOSX1 _20357_ (
    .CLK(CLK_bF$buf79),
    .D(_4697_),
    .Q(\datapath.registers.838[7] [16])
);

DFFPOSX1 _20358_ (
    .CLK(CLK_bF$buf78),
    .D(_4698_),
    .Q(\datapath.registers.838[7] [17])
);

DFFPOSX1 _20359_ (
    .CLK(CLK_bF$buf77),
    .D(_4699_),
    .Q(\datapath.registers.838[7] [18])
);

DFFPOSX1 _20360_ (
    .CLK(CLK_bF$buf76),
    .D(_4700_),
    .Q(\datapath.registers.838[7] [19])
);

DFFPOSX1 _20361_ (
    .CLK(CLK_bF$buf75),
    .D(_4702_),
    .Q(\datapath.registers.838[7] [20])
);

DFFPOSX1 _20362_ (
    .CLK(CLK_bF$buf74),
    .D(_4703_),
    .Q(\datapath.registers.838[7] [21])
);

DFFPOSX1 _20363_ (
    .CLK(CLK_bF$buf73),
    .D(_4704_),
    .Q(\datapath.registers.838[7] [22])
);

DFFPOSX1 _20364_ (
    .CLK(CLK_bF$buf72),
    .D(_4705_),
    .Q(\datapath.registers.838[7] [23])
);

DFFPOSX1 _20365_ (
    .CLK(CLK_bF$buf71),
    .D(_4706_),
    .Q(\datapath.registers.838[7] [24])
);

DFFPOSX1 _20366_ (
    .CLK(CLK_bF$buf70),
    .D(_4707_),
    .Q(\datapath.registers.838[7] [25])
);

DFFPOSX1 _20367_ (
    .CLK(CLK_bF$buf69),
    .D(_4708_),
    .Q(\datapath.registers.838[7] [26])
);

DFFPOSX1 _20368_ (
    .CLK(CLK_bF$buf68),
    .D(_4709_),
    .Q(\datapath.registers.838[7] [27])
);

DFFPOSX1 _20369_ (
    .CLK(CLK_bF$buf67),
    .D(_4710_),
    .Q(\datapath.registers.838[7] [28])
);

DFFPOSX1 _20370_ (
    .CLK(CLK_bF$buf66),
    .D(_4711_),
    .Q(\datapath.registers.838[7] [29])
);

DFFPOSX1 _20371_ (
    .CLK(CLK_bF$buf65),
    .D(_4713_),
    .Q(\datapath.registers.838[7] [30])
);

DFFPOSX1 _20372_ (
    .CLK(CLK_bF$buf64),
    .D(_4714_),
    .Q(\datapath.registers.838[7] [31])
);

DFFPOSX1 _20373_ (
    .CLK(CLK_bF$buf63),
    .D(_3890_),
    .Q(\datapath.registers.838[13] [0])
);

DFFPOSX1 _20374_ (
    .CLK(CLK_bF$buf62),
    .D(_3901_),
    .Q(\datapath.registers.838[13] [1])
);

DFFPOSX1 _20375_ (
    .CLK(CLK_bF$buf61),
    .D(_3912_),
    .Q(\datapath.registers.838[13] [2])
);

DFFPOSX1 _20376_ (
    .CLK(CLK_bF$buf60),
    .D(_3915_),
    .Q(\datapath.registers.838[13] [3])
);

DFFPOSX1 _20377_ (
    .CLK(CLK_bF$buf59),
    .D(_3916_),
    .Q(\datapath.registers.838[13] [4])
);

DFFPOSX1 _20378_ (
    .CLK(CLK_bF$buf58),
    .D(_3917_),
    .Q(\datapath.registers.838[13] [5])
);

DFFPOSX1 _20379_ (
    .CLK(CLK_bF$buf57),
    .D(_3918_),
    .Q(\datapath.registers.838[13] [6])
);

DFFPOSX1 _20380_ (
    .CLK(CLK_bF$buf56),
    .D(_3919_),
    .Q(\datapath.registers.838[13] [7])
);

DFFPOSX1 _20381_ (
    .CLK(CLK_bF$buf55),
    .D(_3920_),
    .Q(\datapath.registers.838[13] [8])
);

DFFPOSX1 _20382_ (
    .CLK(CLK_bF$buf54),
    .D(_3921_),
    .Q(\datapath.registers.838[13] [9])
);

DFFPOSX1 _20383_ (
    .CLK(CLK_bF$buf53),
    .D(_3891_),
    .Q(\datapath.registers.838[13] [10])
);

DFFPOSX1 _20384_ (
    .CLK(CLK_bF$buf52),
    .D(_3892_),
    .Q(\datapath.registers.838[13] [11])
);

DFFPOSX1 _20385_ (
    .CLK(CLK_bF$buf51),
    .D(_3893_),
    .Q(\datapath.registers.838[13] [12])
);

DFFPOSX1 _20386_ (
    .CLK(CLK_bF$buf50),
    .D(_3894_),
    .Q(\datapath.registers.838[13] [13])
);

DFFPOSX1 _20387_ (
    .CLK(CLK_bF$buf49),
    .D(_3895_),
    .Q(\datapath.registers.838[13] [14])
);

DFFPOSX1 _20388_ (
    .CLK(CLK_bF$buf48),
    .D(_3896_),
    .Q(\datapath.registers.838[13] [15])
);

DFFPOSX1 _20389_ (
    .CLK(CLK_bF$buf47),
    .D(_3897_),
    .Q(\datapath.registers.838[13] [16])
);

DFFPOSX1 _20390_ (
    .CLK(CLK_bF$buf46),
    .D(_3898_),
    .Q(\datapath.registers.838[13] [17])
);

DFFPOSX1 _20391_ (
    .CLK(CLK_bF$buf45),
    .D(_3899_),
    .Q(\datapath.registers.838[13] [18])
);

DFFPOSX1 _20392_ (
    .CLK(CLK_bF$buf44),
    .D(_3900_),
    .Q(\datapath.registers.838[13] [19])
);

DFFPOSX1 _20393_ (
    .CLK(CLK_bF$buf43),
    .D(_3902_),
    .Q(\datapath.registers.838[13] [20])
);

DFFPOSX1 _20394_ (
    .CLK(CLK_bF$buf42),
    .D(_3903_),
    .Q(\datapath.registers.838[13] [21])
);

DFFPOSX1 _20395_ (
    .CLK(CLK_bF$buf41),
    .D(_3904_),
    .Q(\datapath.registers.838[13] [22])
);

DFFPOSX1 _20396_ (
    .CLK(CLK_bF$buf40),
    .D(_3905_),
    .Q(\datapath.registers.838[13] [23])
);

DFFPOSX1 _20397_ (
    .CLK(CLK_bF$buf39),
    .D(_3906_),
    .Q(\datapath.registers.838[13] [24])
);

DFFPOSX1 _20398_ (
    .CLK(CLK_bF$buf38),
    .D(_3907_),
    .Q(\datapath.registers.838[13] [25])
);

DFFPOSX1 _20399_ (
    .CLK(CLK_bF$buf37),
    .D(_3908_),
    .Q(\datapath.registers.838[13] [26])
);

DFFPOSX1 _20400_ (
    .CLK(CLK_bF$buf36),
    .D(_3909_),
    .Q(\datapath.registers.838[13] [27])
);

DFFPOSX1 _20401_ (
    .CLK(CLK_bF$buf35),
    .D(_3910_),
    .Q(\datapath.registers.838[13] [28])
);

DFFPOSX1 _20402_ (
    .CLK(CLK_bF$buf34),
    .D(_3911_),
    .Q(\datapath.registers.838[13] [29])
);

DFFPOSX1 _20403_ (
    .CLK(CLK_bF$buf33),
    .D(_3913_),
    .Q(\datapath.registers.838[13] [30])
);

DFFPOSX1 _20404_ (
    .CLK(CLK_bF$buf32),
    .D(_3914_),
    .Q(\datapath.registers.838[13] [31])
);

DFFPOSX1 _20405_ (
    .CLK(CLK_bF$buf31),
    .D(_3858_),
    .Q(\datapath.registers.838[12] [0])
);

DFFPOSX1 _20406_ (
    .CLK(CLK_bF$buf30),
    .D(_3869_),
    .Q(\datapath.registers.838[12] [1])
);

DFFPOSX1 _20407_ (
    .CLK(CLK_bF$buf29),
    .D(_3880_),
    .Q(\datapath.registers.838[12] [2])
);

DFFPOSX1 _20408_ (
    .CLK(CLK_bF$buf28),
    .D(_3883_),
    .Q(\datapath.registers.838[12] [3])
);

DFFPOSX1 _20409_ (
    .CLK(CLK_bF$buf27),
    .D(_3884_),
    .Q(\datapath.registers.838[12] [4])
);

DFFPOSX1 _20410_ (
    .CLK(CLK_bF$buf26),
    .D(_3885_),
    .Q(\datapath.registers.838[12] [5])
);

DFFPOSX1 _20411_ (
    .CLK(CLK_bF$buf25),
    .D(_3886_),
    .Q(\datapath.registers.838[12] [6])
);

DFFPOSX1 _20412_ (
    .CLK(CLK_bF$buf24),
    .D(_3887_),
    .Q(\datapath.registers.838[12] [7])
);

DFFPOSX1 _20413_ (
    .CLK(CLK_bF$buf23),
    .D(_3888_),
    .Q(\datapath.registers.838[12] [8])
);

DFFPOSX1 _20414_ (
    .CLK(CLK_bF$buf22),
    .D(_3889_),
    .Q(\datapath.registers.838[12] [9])
);

DFFPOSX1 _20415_ (
    .CLK(CLK_bF$buf21),
    .D(_3859_),
    .Q(\datapath.registers.838[12] [10])
);

DFFPOSX1 _20416_ (
    .CLK(CLK_bF$buf20),
    .D(_3860_),
    .Q(\datapath.registers.838[12] [11])
);

DFFPOSX1 _20417_ (
    .CLK(CLK_bF$buf19),
    .D(_3861_),
    .Q(\datapath.registers.838[12] [12])
);

DFFPOSX1 _20418_ (
    .CLK(CLK_bF$buf18),
    .D(_3862_),
    .Q(\datapath.registers.838[12] [13])
);

DFFPOSX1 _20419_ (
    .CLK(CLK_bF$buf17),
    .D(_3863_),
    .Q(\datapath.registers.838[12] [14])
);

DFFPOSX1 _20420_ (
    .CLK(CLK_bF$buf16),
    .D(_3864_),
    .Q(\datapath.registers.838[12] [15])
);

DFFPOSX1 _20421_ (
    .CLK(CLK_bF$buf15),
    .D(_3865_),
    .Q(\datapath.registers.838[12] [16])
);

DFFPOSX1 _20422_ (
    .CLK(CLK_bF$buf14),
    .D(_3866_),
    .Q(\datapath.registers.838[12] [17])
);

DFFPOSX1 _20423_ (
    .CLK(CLK_bF$buf13),
    .D(_3867_),
    .Q(\datapath.registers.838[12] [18])
);

DFFPOSX1 _20424_ (
    .CLK(CLK_bF$buf12),
    .D(_3868_),
    .Q(\datapath.registers.838[12] [19])
);

DFFPOSX1 _20425_ (
    .CLK(CLK_bF$buf11),
    .D(_3870_),
    .Q(\datapath.registers.838[12] [20])
);

DFFPOSX1 _20426_ (
    .CLK(CLK_bF$buf10),
    .D(_3871_),
    .Q(\datapath.registers.838[12] [21])
);

DFFPOSX1 _20427_ (
    .CLK(CLK_bF$buf9),
    .D(_3872_),
    .Q(\datapath.registers.838[12] [22])
);

DFFPOSX1 _20428_ (
    .CLK(CLK_bF$buf8),
    .D(_3873_),
    .Q(\datapath.registers.838[12] [23])
);

DFFPOSX1 _20429_ (
    .CLK(CLK_bF$buf7),
    .D(_3874_),
    .Q(\datapath.registers.838[12] [24])
);

DFFPOSX1 _20430_ (
    .CLK(CLK_bF$buf6),
    .D(_3875_),
    .Q(\datapath.registers.838[12] [25])
);

DFFPOSX1 _20431_ (
    .CLK(CLK_bF$buf5),
    .D(_3876_),
    .Q(\datapath.registers.838[12] [26])
);

DFFPOSX1 _20432_ (
    .CLK(CLK_bF$buf4),
    .D(_3877_),
    .Q(\datapath.registers.838[12] [27])
);

DFFPOSX1 _20433_ (
    .CLK(CLK_bF$buf3),
    .D(_3878_),
    .Q(\datapath.registers.838[12] [28])
);

DFFPOSX1 _20434_ (
    .CLK(CLK_bF$buf2),
    .D(_3879_),
    .Q(\datapath.registers.838[12] [29])
);

DFFPOSX1 _20435_ (
    .CLK(CLK_bF$buf1),
    .D(_3881_),
    .Q(\datapath.registers.838[12] [30])
);

DFFPOSX1 _20436_ (
    .CLK(CLK_bF$buf0),
    .D(_3882_),
    .Q(\datapath.registers.838[12] [31])
);

DFFPOSX1 _20437_ (
    .CLK(CLK_bF$buf151),
    .D(_3954_),
    .Q(\datapath.registers.838[15] [0])
);

DFFPOSX1 _20438_ (
    .CLK(CLK_bF$buf150),
    .D(_3965_),
    .Q(\datapath.registers.838[15] [1])
);

DFFPOSX1 _20439_ (
    .CLK(CLK_bF$buf149),
    .D(_3976_),
    .Q(\datapath.registers.838[15] [2])
);

DFFPOSX1 _20440_ (
    .CLK(CLK_bF$buf148),
    .D(_3979_),
    .Q(\datapath.registers.838[15] [3])
);

DFFPOSX1 _20441_ (
    .CLK(CLK_bF$buf147),
    .D(_3980_),
    .Q(\datapath.registers.838[15] [4])
);

DFFPOSX1 _20442_ (
    .CLK(CLK_bF$buf146),
    .D(_3981_),
    .Q(\datapath.registers.838[15] [5])
);

DFFPOSX1 _20443_ (
    .CLK(CLK_bF$buf145),
    .D(_3982_),
    .Q(\datapath.registers.838[15] [6])
);

DFFPOSX1 _20444_ (
    .CLK(CLK_bF$buf144),
    .D(_3983_),
    .Q(\datapath.registers.838[15] [7])
);

DFFPOSX1 _20445_ (
    .CLK(CLK_bF$buf143),
    .D(_3984_),
    .Q(\datapath.registers.838[15] [8])
);

DFFPOSX1 _20446_ (
    .CLK(CLK_bF$buf142),
    .D(_3985_),
    .Q(\datapath.registers.838[15] [9])
);

DFFPOSX1 _20447_ (
    .CLK(CLK_bF$buf141),
    .D(_3955_),
    .Q(\datapath.registers.838[15] [10])
);

DFFPOSX1 _20448_ (
    .CLK(CLK_bF$buf140),
    .D(_3956_),
    .Q(\datapath.registers.838[15] [11])
);

DFFPOSX1 _20449_ (
    .CLK(CLK_bF$buf139),
    .D(_3957_),
    .Q(\datapath.registers.838[15] [12])
);

DFFPOSX1 _20450_ (
    .CLK(CLK_bF$buf138),
    .D(_3958_),
    .Q(\datapath.registers.838[15] [13])
);

DFFPOSX1 _20451_ (
    .CLK(CLK_bF$buf137),
    .D(_3959_),
    .Q(\datapath.registers.838[15] [14])
);

DFFPOSX1 _20452_ (
    .CLK(CLK_bF$buf136),
    .D(_3960_),
    .Q(\datapath.registers.838[15] [15])
);

DFFPOSX1 _20453_ (
    .CLK(CLK_bF$buf135),
    .D(_3961_),
    .Q(\datapath.registers.838[15] [16])
);

DFFPOSX1 _20454_ (
    .CLK(CLK_bF$buf134),
    .D(_3962_),
    .Q(\datapath.registers.838[15] [17])
);

DFFPOSX1 _20455_ (
    .CLK(CLK_bF$buf133),
    .D(_3963_),
    .Q(\datapath.registers.838[15] [18])
);

DFFPOSX1 _20456_ (
    .CLK(CLK_bF$buf132),
    .D(_3964_),
    .Q(\datapath.registers.838[15] [19])
);

DFFPOSX1 _20457_ (
    .CLK(CLK_bF$buf131),
    .D(_3966_),
    .Q(\datapath.registers.838[15] [20])
);

DFFPOSX1 _20458_ (
    .CLK(CLK_bF$buf130),
    .D(_3967_),
    .Q(\datapath.registers.838[15] [21])
);

DFFPOSX1 _20459_ (
    .CLK(CLK_bF$buf129),
    .D(_3968_),
    .Q(\datapath.registers.838[15] [22])
);

DFFPOSX1 _20460_ (
    .CLK(CLK_bF$buf128),
    .D(_3969_),
    .Q(\datapath.registers.838[15] [23])
);

DFFPOSX1 _20461_ (
    .CLK(CLK_bF$buf127),
    .D(_3970_),
    .Q(\datapath.registers.838[15] [24])
);

DFFPOSX1 _20462_ (
    .CLK(CLK_bF$buf126),
    .D(_3971_),
    .Q(\datapath.registers.838[15] [25])
);

DFFPOSX1 _20463_ (
    .CLK(CLK_bF$buf125),
    .D(_3972_),
    .Q(\datapath.registers.838[15] [26])
);

DFFPOSX1 _20464_ (
    .CLK(CLK_bF$buf124),
    .D(_3973_),
    .Q(\datapath.registers.838[15] [27])
);

DFFPOSX1 _20465_ (
    .CLK(CLK_bF$buf123),
    .D(_3974_),
    .Q(\datapath.registers.838[15] [28])
);

DFFPOSX1 _20466_ (
    .CLK(CLK_bF$buf122),
    .D(_3975_),
    .Q(\datapath.registers.838[15] [29])
);

DFFPOSX1 _20467_ (
    .CLK(CLK_bF$buf121),
    .D(_3977_),
    .Q(\datapath.registers.838[15] [30])
);

DFFPOSX1 _20468_ (
    .CLK(CLK_bF$buf120),
    .D(_3978_),
    .Q(\datapath.registers.838[15] [31])
);

DFFPOSX1 _20469_ (
    .CLK(CLK_bF$buf119),
    .D(_3826_),
    .Q(\datapath.registers.838[11] [0])
);

DFFPOSX1 _20470_ (
    .CLK(CLK_bF$buf118),
    .D(_3837_),
    .Q(\datapath.registers.838[11] [1])
);

DFFPOSX1 _20471_ (
    .CLK(CLK_bF$buf117),
    .D(_3848_),
    .Q(\datapath.registers.838[11] [2])
);

DFFPOSX1 _20472_ (
    .CLK(CLK_bF$buf116),
    .D(_3851_),
    .Q(\datapath.registers.838[11] [3])
);

DFFPOSX1 _20473_ (
    .CLK(CLK_bF$buf115),
    .D(_3852_),
    .Q(\datapath.registers.838[11] [4])
);

DFFPOSX1 _20474_ (
    .CLK(CLK_bF$buf114),
    .D(_3853_),
    .Q(\datapath.registers.838[11] [5])
);

DFFPOSX1 _20475_ (
    .CLK(CLK_bF$buf113),
    .D(_3854_),
    .Q(\datapath.registers.838[11] [6])
);

DFFPOSX1 _20476_ (
    .CLK(CLK_bF$buf112),
    .D(_3855_),
    .Q(\datapath.registers.838[11] [7])
);

DFFPOSX1 _20477_ (
    .CLK(CLK_bF$buf111),
    .D(_3856_),
    .Q(\datapath.registers.838[11] [8])
);

DFFPOSX1 _20478_ (
    .CLK(CLK_bF$buf110),
    .D(_3857_),
    .Q(\datapath.registers.838[11] [9])
);

DFFPOSX1 _20479_ (
    .CLK(CLK_bF$buf109),
    .D(_3827_),
    .Q(\datapath.registers.838[11] [10])
);

DFFPOSX1 _20480_ (
    .CLK(CLK_bF$buf108),
    .D(_3828_),
    .Q(\datapath.registers.838[11] [11])
);

DFFPOSX1 _20481_ (
    .CLK(CLK_bF$buf107),
    .D(_3829_),
    .Q(\datapath.registers.838[11] [12])
);

DFFPOSX1 _20482_ (
    .CLK(CLK_bF$buf106),
    .D(_3830_),
    .Q(\datapath.registers.838[11] [13])
);

DFFPOSX1 _20483_ (
    .CLK(CLK_bF$buf105),
    .D(_3831_),
    .Q(\datapath.registers.838[11] [14])
);

DFFPOSX1 _20484_ (
    .CLK(CLK_bF$buf104),
    .D(_3832_),
    .Q(\datapath.registers.838[11] [15])
);

DFFPOSX1 _20485_ (
    .CLK(CLK_bF$buf103),
    .D(_3833_),
    .Q(\datapath.registers.838[11] [16])
);

DFFPOSX1 _20486_ (
    .CLK(CLK_bF$buf102),
    .D(_3834_),
    .Q(\datapath.registers.838[11] [17])
);

DFFPOSX1 _20487_ (
    .CLK(CLK_bF$buf101),
    .D(_3835_),
    .Q(\datapath.registers.838[11] [18])
);

DFFPOSX1 _20488_ (
    .CLK(CLK_bF$buf100),
    .D(_3836_),
    .Q(\datapath.registers.838[11] [19])
);

DFFPOSX1 _20489_ (
    .CLK(CLK_bF$buf99),
    .D(_3838_),
    .Q(\datapath.registers.838[11] [20])
);

DFFPOSX1 _20490_ (
    .CLK(CLK_bF$buf98),
    .D(_3839_),
    .Q(\datapath.registers.838[11] [21])
);

DFFPOSX1 _20491_ (
    .CLK(CLK_bF$buf97),
    .D(_3840_),
    .Q(\datapath.registers.838[11] [22])
);

DFFPOSX1 _20492_ (
    .CLK(CLK_bF$buf96),
    .D(_3841_),
    .Q(\datapath.registers.838[11] [23])
);

DFFPOSX1 _20493_ (
    .CLK(CLK_bF$buf95),
    .D(_3842_),
    .Q(\datapath.registers.838[11] [24])
);

DFFPOSX1 _20494_ (
    .CLK(CLK_bF$buf94),
    .D(_3843_),
    .Q(\datapath.registers.838[11] [25])
);

DFFPOSX1 _20495_ (
    .CLK(CLK_bF$buf93),
    .D(_3844_),
    .Q(\datapath.registers.838[11] [26])
);

DFFPOSX1 _20496_ (
    .CLK(CLK_bF$buf92),
    .D(_3845_),
    .Q(\datapath.registers.838[11] [27])
);

DFFPOSX1 _20497_ (
    .CLK(CLK_bF$buf91),
    .D(_3846_),
    .Q(\datapath.registers.838[11] [28])
);

DFFPOSX1 _20498_ (
    .CLK(CLK_bF$buf90),
    .D(_3847_),
    .Q(\datapath.registers.838[11] [29])
);

DFFPOSX1 _20499_ (
    .CLK(CLK_bF$buf89),
    .D(_3849_),
    .Q(\datapath.registers.838[11] [30])
);

DFFPOSX1 _20500_ (
    .CLK(CLK_bF$buf88),
    .D(_3850_),
    .Q(\datapath.registers.838[11] [31])
);

DFFPOSX1 _20501_ (
    .CLK(CLK_bF$buf87),
    .D(_3794_),
    .Q(\datapath.registers.838[10] [0])
);

DFFPOSX1 _20502_ (
    .CLK(CLK_bF$buf86),
    .D(_3805_),
    .Q(\datapath.registers.838[10] [1])
);

DFFPOSX1 _20503_ (
    .CLK(CLK_bF$buf85),
    .D(_3816_),
    .Q(\datapath.registers.838[10] [2])
);

DFFPOSX1 _20504_ (
    .CLK(CLK_bF$buf84),
    .D(_3819_),
    .Q(\datapath.registers.838[10] [3])
);

DFFPOSX1 _20505_ (
    .CLK(CLK_bF$buf83),
    .D(_3820_),
    .Q(\datapath.registers.838[10] [4])
);

DFFPOSX1 _20506_ (
    .CLK(CLK_bF$buf82),
    .D(_3821_),
    .Q(\datapath.registers.838[10] [5])
);

DFFPOSX1 _20507_ (
    .CLK(CLK_bF$buf81),
    .D(_3822_),
    .Q(\datapath.registers.838[10] [6])
);

DFFPOSX1 _20508_ (
    .CLK(CLK_bF$buf80),
    .D(_3823_),
    .Q(\datapath.registers.838[10] [7])
);

DFFPOSX1 _20509_ (
    .CLK(CLK_bF$buf79),
    .D(_3824_),
    .Q(\datapath.registers.838[10] [8])
);

DFFPOSX1 _20510_ (
    .CLK(CLK_bF$buf78),
    .D(_3825_),
    .Q(\datapath.registers.838[10] [9])
);

DFFPOSX1 _20511_ (
    .CLK(CLK_bF$buf77),
    .D(_3795_),
    .Q(\datapath.registers.838[10] [10])
);

DFFPOSX1 _20512_ (
    .CLK(CLK_bF$buf76),
    .D(_3796_),
    .Q(\datapath.registers.838[10] [11])
);

DFFPOSX1 _20513_ (
    .CLK(CLK_bF$buf75),
    .D(_3797_),
    .Q(\datapath.registers.838[10] [12])
);

DFFPOSX1 _20514_ (
    .CLK(CLK_bF$buf74),
    .D(_3798_),
    .Q(\datapath.registers.838[10] [13])
);

DFFPOSX1 _20515_ (
    .CLK(CLK_bF$buf73),
    .D(_3799_),
    .Q(\datapath.registers.838[10] [14])
);

DFFPOSX1 _20516_ (
    .CLK(CLK_bF$buf72),
    .D(_3800_),
    .Q(\datapath.registers.838[10] [15])
);

DFFPOSX1 _20517_ (
    .CLK(CLK_bF$buf71),
    .D(_3801_),
    .Q(\datapath.registers.838[10] [16])
);

DFFPOSX1 _20518_ (
    .CLK(CLK_bF$buf70),
    .D(_3802_),
    .Q(\datapath.registers.838[10] [17])
);

DFFPOSX1 _20519_ (
    .CLK(CLK_bF$buf69),
    .D(_3803_),
    .Q(\datapath.registers.838[10] [18])
);

DFFPOSX1 _20520_ (
    .CLK(CLK_bF$buf68),
    .D(_3804_),
    .Q(\datapath.registers.838[10] [19])
);

DFFPOSX1 _20521_ (
    .CLK(CLK_bF$buf67),
    .D(_3806_),
    .Q(\datapath.registers.838[10] [20])
);

DFFPOSX1 _20522_ (
    .CLK(CLK_bF$buf66),
    .D(_3807_),
    .Q(\datapath.registers.838[10] [21])
);

DFFPOSX1 _20523_ (
    .CLK(CLK_bF$buf65),
    .D(_3808_),
    .Q(\datapath.registers.838[10] [22])
);

DFFPOSX1 _20524_ (
    .CLK(CLK_bF$buf64),
    .D(_3809_),
    .Q(\datapath.registers.838[10] [23])
);

DFFPOSX1 _20525_ (
    .CLK(CLK_bF$buf63),
    .D(_3810_),
    .Q(\datapath.registers.838[10] [24])
);

DFFPOSX1 _20526_ (
    .CLK(CLK_bF$buf62),
    .D(_3811_),
    .Q(\datapath.registers.838[10] [25])
);

DFFPOSX1 _20527_ (
    .CLK(CLK_bF$buf61),
    .D(_3812_),
    .Q(\datapath.registers.838[10] [26])
);

DFFPOSX1 _20528_ (
    .CLK(CLK_bF$buf60),
    .D(_3813_),
    .Q(\datapath.registers.838[10] [27])
);

DFFPOSX1 _20529_ (
    .CLK(CLK_bF$buf59),
    .D(_3814_),
    .Q(\datapath.registers.838[10] [28])
);

DFFPOSX1 _20530_ (
    .CLK(CLK_bF$buf58),
    .D(_3815_),
    .Q(\datapath.registers.838[10] [29])
);

DFFPOSX1 _20531_ (
    .CLK(CLK_bF$buf57),
    .D(_3817_),
    .Q(\datapath.registers.838[10] [30])
);

DFFPOSX1 _20532_ (
    .CLK(CLK_bF$buf56),
    .D(_3818_),
    .Q(\datapath.registers.838[10] [31])
);

DFFPOSX1 _20533_ (
    .CLK(CLK_bF$buf55),
    .D(_4722_),
    .Q(\datapath.registers.838[8] [0])
);

DFFPOSX1 _20534_ (
    .CLK(CLK_bF$buf54),
    .D(_4733_),
    .Q(\datapath.registers.838[8] [1])
);

DFFPOSX1 _20535_ (
    .CLK(CLK_bF$buf53),
    .D(_4744_),
    .Q(\datapath.registers.838[8] [2])
);

DFFPOSX1 _20536_ (
    .CLK(CLK_bF$buf52),
    .D(_4747_),
    .Q(\datapath.registers.838[8] [3])
);

DFFPOSX1 _20537_ (
    .CLK(CLK_bF$buf51),
    .D(_4748_),
    .Q(\datapath.registers.838[8] [4])
);

DFFPOSX1 _20538_ (
    .CLK(CLK_bF$buf50),
    .D(_4749_),
    .Q(\datapath.registers.838[8] [5])
);

DFFPOSX1 _20539_ (
    .CLK(CLK_bF$buf49),
    .D(_4750_),
    .Q(\datapath.registers.838[8] [6])
);

DFFPOSX1 _20540_ (
    .CLK(CLK_bF$buf48),
    .D(_4751_),
    .Q(\datapath.registers.838[8] [7])
);

DFFPOSX1 _20541_ (
    .CLK(CLK_bF$buf47),
    .D(_4752_),
    .Q(\datapath.registers.838[8] [8])
);

DFFPOSX1 _20542_ (
    .CLK(CLK_bF$buf46),
    .D(_4753_),
    .Q(\datapath.registers.838[8] [9])
);

DFFPOSX1 _20543_ (
    .CLK(CLK_bF$buf45),
    .D(_4723_),
    .Q(\datapath.registers.838[8] [10])
);

DFFPOSX1 _20544_ (
    .CLK(CLK_bF$buf44),
    .D(_4724_),
    .Q(\datapath.registers.838[8] [11])
);

DFFPOSX1 _20545_ (
    .CLK(CLK_bF$buf43),
    .D(_4725_),
    .Q(\datapath.registers.838[8] [12])
);

DFFPOSX1 _20546_ (
    .CLK(CLK_bF$buf42),
    .D(_4726_),
    .Q(\datapath.registers.838[8] [13])
);

DFFPOSX1 _20547_ (
    .CLK(CLK_bF$buf41),
    .D(_4727_),
    .Q(\datapath.registers.838[8] [14])
);

DFFPOSX1 _20548_ (
    .CLK(CLK_bF$buf40),
    .D(_4728_),
    .Q(\datapath.registers.838[8] [15])
);

DFFPOSX1 _20549_ (
    .CLK(CLK_bF$buf39),
    .D(_4729_),
    .Q(\datapath.registers.838[8] [16])
);

DFFPOSX1 _20550_ (
    .CLK(CLK_bF$buf38),
    .D(_4730_),
    .Q(\datapath.registers.838[8] [17])
);

DFFPOSX1 _20551_ (
    .CLK(CLK_bF$buf37),
    .D(_4731_),
    .Q(\datapath.registers.838[8] [18])
);

DFFPOSX1 _20552_ (
    .CLK(CLK_bF$buf36),
    .D(_4732_),
    .Q(\datapath.registers.838[8] [19])
);

DFFPOSX1 _20553_ (
    .CLK(CLK_bF$buf35),
    .D(_4734_),
    .Q(\datapath.registers.838[8] [20])
);

DFFPOSX1 _20554_ (
    .CLK(CLK_bF$buf34),
    .D(_4735_),
    .Q(\datapath.registers.838[8] [21])
);

DFFPOSX1 _20555_ (
    .CLK(CLK_bF$buf33),
    .D(_4736_),
    .Q(\datapath.registers.838[8] [22])
);

DFFPOSX1 _20556_ (
    .CLK(CLK_bF$buf32),
    .D(_4737_),
    .Q(\datapath.registers.838[8] [23])
);

DFFPOSX1 _20557_ (
    .CLK(CLK_bF$buf31),
    .D(_4738_),
    .Q(\datapath.registers.838[8] [24])
);

DFFPOSX1 _20558_ (
    .CLK(CLK_bF$buf30),
    .D(_4739_),
    .Q(\datapath.registers.838[8] [25])
);

DFFPOSX1 _20559_ (
    .CLK(CLK_bF$buf29),
    .D(_4740_),
    .Q(\datapath.registers.838[8] [26])
);

DFFPOSX1 _20560_ (
    .CLK(CLK_bF$buf28),
    .D(_4741_),
    .Q(\datapath.registers.838[8] [27])
);

DFFPOSX1 _20561_ (
    .CLK(CLK_bF$buf27),
    .D(_4742_),
    .Q(\datapath.registers.838[8] [28])
);

DFFPOSX1 _20562_ (
    .CLK(CLK_bF$buf26),
    .D(_4743_),
    .Q(\datapath.registers.838[8] [29])
);

DFFPOSX1 _20563_ (
    .CLK(CLK_bF$buf25),
    .D(_4745_),
    .Q(\datapath.registers.838[8] [30])
);

DFFPOSX1 _20564_ (
    .CLK(CLK_bF$buf24),
    .D(_4746_),
    .Q(\datapath.registers.838[8] [31])
);

DFFPOSX1 _20565_ (
    .CLK(CLK_bF$buf23),
    .D(_4658_),
    .Q(\datapath.registers.838[6] [0])
);

DFFPOSX1 _20566_ (
    .CLK(CLK_bF$buf22),
    .D(_4669_),
    .Q(\datapath.registers.838[6] [1])
);

DFFPOSX1 _20567_ (
    .CLK(CLK_bF$buf21),
    .D(_4680_),
    .Q(\datapath.registers.838[6] [2])
);

DFFPOSX1 _20568_ (
    .CLK(CLK_bF$buf20),
    .D(_4683_),
    .Q(\datapath.registers.838[6] [3])
);

DFFPOSX1 _20569_ (
    .CLK(CLK_bF$buf19),
    .D(_4684_),
    .Q(\datapath.registers.838[6] [4])
);

DFFPOSX1 _20570_ (
    .CLK(CLK_bF$buf18),
    .D(_4685_),
    .Q(\datapath.registers.838[6] [5])
);

DFFPOSX1 _20571_ (
    .CLK(CLK_bF$buf17),
    .D(_4686_),
    .Q(\datapath.registers.838[6] [6])
);

DFFPOSX1 _20572_ (
    .CLK(CLK_bF$buf16),
    .D(_4687_),
    .Q(\datapath.registers.838[6] [7])
);

DFFPOSX1 _20573_ (
    .CLK(CLK_bF$buf15),
    .D(_4688_),
    .Q(\datapath.registers.838[6] [8])
);

DFFPOSX1 _20574_ (
    .CLK(CLK_bF$buf14),
    .D(_4689_),
    .Q(\datapath.registers.838[6] [9])
);

DFFPOSX1 _20575_ (
    .CLK(CLK_bF$buf13),
    .D(_4659_),
    .Q(\datapath.registers.838[6] [10])
);

DFFPOSX1 _20576_ (
    .CLK(CLK_bF$buf12),
    .D(_4660_),
    .Q(\datapath.registers.838[6] [11])
);

DFFPOSX1 _20577_ (
    .CLK(CLK_bF$buf11),
    .D(_4661_),
    .Q(\datapath.registers.838[6] [12])
);

DFFPOSX1 _20578_ (
    .CLK(CLK_bF$buf10),
    .D(_4662_),
    .Q(\datapath.registers.838[6] [13])
);

DFFPOSX1 _20579_ (
    .CLK(CLK_bF$buf9),
    .D(_4663_),
    .Q(\datapath.registers.838[6] [14])
);

DFFPOSX1 _20580_ (
    .CLK(CLK_bF$buf8),
    .D(_4664_),
    .Q(\datapath.registers.838[6] [15])
);

DFFPOSX1 _20581_ (
    .CLK(CLK_bF$buf7),
    .D(_4665_),
    .Q(\datapath.registers.838[6] [16])
);

DFFPOSX1 _20582_ (
    .CLK(CLK_bF$buf6),
    .D(_4666_),
    .Q(\datapath.registers.838[6] [17])
);

DFFPOSX1 _20583_ (
    .CLK(CLK_bF$buf5),
    .D(_4667_),
    .Q(\datapath.registers.838[6] [18])
);

DFFPOSX1 _20584_ (
    .CLK(CLK_bF$buf4),
    .D(_4668_),
    .Q(\datapath.registers.838[6] [19])
);

DFFPOSX1 _20585_ (
    .CLK(CLK_bF$buf3),
    .D(_4670_),
    .Q(\datapath.registers.838[6] [20])
);

DFFPOSX1 _20586_ (
    .CLK(CLK_bF$buf2),
    .D(_4671_),
    .Q(\datapath.registers.838[6] [21])
);

DFFPOSX1 _20587_ (
    .CLK(CLK_bF$buf1),
    .D(_4672_),
    .Q(\datapath.registers.838[6] [22])
);

DFFPOSX1 _20588_ (
    .CLK(CLK_bF$buf0),
    .D(_4673_),
    .Q(\datapath.registers.838[6] [23])
);

DFFPOSX1 _20589_ (
    .CLK(CLK_bF$buf151),
    .D(_4674_),
    .Q(\datapath.registers.838[6] [24])
);

DFFPOSX1 _20590_ (
    .CLK(CLK_bF$buf150),
    .D(_4675_),
    .Q(\datapath.registers.838[6] [25])
);

DFFPOSX1 _20591_ (
    .CLK(CLK_bF$buf149),
    .D(_4676_),
    .Q(\datapath.registers.838[6] [26])
);

DFFPOSX1 _20592_ (
    .CLK(CLK_bF$buf148),
    .D(_4677_),
    .Q(\datapath.registers.838[6] [27])
);

DFFPOSX1 _20593_ (
    .CLK(CLK_bF$buf147),
    .D(_4678_),
    .Q(\datapath.registers.838[6] [28])
);

DFFPOSX1 _20594_ (
    .CLK(CLK_bF$buf146),
    .D(_4679_),
    .Q(\datapath.registers.838[6] [29])
);

DFFPOSX1 _20595_ (
    .CLK(CLK_bF$buf145),
    .D(_4681_),
    .Q(\datapath.registers.838[6] [30])
);

DFFPOSX1 _20596_ (
    .CLK(CLK_bF$buf144),
    .D(_4682_),
    .Q(\datapath.registers.838[6] [31])
);

DFFPOSX1 _20597_ (
    .CLK(CLK_bF$buf143),
    .D(_4146_),
    .Q(\datapath.registers.838[20] [0])
);

DFFPOSX1 _20598_ (
    .CLK(CLK_bF$buf142),
    .D(_4157_),
    .Q(\datapath.registers.838[20] [1])
);

DFFPOSX1 _20599_ (
    .CLK(CLK_bF$buf141),
    .D(_4168_),
    .Q(\datapath.registers.838[20] [2])
);

DFFPOSX1 _20600_ (
    .CLK(CLK_bF$buf140),
    .D(_4171_),
    .Q(\datapath.registers.838[20] [3])
);

DFFPOSX1 _20601_ (
    .CLK(CLK_bF$buf139),
    .D(_4172_),
    .Q(\datapath.registers.838[20] [4])
);

DFFPOSX1 _20602_ (
    .CLK(CLK_bF$buf138),
    .D(_4173_),
    .Q(\datapath.registers.838[20] [5])
);

DFFPOSX1 _20603_ (
    .CLK(CLK_bF$buf137),
    .D(_4174_),
    .Q(\datapath.registers.838[20] [6])
);

DFFPOSX1 _20604_ (
    .CLK(CLK_bF$buf136),
    .D(_4175_),
    .Q(\datapath.registers.838[20] [7])
);

DFFPOSX1 _20605_ (
    .CLK(CLK_bF$buf135),
    .D(_4176_),
    .Q(\datapath.registers.838[20] [8])
);

DFFPOSX1 _20606_ (
    .CLK(CLK_bF$buf134),
    .D(_4177_),
    .Q(\datapath.registers.838[20] [9])
);

DFFPOSX1 _20607_ (
    .CLK(CLK_bF$buf133),
    .D(_4147_),
    .Q(\datapath.registers.838[20] [10])
);

DFFPOSX1 _20608_ (
    .CLK(CLK_bF$buf132),
    .D(_4148_),
    .Q(\datapath.registers.838[20] [11])
);

DFFPOSX1 _20609_ (
    .CLK(CLK_bF$buf131),
    .D(_4149_),
    .Q(\datapath.registers.838[20] [12])
);

DFFPOSX1 _20610_ (
    .CLK(CLK_bF$buf130),
    .D(_4150_),
    .Q(\datapath.registers.838[20] [13])
);

DFFPOSX1 _20611_ (
    .CLK(CLK_bF$buf129),
    .D(_4151_),
    .Q(\datapath.registers.838[20] [14])
);

DFFPOSX1 _20612_ (
    .CLK(CLK_bF$buf128),
    .D(_4152_),
    .Q(\datapath.registers.838[20] [15])
);

DFFPOSX1 _20613_ (
    .CLK(CLK_bF$buf127),
    .D(_4153_),
    .Q(\datapath.registers.838[20] [16])
);

DFFPOSX1 _20614_ (
    .CLK(CLK_bF$buf126),
    .D(_4154_),
    .Q(\datapath.registers.838[20] [17])
);

DFFPOSX1 _20615_ (
    .CLK(CLK_bF$buf125),
    .D(_4155_),
    .Q(\datapath.registers.838[20] [18])
);

DFFPOSX1 _20616_ (
    .CLK(CLK_bF$buf124),
    .D(_4156_),
    .Q(\datapath.registers.838[20] [19])
);

DFFPOSX1 _20617_ (
    .CLK(CLK_bF$buf123),
    .D(_4158_),
    .Q(\datapath.registers.838[20] [20])
);

DFFPOSX1 _20618_ (
    .CLK(CLK_bF$buf122),
    .D(_4159_),
    .Q(\datapath.registers.838[20] [21])
);

DFFPOSX1 _20619_ (
    .CLK(CLK_bF$buf121),
    .D(_4160_),
    .Q(\datapath.registers.838[20] [22])
);

DFFPOSX1 _20620_ (
    .CLK(CLK_bF$buf120),
    .D(_4161_),
    .Q(\datapath.registers.838[20] [23])
);

DFFPOSX1 _20621_ (
    .CLK(CLK_bF$buf119),
    .D(_4162_),
    .Q(\datapath.registers.838[20] [24])
);

DFFPOSX1 _20622_ (
    .CLK(CLK_bF$buf118),
    .D(_4163_),
    .Q(\datapath.registers.838[20] [25])
);

DFFPOSX1 _20623_ (
    .CLK(CLK_bF$buf117),
    .D(_4164_),
    .Q(\datapath.registers.838[20] [26])
);

DFFPOSX1 _20624_ (
    .CLK(CLK_bF$buf116),
    .D(_4165_),
    .Q(\datapath.registers.838[20] [27])
);

DFFPOSX1 _20625_ (
    .CLK(CLK_bF$buf115),
    .D(_4166_),
    .Q(\datapath.registers.838[20] [28])
);

DFFPOSX1 _20626_ (
    .CLK(CLK_bF$buf114),
    .D(_4167_),
    .Q(\datapath.registers.838[20] [29])
);

DFFPOSX1 _20627_ (
    .CLK(CLK_bF$buf113),
    .D(_4169_),
    .Q(\datapath.registers.838[20] [30])
);

DFFPOSX1 _20628_ (
    .CLK(CLK_bF$buf112),
    .D(_4170_),
    .Q(\datapath.registers.838[20] [31])
);

DFFPOSX1 _20629_ (
    .CLK(CLK_bF$buf111),
    .D(_4242_),
    .Q(\datapath.registers.838[23] [0])
);

DFFPOSX1 _20630_ (
    .CLK(CLK_bF$buf110),
    .D(_4253_),
    .Q(\datapath.registers.838[23] [1])
);

DFFPOSX1 _20631_ (
    .CLK(CLK_bF$buf109),
    .D(_4264_),
    .Q(\datapath.registers.838[23] [2])
);

DFFPOSX1 _20632_ (
    .CLK(CLK_bF$buf108),
    .D(_4267_),
    .Q(\datapath.registers.838[23] [3])
);

DFFPOSX1 _20633_ (
    .CLK(CLK_bF$buf107),
    .D(_4268_),
    .Q(\datapath.registers.838[23] [4])
);

DFFPOSX1 _20634_ (
    .CLK(CLK_bF$buf106),
    .D(_4269_),
    .Q(\datapath.registers.838[23] [5])
);

DFFPOSX1 _20635_ (
    .CLK(CLK_bF$buf105),
    .D(_4270_),
    .Q(\datapath.registers.838[23] [6])
);

DFFPOSX1 _20636_ (
    .CLK(CLK_bF$buf104),
    .D(_4271_),
    .Q(\datapath.registers.838[23] [7])
);

DFFPOSX1 _20637_ (
    .CLK(CLK_bF$buf103),
    .D(_4272_),
    .Q(\datapath.registers.838[23] [8])
);

DFFPOSX1 _20638_ (
    .CLK(CLK_bF$buf102),
    .D(_4273_),
    .Q(\datapath.registers.838[23] [9])
);

DFFPOSX1 _20639_ (
    .CLK(CLK_bF$buf101),
    .D(_4243_),
    .Q(\datapath.registers.838[23] [10])
);

DFFPOSX1 _20640_ (
    .CLK(CLK_bF$buf100),
    .D(_4244_),
    .Q(\datapath.registers.838[23] [11])
);

DFFPOSX1 _20641_ (
    .CLK(CLK_bF$buf99),
    .D(_4245_),
    .Q(\datapath.registers.838[23] [12])
);

DFFPOSX1 _20642_ (
    .CLK(CLK_bF$buf98),
    .D(_4246_),
    .Q(\datapath.registers.838[23] [13])
);

DFFPOSX1 _20643_ (
    .CLK(CLK_bF$buf97),
    .D(_4247_),
    .Q(\datapath.registers.838[23] [14])
);

DFFPOSX1 _20644_ (
    .CLK(CLK_bF$buf96),
    .D(_4248_),
    .Q(\datapath.registers.838[23] [15])
);

DFFPOSX1 _20645_ (
    .CLK(CLK_bF$buf95),
    .D(_4249_),
    .Q(\datapath.registers.838[23] [16])
);

DFFPOSX1 _20646_ (
    .CLK(CLK_bF$buf94),
    .D(_4250_),
    .Q(\datapath.registers.838[23] [17])
);

DFFPOSX1 _20647_ (
    .CLK(CLK_bF$buf93),
    .D(_4251_),
    .Q(\datapath.registers.838[23] [18])
);

DFFPOSX1 _20648_ (
    .CLK(CLK_bF$buf92),
    .D(_4252_),
    .Q(\datapath.registers.838[23] [19])
);

DFFPOSX1 _20649_ (
    .CLK(CLK_bF$buf91),
    .D(_4254_),
    .Q(\datapath.registers.838[23] [20])
);

DFFPOSX1 _20650_ (
    .CLK(CLK_bF$buf90),
    .D(_4255_),
    .Q(\datapath.registers.838[23] [21])
);

DFFPOSX1 _20651_ (
    .CLK(CLK_bF$buf89),
    .D(_4256_),
    .Q(\datapath.registers.838[23] [22])
);

DFFPOSX1 _20652_ (
    .CLK(CLK_bF$buf88),
    .D(_4257_),
    .Q(\datapath.registers.838[23] [23])
);

DFFPOSX1 _20653_ (
    .CLK(CLK_bF$buf87),
    .D(_4258_),
    .Q(\datapath.registers.838[23] [24])
);

DFFPOSX1 _20654_ (
    .CLK(CLK_bF$buf86),
    .D(_4259_),
    .Q(\datapath.registers.838[23] [25])
);

DFFPOSX1 _20655_ (
    .CLK(CLK_bF$buf85),
    .D(_4260_),
    .Q(\datapath.registers.838[23] [26])
);

DFFPOSX1 _20656_ (
    .CLK(CLK_bF$buf84),
    .D(_4261_),
    .Q(\datapath.registers.838[23] [27])
);

DFFPOSX1 _20657_ (
    .CLK(CLK_bF$buf83),
    .D(_4262_),
    .Q(\datapath.registers.838[23] [28])
);

DFFPOSX1 _20658_ (
    .CLK(CLK_bF$buf82),
    .D(_4263_),
    .Q(\datapath.registers.838[23] [29])
);

DFFPOSX1 _20659_ (
    .CLK(CLK_bF$buf81),
    .D(_4265_),
    .Q(\datapath.registers.838[23] [30])
);

DFFPOSX1 _20660_ (
    .CLK(CLK_bF$buf80),
    .D(_4266_),
    .Q(\datapath.registers.838[23] [31])
);

DFFPOSX1 _20661_ (
    .CLK(CLK_bF$buf79),
    .D(_3922_),
    .Q(\datapath.registers.838[14] [0])
);

DFFPOSX1 _20662_ (
    .CLK(CLK_bF$buf78),
    .D(_3933_),
    .Q(\datapath.registers.838[14] [1])
);

DFFPOSX1 _20663_ (
    .CLK(CLK_bF$buf77),
    .D(_3944_),
    .Q(\datapath.registers.838[14] [2])
);

DFFPOSX1 _20664_ (
    .CLK(CLK_bF$buf76),
    .D(_3947_),
    .Q(\datapath.registers.838[14] [3])
);

DFFPOSX1 _20665_ (
    .CLK(CLK_bF$buf75),
    .D(_3948_),
    .Q(\datapath.registers.838[14] [4])
);

DFFPOSX1 _20666_ (
    .CLK(CLK_bF$buf74),
    .D(_3949_),
    .Q(\datapath.registers.838[14] [5])
);

DFFPOSX1 _20667_ (
    .CLK(CLK_bF$buf73),
    .D(_3950_),
    .Q(\datapath.registers.838[14] [6])
);

DFFPOSX1 _20668_ (
    .CLK(CLK_bF$buf72),
    .D(_3951_),
    .Q(\datapath.registers.838[14] [7])
);

DFFPOSX1 _20669_ (
    .CLK(CLK_bF$buf71),
    .D(_3952_),
    .Q(\datapath.registers.838[14] [8])
);

DFFPOSX1 _20670_ (
    .CLK(CLK_bF$buf70),
    .D(_3953_),
    .Q(\datapath.registers.838[14] [9])
);

DFFPOSX1 _20671_ (
    .CLK(CLK_bF$buf69),
    .D(_3923_),
    .Q(\datapath.registers.838[14] [10])
);

DFFPOSX1 _20672_ (
    .CLK(CLK_bF$buf68),
    .D(_3924_),
    .Q(\datapath.registers.838[14] [11])
);

DFFPOSX1 _20673_ (
    .CLK(CLK_bF$buf67),
    .D(_3925_),
    .Q(\datapath.registers.838[14] [12])
);

DFFPOSX1 _20674_ (
    .CLK(CLK_bF$buf66),
    .D(_3926_),
    .Q(\datapath.registers.838[14] [13])
);

DFFPOSX1 _20675_ (
    .CLK(CLK_bF$buf65),
    .D(_3927_),
    .Q(\datapath.registers.838[14] [14])
);

DFFPOSX1 _20676_ (
    .CLK(CLK_bF$buf64),
    .D(_3928_),
    .Q(\datapath.registers.838[14] [15])
);

DFFPOSX1 _20677_ (
    .CLK(CLK_bF$buf63),
    .D(_3929_),
    .Q(\datapath.registers.838[14] [16])
);

DFFPOSX1 _20678_ (
    .CLK(CLK_bF$buf62),
    .D(_3930_),
    .Q(\datapath.registers.838[14] [17])
);

DFFPOSX1 _20679_ (
    .CLK(CLK_bF$buf61),
    .D(_3931_),
    .Q(\datapath.registers.838[14] [18])
);

DFFPOSX1 _20680_ (
    .CLK(CLK_bF$buf60),
    .D(_3932_),
    .Q(\datapath.registers.838[14] [19])
);

DFFPOSX1 _20681_ (
    .CLK(CLK_bF$buf59),
    .D(_3934_),
    .Q(\datapath.registers.838[14] [20])
);

DFFPOSX1 _20682_ (
    .CLK(CLK_bF$buf58),
    .D(_3935_),
    .Q(\datapath.registers.838[14] [21])
);

DFFPOSX1 _20683_ (
    .CLK(CLK_bF$buf57),
    .D(_3936_),
    .Q(\datapath.registers.838[14] [22])
);

DFFPOSX1 _20684_ (
    .CLK(CLK_bF$buf56),
    .D(_3937_),
    .Q(\datapath.registers.838[14] [23])
);

DFFPOSX1 _20685_ (
    .CLK(CLK_bF$buf55),
    .D(_3938_),
    .Q(\datapath.registers.838[14] [24])
);

DFFPOSX1 _20686_ (
    .CLK(CLK_bF$buf54),
    .D(_3939_),
    .Q(\datapath.registers.838[14] [25])
);

DFFPOSX1 _20687_ (
    .CLK(CLK_bF$buf53),
    .D(_3940_),
    .Q(\datapath.registers.838[14] [26])
);

DFFPOSX1 _20688_ (
    .CLK(CLK_bF$buf52),
    .D(_3941_),
    .Q(\datapath.registers.838[14] [27])
);

DFFPOSX1 _20689_ (
    .CLK(CLK_bF$buf51),
    .D(_3942_),
    .Q(\datapath.registers.838[14] [28])
);

DFFPOSX1 _20690_ (
    .CLK(CLK_bF$buf50),
    .D(_3943_),
    .Q(\datapath.registers.838[14] [29])
);

DFFPOSX1 _20691_ (
    .CLK(CLK_bF$buf49),
    .D(_3945_),
    .Q(\datapath.registers.838[14] [30])
);

DFFPOSX1 _20692_ (
    .CLK(CLK_bF$buf48),
    .D(_3946_),
    .Q(\datapath.registers.838[14] [31])
);

DFFPOSX1 _20693_ (
    .CLK(CLK_bF$buf47),
    .D(_4754_),
    .Q(\datapath.registers.838[9] [0])
);

DFFPOSX1 _20694_ (
    .CLK(CLK_bF$buf46),
    .D(_4765_),
    .Q(\datapath.registers.838[9] [1])
);

DFFPOSX1 _20695_ (
    .CLK(CLK_bF$buf45),
    .D(_4776_),
    .Q(\datapath.registers.838[9] [2])
);

DFFPOSX1 _20696_ (
    .CLK(CLK_bF$buf44),
    .D(_4779_),
    .Q(\datapath.registers.838[9] [3])
);

DFFPOSX1 _20697_ (
    .CLK(CLK_bF$buf43),
    .D(_4780_),
    .Q(\datapath.registers.838[9] [4])
);

DFFPOSX1 _20698_ (
    .CLK(CLK_bF$buf42),
    .D(_4781_),
    .Q(\datapath.registers.838[9] [5])
);

DFFPOSX1 _20699_ (
    .CLK(CLK_bF$buf41),
    .D(_4782_),
    .Q(\datapath.registers.838[9] [6])
);

DFFPOSX1 _20700_ (
    .CLK(CLK_bF$buf40),
    .D(_4783_),
    .Q(\datapath.registers.838[9] [7])
);

DFFPOSX1 _20701_ (
    .CLK(CLK_bF$buf39),
    .D(_4784_),
    .Q(\datapath.registers.838[9] [8])
);

DFFPOSX1 _20702_ (
    .CLK(CLK_bF$buf38),
    .D(_4785_),
    .Q(\datapath.registers.838[9] [9])
);

DFFPOSX1 _20703_ (
    .CLK(CLK_bF$buf37),
    .D(_4755_),
    .Q(\datapath.registers.838[9] [10])
);

DFFPOSX1 _20704_ (
    .CLK(CLK_bF$buf36),
    .D(_4756_),
    .Q(\datapath.registers.838[9] [11])
);

DFFPOSX1 _20705_ (
    .CLK(CLK_bF$buf35),
    .D(_4757_),
    .Q(\datapath.registers.838[9] [12])
);

DFFPOSX1 _20706_ (
    .CLK(CLK_bF$buf34),
    .D(_4758_),
    .Q(\datapath.registers.838[9] [13])
);

DFFPOSX1 _20707_ (
    .CLK(CLK_bF$buf33),
    .D(_4759_),
    .Q(\datapath.registers.838[9] [14])
);

DFFPOSX1 _20708_ (
    .CLK(CLK_bF$buf32),
    .D(_4760_),
    .Q(\datapath.registers.838[9] [15])
);

DFFPOSX1 _20709_ (
    .CLK(CLK_bF$buf31),
    .D(_4761_),
    .Q(\datapath.registers.838[9] [16])
);

DFFPOSX1 _20710_ (
    .CLK(CLK_bF$buf30),
    .D(_4762_),
    .Q(\datapath.registers.838[9] [17])
);

DFFPOSX1 _20711_ (
    .CLK(CLK_bF$buf29),
    .D(_4763_),
    .Q(\datapath.registers.838[9] [18])
);

DFFPOSX1 _20712_ (
    .CLK(CLK_bF$buf28),
    .D(_4764_),
    .Q(\datapath.registers.838[9] [19])
);

DFFPOSX1 _20713_ (
    .CLK(CLK_bF$buf27),
    .D(_4766_),
    .Q(\datapath.registers.838[9] [20])
);

DFFPOSX1 _20714_ (
    .CLK(CLK_bF$buf26),
    .D(_4767_),
    .Q(\datapath.registers.838[9] [21])
);

DFFPOSX1 _20715_ (
    .CLK(CLK_bF$buf25),
    .D(_4768_),
    .Q(\datapath.registers.838[9] [22])
);

DFFPOSX1 _20716_ (
    .CLK(CLK_bF$buf24),
    .D(_4769_),
    .Q(\datapath.registers.838[9] [23])
);

DFFPOSX1 _20717_ (
    .CLK(CLK_bF$buf23),
    .D(_4770_),
    .Q(\datapath.registers.838[9] [24])
);

DFFPOSX1 _20718_ (
    .CLK(CLK_bF$buf22),
    .D(_4771_),
    .Q(\datapath.registers.838[9] [25])
);

DFFPOSX1 _20719_ (
    .CLK(CLK_bF$buf21),
    .D(_4772_),
    .Q(\datapath.registers.838[9] [26])
);

DFFPOSX1 _20720_ (
    .CLK(CLK_bF$buf20),
    .D(_4773_),
    .Q(\datapath.registers.838[9] [27])
);

DFFPOSX1 _20721_ (
    .CLK(CLK_bF$buf19),
    .D(_4774_),
    .Q(\datapath.registers.838[9] [28])
);

DFFPOSX1 _20722_ (
    .CLK(CLK_bF$buf18),
    .D(_4775_),
    .Q(\datapath.registers.838[9] [29])
);

DFFPOSX1 _20723_ (
    .CLK(CLK_bF$buf17),
    .D(_4777_),
    .Q(\datapath.registers.838[9] [30])
);

DFFPOSX1 _20724_ (
    .CLK(CLK_bF$buf16),
    .D(_4778_),
    .Q(\datapath.registers.838[9] [31])
);

DFFPOSX1 _20725_ (
    .CLK(CLK_bF$buf15),
    .D(_3762_),
    .Q(\datapath.registers.838[0] [0])
);

DFFPOSX1 _20726_ (
    .CLK(CLK_bF$buf14),
    .D(_3773_),
    .Q(\datapath.registers.838[0] [1])
);

DFFPOSX1 _20727_ (
    .CLK(CLK_bF$buf13),
    .D(_3784_),
    .Q(\datapath.registers.838[0] [2])
);

DFFPOSX1 _20728_ (
    .CLK(CLK_bF$buf12),
    .D(_3787_),
    .Q(\datapath.registers.838[0] [3])
);

DFFPOSX1 _20729_ (
    .CLK(CLK_bF$buf11),
    .D(_3788_),
    .Q(\datapath.registers.838[0] [4])
);

DFFPOSX1 _20730_ (
    .CLK(CLK_bF$buf10),
    .D(_3789_),
    .Q(\datapath.registers.838[0] [5])
);

DFFPOSX1 _20731_ (
    .CLK(CLK_bF$buf9),
    .D(_3790_),
    .Q(\datapath.registers.838[0] [6])
);

DFFPOSX1 _20732_ (
    .CLK(CLK_bF$buf8),
    .D(_3791_),
    .Q(\datapath.registers.838[0] [7])
);

DFFPOSX1 _20733_ (
    .CLK(CLK_bF$buf7),
    .D(_3792_),
    .Q(\datapath.registers.838[0] [8])
);

DFFPOSX1 _20734_ (
    .CLK(CLK_bF$buf6),
    .D(_3793_),
    .Q(\datapath.registers.838[0] [9])
);

DFFPOSX1 _20735_ (
    .CLK(CLK_bF$buf5),
    .D(_3763_),
    .Q(\datapath.registers.838[0] [10])
);

DFFPOSX1 _20736_ (
    .CLK(CLK_bF$buf4),
    .D(_3764_),
    .Q(\datapath.registers.838[0] [11])
);

DFFPOSX1 _20737_ (
    .CLK(CLK_bF$buf3),
    .D(_3765_),
    .Q(\datapath.registers.838[0] [12])
);

DFFPOSX1 _20738_ (
    .CLK(CLK_bF$buf2),
    .D(_3766_),
    .Q(\datapath.registers.838[0] [13])
);

DFFPOSX1 _20739_ (
    .CLK(CLK_bF$buf1),
    .D(_3767_),
    .Q(\datapath.registers.838[0] [14])
);

DFFPOSX1 _20740_ (
    .CLK(CLK_bF$buf0),
    .D(_3768_),
    .Q(\datapath.registers.838[0] [15])
);

DFFPOSX1 _20741_ (
    .CLK(CLK_bF$buf151),
    .D(_3769_),
    .Q(\datapath.registers.838[0] [16])
);

DFFPOSX1 _20742_ (
    .CLK(CLK_bF$buf150),
    .D(_3770_),
    .Q(\datapath.registers.838[0] [17])
);

DFFPOSX1 _20743_ (
    .CLK(CLK_bF$buf149),
    .D(_3771_),
    .Q(\datapath.registers.838[0] [18])
);

DFFPOSX1 _20744_ (
    .CLK(CLK_bF$buf148),
    .D(_3772_),
    .Q(\datapath.registers.838[0] [19])
);

DFFPOSX1 _20745_ (
    .CLK(CLK_bF$buf147),
    .D(_3774_),
    .Q(\datapath.registers.838[0] [20])
);

DFFPOSX1 _20746_ (
    .CLK(CLK_bF$buf146),
    .D(_3775_),
    .Q(\datapath.registers.838[0] [21])
);

DFFPOSX1 _20747_ (
    .CLK(CLK_bF$buf145),
    .D(_3776_),
    .Q(\datapath.registers.838[0] [22])
);

DFFPOSX1 _20748_ (
    .CLK(CLK_bF$buf144),
    .D(_3777_),
    .Q(\datapath.registers.838[0] [23])
);

DFFPOSX1 _20749_ (
    .CLK(CLK_bF$buf143),
    .D(_3778_),
    .Q(\datapath.registers.838[0] [24])
);

DFFPOSX1 _20750_ (
    .CLK(CLK_bF$buf142),
    .D(_3779_),
    .Q(\datapath.registers.838[0] [25])
);

DFFPOSX1 _20751_ (
    .CLK(CLK_bF$buf141),
    .D(_3780_),
    .Q(\datapath.registers.838[0] [26])
);

DFFPOSX1 _20752_ (
    .CLK(CLK_bF$buf140),
    .D(_3781_),
    .Q(\datapath.registers.838[0] [27])
);

DFFPOSX1 _20753_ (
    .CLK(CLK_bF$buf139),
    .D(_3782_),
    .Q(\datapath.registers.838[0] [28])
);

DFFPOSX1 _20754_ (
    .CLK(CLK_bF$buf138),
    .D(_3783_),
    .Q(\datapath.registers.838[0] [29])
);

DFFPOSX1 _20755_ (
    .CLK(CLK_bF$buf137),
    .D(_3785_),
    .Q(\datapath.registers.838[0] [30])
);

DFFPOSX1 _20756_ (
    .CLK(CLK_bF$buf136),
    .D(_3786_),
    .Q(\datapath.registers.838[0] [31])
);

DFFPOSX1 _20757_ (
    .CLK(CLK_bF$buf135),
    .D(_4626_),
    .Q(\datapath.registers.838[5] [0])
);

DFFPOSX1 _20758_ (
    .CLK(CLK_bF$buf134),
    .D(_4637_),
    .Q(\datapath.registers.838[5] [1])
);

DFFPOSX1 _20759_ (
    .CLK(CLK_bF$buf133),
    .D(_4648_),
    .Q(\datapath.registers.838[5] [2])
);

DFFPOSX1 _20760_ (
    .CLK(CLK_bF$buf132),
    .D(_4651_),
    .Q(\datapath.registers.838[5] [3])
);

DFFPOSX1 _20761_ (
    .CLK(CLK_bF$buf131),
    .D(_4652_),
    .Q(\datapath.registers.838[5] [4])
);

DFFPOSX1 _20762_ (
    .CLK(CLK_bF$buf130),
    .D(_4653_),
    .Q(\datapath.registers.838[5] [5])
);

DFFPOSX1 _20763_ (
    .CLK(CLK_bF$buf129),
    .D(_4654_),
    .Q(\datapath.registers.838[5] [6])
);

DFFPOSX1 _20764_ (
    .CLK(CLK_bF$buf128),
    .D(_4655_),
    .Q(\datapath.registers.838[5] [7])
);

DFFPOSX1 _20765_ (
    .CLK(CLK_bF$buf127),
    .D(_4656_),
    .Q(\datapath.registers.838[5] [8])
);

DFFPOSX1 _20766_ (
    .CLK(CLK_bF$buf126),
    .D(_4657_),
    .Q(\datapath.registers.838[5] [9])
);

DFFPOSX1 _20767_ (
    .CLK(CLK_bF$buf125),
    .D(_4627_),
    .Q(\datapath.registers.838[5] [10])
);

DFFPOSX1 _20768_ (
    .CLK(CLK_bF$buf124),
    .D(_4628_),
    .Q(\datapath.registers.838[5] [11])
);

DFFPOSX1 _20769_ (
    .CLK(CLK_bF$buf123),
    .D(_4629_),
    .Q(\datapath.registers.838[5] [12])
);

DFFPOSX1 _20770_ (
    .CLK(CLK_bF$buf122),
    .D(_4630_),
    .Q(\datapath.registers.838[5] [13])
);

DFFPOSX1 _20771_ (
    .CLK(CLK_bF$buf121),
    .D(_4631_),
    .Q(\datapath.registers.838[5] [14])
);

DFFPOSX1 _20772_ (
    .CLK(CLK_bF$buf120),
    .D(_4632_),
    .Q(\datapath.registers.838[5] [15])
);

DFFPOSX1 _20773_ (
    .CLK(CLK_bF$buf119),
    .D(_4633_),
    .Q(\datapath.registers.838[5] [16])
);

DFFPOSX1 _20774_ (
    .CLK(CLK_bF$buf118),
    .D(_4634_),
    .Q(\datapath.registers.838[5] [17])
);

DFFPOSX1 _20775_ (
    .CLK(CLK_bF$buf117),
    .D(_4635_),
    .Q(\datapath.registers.838[5] [18])
);

DFFPOSX1 _20776_ (
    .CLK(CLK_bF$buf116),
    .D(_4636_),
    .Q(\datapath.registers.838[5] [19])
);

DFFPOSX1 _20777_ (
    .CLK(CLK_bF$buf115),
    .D(_4638_),
    .Q(\datapath.registers.838[5] [20])
);

DFFPOSX1 _20778_ (
    .CLK(CLK_bF$buf114),
    .D(_4639_),
    .Q(\datapath.registers.838[5] [21])
);

DFFPOSX1 _20779_ (
    .CLK(CLK_bF$buf113),
    .D(_4640_),
    .Q(\datapath.registers.838[5] [22])
);

DFFPOSX1 _20780_ (
    .CLK(CLK_bF$buf112),
    .D(_4641_),
    .Q(\datapath.registers.838[5] [23])
);

DFFPOSX1 _20781_ (
    .CLK(CLK_bF$buf111),
    .D(_4642_),
    .Q(\datapath.registers.838[5] [24])
);

DFFPOSX1 _20782_ (
    .CLK(CLK_bF$buf110),
    .D(_4643_),
    .Q(\datapath.registers.838[5] [25])
);

DFFPOSX1 _20783_ (
    .CLK(CLK_bF$buf109),
    .D(_4644_),
    .Q(\datapath.registers.838[5] [26])
);

DFFPOSX1 _20784_ (
    .CLK(CLK_bF$buf108),
    .D(_4645_),
    .Q(\datapath.registers.838[5] [27])
);

DFFPOSX1 _20785_ (
    .CLK(CLK_bF$buf107),
    .D(_4646_),
    .Q(\datapath.registers.838[5] [28])
);

DFFPOSX1 _20786_ (
    .CLK(CLK_bF$buf106),
    .D(_4647_),
    .Q(\datapath.registers.838[5] [29])
);

DFFPOSX1 _20787_ (
    .CLK(CLK_bF$buf105),
    .D(_4649_),
    .Q(\datapath.registers.838[5] [30])
);

DFFPOSX1 _20788_ (
    .CLK(CLK_bF$buf104),
    .D(_4650_),
    .Q(\datapath.registers.838[5] [31])
);

DFFPOSX1 _20789_ (
    .CLK(CLK_bF$buf103),
    .D(_4530_),
    .Q(\datapath.registers.838[31] [0])
);

DFFPOSX1 _20790_ (
    .CLK(CLK_bF$buf102),
    .D(_4541_),
    .Q(\datapath.registers.838[31] [1])
);

DFFPOSX1 _20791_ (
    .CLK(CLK_bF$buf101),
    .D(_4552_),
    .Q(\datapath.registers.838[31] [2])
);

DFFPOSX1 _20792_ (
    .CLK(CLK_bF$buf100),
    .D(_4555_),
    .Q(\datapath.registers.838[31] [3])
);

DFFPOSX1 _20793_ (
    .CLK(CLK_bF$buf99),
    .D(_4556_),
    .Q(\datapath.registers.838[31] [4])
);

DFFPOSX1 _20794_ (
    .CLK(CLK_bF$buf98),
    .D(_4557_),
    .Q(\datapath.registers.838[31] [5])
);

DFFPOSX1 _20795_ (
    .CLK(CLK_bF$buf97),
    .D(_4558_),
    .Q(\datapath.registers.838[31] [6])
);

DFFPOSX1 _20796_ (
    .CLK(CLK_bF$buf96),
    .D(_4559_),
    .Q(\datapath.registers.838[31] [7])
);

DFFPOSX1 _20797_ (
    .CLK(CLK_bF$buf95),
    .D(_4560_),
    .Q(\datapath.registers.838[31] [8])
);

DFFPOSX1 _20798_ (
    .CLK(CLK_bF$buf94),
    .D(_4561_),
    .Q(\datapath.registers.838[31] [9])
);

DFFPOSX1 _20799_ (
    .CLK(CLK_bF$buf93),
    .D(_4531_),
    .Q(\datapath.registers.838[31] [10])
);

DFFPOSX1 _20800_ (
    .CLK(CLK_bF$buf92),
    .D(_4532_),
    .Q(\datapath.registers.838[31] [11])
);

DFFPOSX1 _20801_ (
    .CLK(CLK_bF$buf91),
    .D(_4533_),
    .Q(\datapath.registers.838[31] [12])
);

DFFPOSX1 _20802_ (
    .CLK(CLK_bF$buf90),
    .D(_4534_),
    .Q(\datapath.registers.838[31] [13])
);

DFFPOSX1 _20803_ (
    .CLK(CLK_bF$buf89),
    .D(_4535_),
    .Q(\datapath.registers.838[31] [14])
);

DFFPOSX1 _20804_ (
    .CLK(CLK_bF$buf88),
    .D(_4536_),
    .Q(\datapath.registers.838[31] [15])
);

DFFPOSX1 _20805_ (
    .CLK(CLK_bF$buf87),
    .D(_4537_),
    .Q(\datapath.registers.838[31] [16])
);

DFFPOSX1 _20806_ (
    .CLK(CLK_bF$buf86),
    .D(_4538_),
    .Q(\datapath.registers.838[31] [17])
);

DFFPOSX1 _20807_ (
    .CLK(CLK_bF$buf85),
    .D(_4539_),
    .Q(\datapath.registers.838[31] [18])
);

DFFPOSX1 _20808_ (
    .CLK(CLK_bF$buf84),
    .D(_4540_),
    .Q(\datapath.registers.838[31] [19])
);

DFFPOSX1 _20809_ (
    .CLK(CLK_bF$buf83),
    .D(_4542_),
    .Q(\datapath.registers.838[31] [20])
);

DFFPOSX1 _20810_ (
    .CLK(CLK_bF$buf82),
    .D(_4543_),
    .Q(\datapath.registers.838[31] [21])
);

DFFPOSX1 _20811_ (
    .CLK(CLK_bF$buf81),
    .D(_4544_),
    .Q(\datapath.registers.838[31] [22])
);

DFFPOSX1 _20812_ (
    .CLK(CLK_bF$buf80),
    .D(_4545_),
    .Q(\datapath.registers.838[31] [23])
);

DFFPOSX1 _20813_ (
    .CLK(CLK_bF$buf79),
    .D(_4546_),
    .Q(\datapath.registers.838[31] [24])
);

DFFPOSX1 _20814_ (
    .CLK(CLK_bF$buf78),
    .D(_4547_),
    .Q(\datapath.registers.838[31] [25])
);

DFFPOSX1 _20815_ (
    .CLK(CLK_bF$buf77),
    .D(_4548_),
    .Q(\datapath.registers.838[31] [26])
);

DFFPOSX1 _20816_ (
    .CLK(CLK_bF$buf76),
    .D(_4549_),
    .Q(\datapath.registers.838[31] [27])
);

DFFPOSX1 _20817_ (
    .CLK(CLK_bF$buf75),
    .D(_4550_),
    .Q(\datapath.registers.838[31] [28])
);

DFFPOSX1 _20818_ (
    .CLK(CLK_bF$buf74),
    .D(_4551_),
    .Q(\datapath.registers.838[31] [29])
);

DFFPOSX1 _20819_ (
    .CLK(CLK_bF$buf73),
    .D(_4553_),
    .Q(\datapath.registers.838[31] [30])
);

DFFPOSX1 _20820_ (
    .CLK(CLK_bF$buf72),
    .D(_4554_),
    .Q(\datapath.registers.838[31] [31])
);

DFFPOSX1 _20821_ (
    .CLK(CLK_bF$buf71),
    .D(_4498_),
    .Q(\datapath.registers.838[30] [0])
);

DFFPOSX1 _20822_ (
    .CLK(CLK_bF$buf70),
    .D(_4509_),
    .Q(\datapath.registers.838[30] [1])
);

DFFPOSX1 _20823_ (
    .CLK(CLK_bF$buf69),
    .D(_4520_),
    .Q(\datapath.registers.838[30] [2])
);

DFFPOSX1 _20824_ (
    .CLK(CLK_bF$buf68),
    .D(_4523_),
    .Q(\datapath.registers.838[30] [3])
);

DFFPOSX1 _20825_ (
    .CLK(CLK_bF$buf67),
    .D(_4524_),
    .Q(\datapath.registers.838[30] [4])
);

DFFPOSX1 _20826_ (
    .CLK(CLK_bF$buf66),
    .D(_4525_),
    .Q(\datapath.registers.838[30] [5])
);

DFFPOSX1 _20827_ (
    .CLK(CLK_bF$buf65),
    .D(_4526_),
    .Q(\datapath.registers.838[30] [6])
);

DFFPOSX1 _20828_ (
    .CLK(CLK_bF$buf64),
    .D(_4527_),
    .Q(\datapath.registers.838[30] [7])
);

DFFPOSX1 _20829_ (
    .CLK(CLK_bF$buf63),
    .D(_4528_),
    .Q(\datapath.registers.838[30] [8])
);

DFFPOSX1 _20830_ (
    .CLK(CLK_bF$buf62),
    .D(_4529_),
    .Q(\datapath.registers.838[30] [9])
);

DFFPOSX1 _20831_ (
    .CLK(CLK_bF$buf61),
    .D(_4499_),
    .Q(\datapath.registers.838[30] [10])
);

DFFPOSX1 _20832_ (
    .CLK(CLK_bF$buf60),
    .D(_4500_),
    .Q(\datapath.registers.838[30] [11])
);

DFFPOSX1 _20833_ (
    .CLK(CLK_bF$buf59),
    .D(_4501_),
    .Q(\datapath.registers.838[30] [12])
);

DFFPOSX1 _20834_ (
    .CLK(CLK_bF$buf58),
    .D(_4502_),
    .Q(\datapath.registers.838[30] [13])
);

DFFPOSX1 _20835_ (
    .CLK(CLK_bF$buf57),
    .D(_4503_),
    .Q(\datapath.registers.838[30] [14])
);

DFFPOSX1 _20836_ (
    .CLK(CLK_bF$buf56),
    .D(_4504_),
    .Q(\datapath.registers.838[30] [15])
);

DFFPOSX1 _20837_ (
    .CLK(CLK_bF$buf55),
    .D(_4505_),
    .Q(\datapath.registers.838[30] [16])
);

DFFPOSX1 _20838_ (
    .CLK(CLK_bF$buf54),
    .D(_4506_),
    .Q(\datapath.registers.838[30] [17])
);

DFFPOSX1 _20839_ (
    .CLK(CLK_bF$buf53),
    .D(_4507_),
    .Q(\datapath.registers.838[30] [18])
);

DFFPOSX1 _20840_ (
    .CLK(CLK_bF$buf52),
    .D(_4508_),
    .Q(\datapath.registers.838[30] [19])
);

DFFPOSX1 _20841_ (
    .CLK(CLK_bF$buf51),
    .D(_4510_),
    .Q(\datapath.registers.838[30] [20])
);

DFFPOSX1 _20842_ (
    .CLK(CLK_bF$buf50),
    .D(_4511_),
    .Q(\datapath.registers.838[30] [21])
);

DFFPOSX1 _20843_ (
    .CLK(CLK_bF$buf49),
    .D(_4512_),
    .Q(\datapath.registers.838[30] [22])
);

DFFPOSX1 _20844_ (
    .CLK(CLK_bF$buf48),
    .D(_4513_),
    .Q(\datapath.registers.838[30] [23])
);

DFFPOSX1 _20845_ (
    .CLK(CLK_bF$buf47),
    .D(_4514_),
    .Q(\datapath.registers.838[30] [24])
);

DFFPOSX1 _20846_ (
    .CLK(CLK_bF$buf46),
    .D(_4515_),
    .Q(\datapath.registers.838[30] [25])
);

DFFPOSX1 _20847_ (
    .CLK(CLK_bF$buf45),
    .D(_4516_),
    .Q(\datapath.registers.838[30] [26])
);

DFFPOSX1 _20848_ (
    .CLK(CLK_bF$buf44),
    .D(_4517_),
    .Q(\datapath.registers.838[30] [27])
);

DFFPOSX1 _20849_ (
    .CLK(CLK_bF$buf43),
    .D(_4518_),
    .Q(\datapath.registers.838[30] [28])
);

DFFPOSX1 _20850_ (
    .CLK(CLK_bF$buf42),
    .D(_4519_),
    .Q(\datapath.registers.838[30] [29])
);

DFFPOSX1 _20851_ (
    .CLK(CLK_bF$buf41),
    .D(_4521_),
    .Q(\datapath.registers.838[30] [30])
);

DFFPOSX1 _20852_ (
    .CLK(CLK_bF$buf40),
    .D(_4522_),
    .Q(\datapath.registers.838[30] [31])
);

DFFPOSX1 _20853_ (
    .CLK(CLK_bF$buf39),
    .D(_4434_),
    .Q(\datapath.registers.838[29] [0])
);

DFFPOSX1 _20854_ (
    .CLK(CLK_bF$buf38),
    .D(_4445_),
    .Q(\datapath.registers.838[29] [1])
);

DFFPOSX1 _20855_ (
    .CLK(CLK_bF$buf37),
    .D(_4456_),
    .Q(\datapath.registers.838[29] [2])
);

DFFPOSX1 _20856_ (
    .CLK(CLK_bF$buf36),
    .D(_4459_),
    .Q(\datapath.registers.838[29] [3])
);

DFFPOSX1 _20857_ (
    .CLK(CLK_bF$buf35),
    .D(_4460_),
    .Q(\datapath.registers.838[29] [4])
);

DFFPOSX1 _20858_ (
    .CLK(CLK_bF$buf34),
    .D(_4461_),
    .Q(\datapath.registers.838[29] [5])
);

DFFPOSX1 _20859_ (
    .CLK(CLK_bF$buf33),
    .D(_4462_),
    .Q(\datapath.registers.838[29] [6])
);

DFFPOSX1 _20860_ (
    .CLK(CLK_bF$buf32),
    .D(_4463_),
    .Q(\datapath.registers.838[29] [7])
);

DFFPOSX1 _20861_ (
    .CLK(CLK_bF$buf31),
    .D(_4464_),
    .Q(\datapath.registers.838[29] [8])
);

DFFPOSX1 _20862_ (
    .CLK(CLK_bF$buf30),
    .D(_4465_),
    .Q(\datapath.registers.838[29] [9])
);

DFFPOSX1 _20863_ (
    .CLK(CLK_bF$buf29),
    .D(_4435_),
    .Q(\datapath.registers.838[29] [10])
);

DFFPOSX1 _20864_ (
    .CLK(CLK_bF$buf28),
    .D(_4436_),
    .Q(\datapath.registers.838[29] [11])
);

DFFPOSX1 _20865_ (
    .CLK(CLK_bF$buf27),
    .D(_4437_),
    .Q(\datapath.registers.838[29] [12])
);

DFFPOSX1 _20866_ (
    .CLK(CLK_bF$buf26),
    .D(_4438_),
    .Q(\datapath.registers.838[29] [13])
);

DFFPOSX1 _20867_ (
    .CLK(CLK_bF$buf25),
    .D(_4439_),
    .Q(\datapath.registers.838[29] [14])
);

DFFPOSX1 _20868_ (
    .CLK(CLK_bF$buf24),
    .D(_4440_),
    .Q(\datapath.registers.838[29] [15])
);

DFFPOSX1 _20869_ (
    .CLK(CLK_bF$buf23),
    .D(_4441_),
    .Q(\datapath.registers.838[29] [16])
);

DFFPOSX1 _20870_ (
    .CLK(CLK_bF$buf22),
    .D(_4442_),
    .Q(\datapath.registers.838[29] [17])
);

DFFPOSX1 _20871_ (
    .CLK(CLK_bF$buf21),
    .D(_4443_),
    .Q(\datapath.registers.838[29] [18])
);

DFFPOSX1 _20872_ (
    .CLK(CLK_bF$buf20),
    .D(_4444_),
    .Q(\datapath.registers.838[29] [19])
);

DFFPOSX1 _20873_ (
    .CLK(CLK_bF$buf19),
    .D(_4446_),
    .Q(\datapath.registers.838[29] [20])
);

DFFPOSX1 _20874_ (
    .CLK(CLK_bF$buf18),
    .D(_4447_),
    .Q(\datapath.registers.838[29] [21])
);

DFFPOSX1 _20875_ (
    .CLK(CLK_bF$buf17),
    .D(_4448_),
    .Q(\datapath.registers.838[29] [22])
);

DFFPOSX1 _20876_ (
    .CLK(CLK_bF$buf16),
    .D(_4449_),
    .Q(\datapath.registers.838[29] [23])
);

DFFPOSX1 _20877_ (
    .CLK(CLK_bF$buf15),
    .D(_4450_),
    .Q(\datapath.registers.838[29] [24])
);

DFFPOSX1 _20878_ (
    .CLK(CLK_bF$buf14),
    .D(_4451_),
    .Q(\datapath.registers.838[29] [25])
);

DFFPOSX1 _20879_ (
    .CLK(CLK_bF$buf13),
    .D(_4452_),
    .Q(\datapath.registers.838[29] [26])
);

DFFPOSX1 _20880_ (
    .CLK(CLK_bF$buf12),
    .D(_4453_),
    .Q(\datapath.registers.838[29] [27])
);

DFFPOSX1 _20881_ (
    .CLK(CLK_bF$buf11),
    .D(_4454_),
    .Q(\datapath.registers.838[29] [28])
);

DFFPOSX1 _20882_ (
    .CLK(CLK_bF$buf10),
    .D(_4455_),
    .Q(\datapath.registers.838[29] [29])
);

DFFPOSX1 _20883_ (
    .CLK(CLK_bF$buf9),
    .D(_4457_),
    .Q(\datapath.registers.838[29] [30])
);

DFFPOSX1 _20884_ (
    .CLK(CLK_bF$buf8),
    .D(_4458_),
    .Q(\datapath.registers.838[29] [31])
);

DFFPOSX1 _20885_ (
    .CLK(CLK_bF$buf7),
    .D(_4562_),
    .Q(\datapath.registers.838[3] [0])
);

DFFPOSX1 _20886_ (
    .CLK(CLK_bF$buf6),
    .D(_4573_),
    .Q(\datapath.registers.838[3] [1])
);

DFFPOSX1 _20887_ (
    .CLK(CLK_bF$buf5),
    .D(_4584_),
    .Q(\datapath.registers.838[3] [2])
);

DFFPOSX1 _20888_ (
    .CLK(CLK_bF$buf4),
    .D(_4587_),
    .Q(\datapath.registers.838[3] [3])
);

DFFPOSX1 _20889_ (
    .CLK(CLK_bF$buf3),
    .D(_4588_),
    .Q(\datapath.registers.838[3] [4])
);

DFFPOSX1 _20890_ (
    .CLK(CLK_bF$buf2),
    .D(_4589_),
    .Q(\datapath.registers.838[3] [5])
);

DFFPOSX1 _20891_ (
    .CLK(CLK_bF$buf1),
    .D(_4590_),
    .Q(\datapath.registers.838[3] [6])
);

DFFPOSX1 _20892_ (
    .CLK(CLK_bF$buf0),
    .D(_4591_),
    .Q(\datapath.registers.838[3] [7])
);

DFFPOSX1 _20893_ (
    .CLK(CLK_bF$buf151),
    .D(_4592_),
    .Q(\datapath.registers.838[3] [8])
);

DFFPOSX1 _20894_ (
    .CLK(CLK_bF$buf150),
    .D(_4593_),
    .Q(\datapath.registers.838[3] [9])
);

DFFPOSX1 _20895_ (
    .CLK(CLK_bF$buf149),
    .D(_4563_),
    .Q(\datapath.registers.838[3] [10])
);

DFFPOSX1 _20896_ (
    .CLK(CLK_bF$buf148),
    .D(_4564_),
    .Q(\datapath.registers.838[3] [11])
);

DFFPOSX1 _20897_ (
    .CLK(CLK_bF$buf147),
    .D(_4565_),
    .Q(\datapath.registers.838[3] [12])
);

DFFPOSX1 _20898_ (
    .CLK(CLK_bF$buf146),
    .D(_4566_),
    .Q(\datapath.registers.838[3] [13])
);

DFFPOSX1 _20899_ (
    .CLK(CLK_bF$buf145),
    .D(_4567_),
    .Q(\datapath.registers.838[3] [14])
);

DFFPOSX1 _20900_ (
    .CLK(CLK_bF$buf144),
    .D(_4568_),
    .Q(\datapath.registers.838[3] [15])
);

DFFPOSX1 _20901_ (
    .CLK(CLK_bF$buf143),
    .D(_4569_),
    .Q(\datapath.registers.838[3] [16])
);

DFFPOSX1 _20902_ (
    .CLK(CLK_bF$buf142),
    .D(_4570_),
    .Q(\datapath.registers.838[3] [17])
);

DFFPOSX1 _20903_ (
    .CLK(CLK_bF$buf141),
    .D(_4571_),
    .Q(\datapath.registers.838[3] [18])
);

DFFPOSX1 _20904_ (
    .CLK(CLK_bF$buf140),
    .D(_4572_),
    .Q(\datapath.registers.838[3] [19])
);

DFFPOSX1 _20905_ (
    .CLK(CLK_bF$buf139),
    .D(_4574_),
    .Q(\datapath.registers.838[3] [20])
);

DFFPOSX1 _20906_ (
    .CLK(CLK_bF$buf138),
    .D(_4575_),
    .Q(\datapath.registers.838[3] [21])
);

DFFPOSX1 _20907_ (
    .CLK(CLK_bF$buf137),
    .D(_4576_),
    .Q(\datapath.registers.838[3] [22])
);

DFFPOSX1 _20908_ (
    .CLK(CLK_bF$buf136),
    .D(_4577_),
    .Q(\datapath.registers.838[3] [23])
);

DFFPOSX1 _20909_ (
    .CLK(CLK_bF$buf135),
    .D(_4578_),
    .Q(\datapath.registers.838[3] [24])
);

DFFPOSX1 _20910_ (
    .CLK(CLK_bF$buf134),
    .D(_4579_),
    .Q(\datapath.registers.838[3] [25])
);

DFFPOSX1 _20911_ (
    .CLK(CLK_bF$buf133),
    .D(_4580_),
    .Q(\datapath.registers.838[3] [26])
);

DFFPOSX1 _20912_ (
    .CLK(CLK_bF$buf132),
    .D(_4581_),
    .Q(\datapath.registers.838[3] [27])
);

DFFPOSX1 _20913_ (
    .CLK(CLK_bF$buf131),
    .D(_4582_),
    .Q(\datapath.registers.838[3] [28])
);

DFFPOSX1 _20914_ (
    .CLK(CLK_bF$buf130),
    .D(_4583_),
    .Q(\datapath.registers.838[3] [29])
);

DFFPOSX1 _20915_ (
    .CLK(CLK_bF$buf129),
    .D(_4585_),
    .Q(\datapath.registers.838[3] [30])
);

DFFPOSX1 _20916_ (
    .CLK(CLK_bF$buf128),
    .D(_4586_),
    .Q(\datapath.registers.838[3] [31])
);

DFFPOSX1 _20917_ (
    .CLK(CLK_bF$buf127),
    .D(_4114_),
    .Q(\datapath.registers.838[1] [0])
);

DFFPOSX1 _20918_ (
    .CLK(CLK_bF$buf126),
    .D(_4125_),
    .Q(\datapath.registers.838[1] [1])
);

DFFPOSX1 _20919_ (
    .CLK(CLK_bF$buf125),
    .D(_4136_),
    .Q(\datapath.registers.838[1] [2])
);

DFFPOSX1 _20920_ (
    .CLK(CLK_bF$buf124),
    .D(_4139_),
    .Q(\datapath.registers.838[1] [3])
);

DFFPOSX1 _20921_ (
    .CLK(CLK_bF$buf123),
    .D(_4140_),
    .Q(\datapath.registers.838[1] [4])
);

DFFPOSX1 _20922_ (
    .CLK(CLK_bF$buf122),
    .D(_4141_),
    .Q(\datapath.registers.838[1] [5])
);

DFFPOSX1 _20923_ (
    .CLK(CLK_bF$buf121),
    .D(_4142_),
    .Q(\datapath.registers.838[1] [6])
);

DFFPOSX1 _20924_ (
    .CLK(CLK_bF$buf120),
    .D(_4143_),
    .Q(\datapath.registers.838[1] [7])
);

DFFPOSX1 _20925_ (
    .CLK(CLK_bF$buf119),
    .D(_4144_),
    .Q(\datapath.registers.838[1] [8])
);

DFFPOSX1 _20926_ (
    .CLK(CLK_bF$buf118),
    .D(_4145_),
    .Q(\datapath.registers.838[1] [9])
);

DFFPOSX1 _20927_ (
    .CLK(CLK_bF$buf117),
    .D(_4115_),
    .Q(\datapath.registers.838[1] [10])
);

DFFPOSX1 _20928_ (
    .CLK(CLK_bF$buf116),
    .D(_4116_),
    .Q(\datapath.registers.838[1] [11])
);

DFFPOSX1 _20929_ (
    .CLK(CLK_bF$buf115),
    .D(_4117_),
    .Q(\datapath.registers.838[1] [12])
);

DFFPOSX1 _20930_ (
    .CLK(CLK_bF$buf114),
    .D(_4118_),
    .Q(\datapath.registers.838[1] [13])
);

DFFPOSX1 _20931_ (
    .CLK(CLK_bF$buf113),
    .D(_4119_),
    .Q(\datapath.registers.838[1] [14])
);

DFFPOSX1 _20932_ (
    .CLK(CLK_bF$buf112),
    .D(_4120_),
    .Q(\datapath.registers.838[1] [15])
);

DFFPOSX1 _20933_ (
    .CLK(CLK_bF$buf111),
    .D(_4121_),
    .Q(\datapath.registers.838[1] [16])
);

DFFPOSX1 _20934_ (
    .CLK(CLK_bF$buf110),
    .D(_4122_),
    .Q(\datapath.registers.838[1] [17])
);

DFFPOSX1 _20935_ (
    .CLK(CLK_bF$buf109),
    .D(_4123_),
    .Q(\datapath.registers.838[1] [18])
);

DFFPOSX1 _20936_ (
    .CLK(CLK_bF$buf108),
    .D(_4124_),
    .Q(\datapath.registers.838[1] [19])
);

DFFPOSX1 _20937_ (
    .CLK(CLK_bF$buf107),
    .D(_4126_),
    .Q(\datapath.registers.838[1] [20])
);

DFFPOSX1 _20938_ (
    .CLK(CLK_bF$buf106),
    .D(_4127_),
    .Q(\datapath.registers.838[1] [21])
);

DFFPOSX1 _20939_ (
    .CLK(CLK_bF$buf105),
    .D(_4128_),
    .Q(\datapath.registers.838[1] [22])
);

DFFPOSX1 _20940_ (
    .CLK(CLK_bF$buf104),
    .D(_4129_),
    .Q(\datapath.registers.838[1] [23])
);

DFFPOSX1 _20941_ (
    .CLK(CLK_bF$buf103),
    .D(_4130_),
    .Q(\datapath.registers.838[1] [24])
);

DFFPOSX1 _20942_ (
    .CLK(CLK_bF$buf102),
    .D(_4131_),
    .Q(\datapath.registers.838[1] [25])
);

DFFPOSX1 _20943_ (
    .CLK(CLK_bF$buf101),
    .D(_4132_),
    .Q(\datapath.registers.838[1] [26])
);

DFFPOSX1 _20944_ (
    .CLK(CLK_bF$buf100),
    .D(_4133_),
    .Q(\datapath.registers.838[1] [27])
);

DFFPOSX1 _20945_ (
    .CLK(CLK_bF$buf99),
    .D(_4134_),
    .Q(\datapath.registers.838[1] [28])
);

DFFPOSX1 _20946_ (
    .CLK(CLK_bF$buf98),
    .D(_4135_),
    .Q(\datapath.registers.838[1] [29])
);

DFFPOSX1 _20947_ (
    .CLK(CLK_bF$buf97),
    .D(_4137_),
    .Q(\datapath.registers.838[1] [30])
);

DFFPOSX1 _20948_ (
    .CLK(CLK_bF$buf96),
    .D(_4138_),
    .Q(\datapath.registers.838[1] [31])
);

DFFPOSX1 _20949_ (
    .CLK(CLK_bF$buf95),
    .D(_4178_),
    .Q(\datapath.registers.838[21] [0])
);

DFFPOSX1 _20950_ (
    .CLK(CLK_bF$buf94),
    .D(_4189_),
    .Q(\datapath.registers.838[21] [1])
);

DFFPOSX1 _20951_ (
    .CLK(CLK_bF$buf93),
    .D(_4200_),
    .Q(\datapath.registers.838[21] [2])
);

DFFPOSX1 _20952_ (
    .CLK(CLK_bF$buf92),
    .D(_4203_),
    .Q(\datapath.registers.838[21] [3])
);

DFFPOSX1 _20953_ (
    .CLK(CLK_bF$buf91),
    .D(_4204_),
    .Q(\datapath.registers.838[21] [4])
);

DFFPOSX1 _20954_ (
    .CLK(CLK_bF$buf90),
    .D(_4205_),
    .Q(\datapath.registers.838[21] [5])
);

DFFPOSX1 _20955_ (
    .CLK(CLK_bF$buf89),
    .D(_4206_),
    .Q(\datapath.registers.838[21] [6])
);

DFFPOSX1 _20956_ (
    .CLK(CLK_bF$buf88),
    .D(_4207_),
    .Q(\datapath.registers.838[21] [7])
);

DFFPOSX1 _20957_ (
    .CLK(CLK_bF$buf87),
    .D(_4208_),
    .Q(\datapath.registers.838[21] [8])
);

DFFPOSX1 _20958_ (
    .CLK(CLK_bF$buf86),
    .D(_4209_),
    .Q(\datapath.registers.838[21] [9])
);

DFFPOSX1 _20959_ (
    .CLK(CLK_bF$buf85),
    .D(_4179_),
    .Q(\datapath.registers.838[21] [10])
);

DFFPOSX1 _20960_ (
    .CLK(CLK_bF$buf84),
    .D(_4180_),
    .Q(\datapath.registers.838[21] [11])
);

DFFPOSX1 _20961_ (
    .CLK(CLK_bF$buf83),
    .D(_4181_),
    .Q(\datapath.registers.838[21] [12])
);

DFFPOSX1 _20962_ (
    .CLK(CLK_bF$buf82),
    .D(_4182_),
    .Q(\datapath.registers.838[21] [13])
);

DFFPOSX1 _20963_ (
    .CLK(CLK_bF$buf81),
    .D(_4183_),
    .Q(\datapath.registers.838[21] [14])
);

DFFPOSX1 _20964_ (
    .CLK(CLK_bF$buf80),
    .D(_4184_),
    .Q(\datapath.registers.838[21] [15])
);

DFFPOSX1 _20965_ (
    .CLK(CLK_bF$buf79),
    .D(_4185_),
    .Q(\datapath.registers.838[21] [16])
);

DFFPOSX1 _20966_ (
    .CLK(CLK_bF$buf78),
    .D(_4186_),
    .Q(\datapath.registers.838[21] [17])
);

DFFPOSX1 _20967_ (
    .CLK(CLK_bF$buf77),
    .D(_4187_),
    .Q(\datapath.registers.838[21] [18])
);

DFFPOSX1 _20968_ (
    .CLK(CLK_bF$buf76),
    .D(_4188_),
    .Q(\datapath.registers.838[21] [19])
);

DFFPOSX1 _20969_ (
    .CLK(CLK_bF$buf75),
    .D(_4190_),
    .Q(\datapath.registers.838[21] [20])
);

DFFPOSX1 _20970_ (
    .CLK(CLK_bF$buf74),
    .D(_4191_),
    .Q(\datapath.registers.838[21] [21])
);

DFFPOSX1 _20971_ (
    .CLK(CLK_bF$buf73),
    .D(_4192_),
    .Q(\datapath.registers.838[21] [22])
);

DFFPOSX1 _20972_ (
    .CLK(CLK_bF$buf72),
    .D(_4193_),
    .Q(\datapath.registers.838[21] [23])
);

DFFPOSX1 _20973_ (
    .CLK(CLK_bF$buf71),
    .D(_4194_),
    .Q(\datapath.registers.838[21] [24])
);

DFFPOSX1 _20974_ (
    .CLK(CLK_bF$buf70),
    .D(_4195_),
    .Q(\datapath.registers.838[21] [25])
);

DFFPOSX1 _20975_ (
    .CLK(CLK_bF$buf69),
    .D(_4196_),
    .Q(\datapath.registers.838[21] [26])
);

DFFPOSX1 _20976_ (
    .CLK(CLK_bF$buf68),
    .D(_4197_),
    .Q(\datapath.registers.838[21] [27])
);

DFFPOSX1 _20977_ (
    .CLK(CLK_bF$buf67),
    .D(_4198_),
    .Q(\datapath.registers.838[21] [28])
);

DFFPOSX1 _20978_ (
    .CLK(CLK_bF$buf66),
    .D(_4199_),
    .Q(\datapath.registers.838[21] [29])
);

DFFPOSX1 _20979_ (
    .CLK(CLK_bF$buf65),
    .D(_4201_),
    .Q(\datapath.registers.838[21] [30])
);

DFFPOSX1 _20980_ (
    .CLK(CLK_bF$buf64),
    .D(_4202_),
    .Q(\datapath.registers.838[21] [31])
);

DFFPOSX1 _20981_ (
    .CLK(CLK_bF$buf63),
    .D(_4050_),
    .Q(\datapath.registers.838[18] [0])
);

DFFPOSX1 _20982_ (
    .CLK(CLK_bF$buf62),
    .D(_4061_),
    .Q(\datapath.registers.838[18] [1])
);

DFFPOSX1 _20983_ (
    .CLK(CLK_bF$buf61),
    .D(_4072_),
    .Q(\datapath.registers.838[18] [2])
);

DFFPOSX1 _20984_ (
    .CLK(CLK_bF$buf60),
    .D(_4075_),
    .Q(\datapath.registers.838[18] [3])
);

DFFPOSX1 _20985_ (
    .CLK(CLK_bF$buf59),
    .D(_4076_),
    .Q(\datapath.registers.838[18] [4])
);

DFFPOSX1 _20986_ (
    .CLK(CLK_bF$buf58),
    .D(_4077_),
    .Q(\datapath.registers.838[18] [5])
);

DFFPOSX1 _20987_ (
    .CLK(CLK_bF$buf57),
    .D(_4078_),
    .Q(\datapath.registers.838[18] [6])
);

DFFPOSX1 _20988_ (
    .CLK(CLK_bF$buf56),
    .D(_4079_),
    .Q(\datapath.registers.838[18] [7])
);

DFFPOSX1 _20989_ (
    .CLK(CLK_bF$buf55),
    .D(_4080_),
    .Q(\datapath.registers.838[18] [8])
);

DFFPOSX1 _20990_ (
    .CLK(CLK_bF$buf54),
    .D(_4081_),
    .Q(\datapath.registers.838[18] [9])
);

DFFPOSX1 _20991_ (
    .CLK(CLK_bF$buf53),
    .D(_4051_),
    .Q(\datapath.registers.838[18] [10])
);

DFFPOSX1 _20992_ (
    .CLK(CLK_bF$buf52),
    .D(_4052_),
    .Q(\datapath.registers.838[18] [11])
);

DFFPOSX1 _20993_ (
    .CLK(CLK_bF$buf51),
    .D(_4053_),
    .Q(\datapath.registers.838[18] [12])
);

DFFPOSX1 _20994_ (
    .CLK(CLK_bF$buf50),
    .D(_4054_),
    .Q(\datapath.registers.838[18] [13])
);

DFFPOSX1 _20995_ (
    .CLK(CLK_bF$buf49),
    .D(_4055_),
    .Q(\datapath.registers.838[18] [14])
);

DFFPOSX1 _20996_ (
    .CLK(CLK_bF$buf48),
    .D(_4056_),
    .Q(\datapath.registers.838[18] [15])
);

DFFPOSX1 _20997_ (
    .CLK(CLK_bF$buf47),
    .D(_4057_),
    .Q(\datapath.registers.838[18] [16])
);

DFFPOSX1 _20998_ (
    .CLK(CLK_bF$buf46),
    .D(_4058_),
    .Q(\datapath.registers.838[18] [17])
);

DFFPOSX1 _20999_ (
    .CLK(CLK_bF$buf45),
    .D(_4059_),
    .Q(\datapath.registers.838[18] [18])
);

DFFPOSX1 _21000_ (
    .CLK(CLK_bF$buf44),
    .D(_4060_),
    .Q(\datapath.registers.838[18] [19])
);

DFFPOSX1 _21001_ (
    .CLK(CLK_bF$buf43),
    .D(_4062_),
    .Q(\datapath.registers.838[18] [20])
);

DFFPOSX1 _21002_ (
    .CLK(CLK_bF$buf42),
    .D(_4063_),
    .Q(\datapath.registers.838[18] [21])
);

DFFPOSX1 _21003_ (
    .CLK(CLK_bF$buf41),
    .D(_4064_),
    .Q(\datapath.registers.838[18] [22])
);

DFFPOSX1 _21004_ (
    .CLK(CLK_bF$buf40),
    .D(_4065_),
    .Q(\datapath.registers.838[18] [23])
);

DFFPOSX1 _21005_ (
    .CLK(CLK_bF$buf39),
    .D(_4066_),
    .Q(\datapath.registers.838[18] [24])
);

DFFPOSX1 _21006_ (
    .CLK(CLK_bF$buf38),
    .D(_4067_),
    .Q(\datapath.registers.838[18] [25])
);

DFFPOSX1 _21007_ (
    .CLK(CLK_bF$buf37),
    .D(_4068_),
    .Q(\datapath.registers.838[18] [26])
);

DFFPOSX1 _21008_ (
    .CLK(CLK_bF$buf36),
    .D(_4069_),
    .Q(\datapath.registers.838[18] [27])
);

DFFPOSX1 _21009_ (
    .CLK(CLK_bF$buf35),
    .D(_4070_),
    .Q(\datapath.registers.838[18] [28])
);

DFFPOSX1 _21010_ (
    .CLK(CLK_bF$buf34),
    .D(_4071_),
    .Q(\datapath.registers.838[18] [29])
);

DFFPOSX1 _21011_ (
    .CLK(CLK_bF$buf33),
    .D(_4073_),
    .Q(\datapath.registers.838[18] [30])
);

DFFPOSX1 _21012_ (
    .CLK(CLK_bF$buf32),
    .D(_4074_),
    .Q(\datapath.registers.838[18] [31])
);

DFFPOSX1 _21013_ (
    .CLK(CLK_bF$buf31),
    .D(_4082_),
    .Q(\datapath.registers.838[19] [0])
);

DFFPOSX1 _21014_ (
    .CLK(CLK_bF$buf30),
    .D(_4093_),
    .Q(\datapath.registers.838[19] [1])
);

DFFPOSX1 _21015_ (
    .CLK(CLK_bF$buf29),
    .D(_4104_),
    .Q(\datapath.registers.838[19] [2])
);

DFFPOSX1 _21016_ (
    .CLK(CLK_bF$buf28),
    .D(_4107_),
    .Q(\datapath.registers.838[19] [3])
);

DFFPOSX1 _21017_ (
    .CLK(CLK_bF$buf27),
    .D(_4108_),
    .Q(\datapath.registers.838[19] [4])
);

DFFPOSX1 _21018_ (
    .CLK(CLK_bF$buf26),
    .D(_4109_),
    .Q(\datapath.registers.838[19] [5])
);

DFFPOSX1 _21019_ (
    .CLK(CLK_bF$buf25),
    .D(_4110_),
    .Q(\datapath.registers.838[19] [6])
);

DFFPOSX1 _21020_ (
    .CLK(CLK_bF$buf24),
    .D(_4111_),
    .Q(\datapath.registers.838[19] [7])
);

DFFPOSX1 _21021_ (
    .CLK(CLK_bF$buf23),
    .D(_4112_),
    .Q(\datapath.registers.838[19] [8])
);

DFFPOSX1 _21022_ (
    .CLK(CLK_bF$buf22),
    .D(_4113_),
    .Q(\datapath.registers.838[19] [9])
);

DFFPOSX1 _21023_ (
    .CLK(CLK_bF$buf21),
    .D(_4083_),
    .Q(\datapath.registers.838[19] [10])
);

DFFPOSX1 _21024_ (
    .CLK(CLK_bF$buf20),
    .D(_4084_),
    .Q(\datapath.registers.838[19] [11])
);

DFFPOSX1 _21025_ (
    .CLK(CLK_bF$buf19),
    .D(_4085_),
    .Q(\datapath.registers.838[19] [12])
);

DFFPOSX1 _21026_ (
    .CLK(CLK_bF$buf18),
    .D(_4086_),
    .Q(\datapath.registers.838[19] [13])
);

DFFPOSX1 _21027_ (
    .CLK(CLK_bF$buf17),
    .D(_4087_),
    .Q(\datapath.registers.838[19] [14])
);

DFFPOSX1 _21028_ (
    .CLK(CLK_bF$buf16),
    .D(_4088_),
    .Q(\datapath.registers.838[19] [15])
);

DFFPOSX1 _21029_ (
    .CLK(CLK_bF$buf15),
    .D(_4089_),
    .Q(\datapath.registers.838[19] [16])
);

DFFPOSX1 _21030_ (
    .CLK(CLK_bF$buf14),
    .D(_4090_),
    .Q(\datapath.registers.838[19] [17])
);

DFFPOSX1 _21031_ (
    .CLK(CLK_bF$buf13),
    .D(_4091_),
    .Q(\datapath.registers.838[19] [18])
);

DFFPOSX1 _21032_ (
    .CLK(CLK_bF$buf12),
    .D(_4092_),
    .Q(\datapath.registers.838[19] [19])
);

DFFPOSX1 _21033_ (
    .CLK(CLK_bF$buf11),
    .D(_4094_),
    .Q(\datapath.registers.838[19] [20])
);

DFFPOSX1 _21034_ (
    .CLK(CLK_bF$buf10),
    .D(_4095_),
    .Q(\datapath.registers.838[19] [21])
);

DFFPOSX1 _21035_ (
    .CLK(CLK_bF$buf9),
    .D(_4096_),
    .Q(\datapath.registers.838[19] [22])
);

DFFPOSX1 _21036_ (
    .CLK(CLK_bF$buf8),
    .D(_4097_),
    .Q(\datapath.registers.838[19] [23])
);

DFFPOSX1 _21037_ (
    .CLK(CLK_bF$buf7),
    .D(_4098_),
    .Q(\datapath.registers.838[19] [24])
);

DFFPOSX1 _21038_ (
    .CLK(CLK_bF$buf6),
    .D(_4099_),
    .Q(\datapath.registers.838[19] [25])
);

DFFPOSX1 _21039_ (
    .CLK(CLK_bF$buf5),
    .D(_4100_),
    .Q(\datapath.registers.838[19] [26])
);

DFFPOSX1 _21040_ (
    .CLK(CLK_bF$buf4),
    .D(_4101_),
    .Q(\datapath.registers.838[19] [27])
);

DFFPOSX1 _21041_ (
    .CLK(CLK_bF$buf3),
    .D(_4102_),
    .Q(\datapath.registers.838[19] [28])
);

DFFPOSX1 _21042_ (
    .CLK(CLK_bF$buf2),
    .D(_4103_),
    .Q(\datapath.registers.838[19] [29])
);

DFFPOSX1 _21043_ (
    .CLK(CLK_bF$buf1),
    .D(_4105_),
    .Q(\datapath.registers.838[19] [30])
);

DFFPOSX1 _21044_ (
    .CLK(CLK_bF$buf0),
    .D(_4106_),
    .Q(\datapath.registers.838[19] [31])
);

DFFPOSX1 _21045_ (
    .CLK(CLK_bF$buf151),
    .D(_4018_),
    .Q(\datapath.registers.838[17] [0])
);

DFFPOSX1 _21046_ (
    .CLK(CLK_bF$buf150),
    .D(_4029_),
    .Q(\datapath.registers.838[17] [1])
);

DFFPOSX1 _21047_ (
    .CLK(CLK_bF$buf149),
    .D(_4040_),
    .Q(\datapath.registers.838[17] [2])
);

DFFPOSX1 _21048_ (
    .CLK(CLK_bF$buf148),
    .D(_4043_),
    .Q(\datapath.registers.838[17] [3])
);

DFFPOSX1 _21049_ (
    .CLK(CLK_bF$buf147),
    .D(_4044_),
    .Q(\datapath.registers.838[17] [4])
);

DFFPOSX1 _21050_ (
    .CLK(CLK_bF$buf146),
    .D(_4045_),
    .Q(\datapath.registers.838[17] [5])
);

DFFPOSX1 _21051_ (
    .CLK(CLK_bF$buf145),
    .D(_4046_),
    .Q(\datapath.registers.838[17] [6])
);

DFFPOSX1 _21052_ (
    .CLK(CLK_bF$buf144),
    .D(_4047_),
    .Q(\datapath.registers.838[17] [7])
);

DFFPOSX1 _21053_ (
    .CLK(CLK_bF$buf143),
    .D(_4048_),
    .Q(\datapath.registers.838[17] [8])
);

DFFPOSX1 _21054_ (
    .CLK(CLK_bF$buf142),
    .D(_4049_),
    .Q(\datapath.registers.838[17] [9])
);

DFFPOSX1 _21055_ (
    .CLK(CLK_bF$buf141),
    .D(_4019_),
    .Q(\datapath.registers.838[17] [10])
);

DFFPOSX1 _21056_ (
    .CLK(CLK_bF$buf140),
    .D(_4020_),
    .Q(\datapath.registers.838[17] [11])
);

DFFPOSX1 _21057_ (
    .CLK(CLK_bF$buf139),
    .D(_4021_),
    .Q(\datapath.registers.838[17] [12])
);

DFFPOSX1 _21058_ (
    .CLK(CLK_bF$buf138),
    .D(_4022_),
    .Q(\datapath.registers.838[17] [13])
);

DFFPOSX1 _21059_ (
    .CLK(CLK_bF$buf137),
    .D(_4023_),
    .Q(\datapath.registers.838[17] [14])
);

DFFPOSX1 _21060_ (
    .CLK(CLK_bF$buf136),
    .D(_4024_),
    .Q(\datapath.registers.838[17] [15])
);

DFFPOSX1 _21061_ (
    .CLK(CLK_bF$buf135),
    .D(_4025_),
    .Q(\datapath.registers.838[17] [16])
);

DFFPOSX1 _21062_ (
    .CLK(CLK_bF$buf134),
    .D(_4026_),
    .Q(\datapath.registers.838[17] [17])
);

DFFPOSX1 _21063_ (
    .CLK(CLK_bF$buf133),
    .D(_4027_),
    .Q(\datapath.registers.838[17] [18])
);

DFFPOSX1 _21064_ (
    .CLK(CLK_bF$buf132),
    .D(_4028_),
    .Q(\datapath.registers.838[17] [19])
);

DFFPOSX1 _21065_ (
    .CLK(CLK_bF$buf131),
    .D(_4030_),
    .Q(\datapath.registers.838[17] [20])
);

DFFPOSX1 _21066_ (
    .CLK(CLK_bF$buf130),
    .D(_4031_),
    .Q(\datapath.registers.838[17] [21])
);

DFFPOSX1 _21067_ (
    .CLK(CLK_bF$buf129),
    .D(_4032_),
    .Q(\datapath.registers.838[17] [22])
);

DFFPOSX1 _21068_ (
    .CLK(CLK_bF$buf128),
    .D(_4033_),
    .Q(\datapath.registers.838[17] [23])
);

DFFPOSX1 _21069_ (
    .CLK(CLK_bF$buf127),
    .D(_4034_),
    .Q(\datapath.registers.838[17] [24])
);

DFFPOSX1 _21070_ (
    .CLK(CLK_bF$buf126),
    .D(_4035_),
    .Q(\datapath.registers.838[17] [25])
);

DFFPOSX1 _21071_ (
    .CLK(CLK_bF$buf125),
    .D(_4036_),
    .Q(\datapath.registers.838[17] [26])
);

DFFPOSX1 _21072_ (
    .CLK(CLK_bF$buf124),
    .D(_4037_),
    .Q(\datapath.registers.838[17] [27])
);

DFFPOSX1 _21073_ (
    .CLK(CLK_bF$buf123),
    .D(_4038_),
    .Q(\datapath.registers.838[17] [28])
);

DFFPOSX1 _21074_ (
    .CLK(CLK_bF$buf122),
    .D(_4039_),
    .Q(\datapath.registers.838[17] [29])
);

DFFPOSX1 _21075_ (
    .CLK(CLK_bF$buf121),
    .D(_4041_),
    .Q(\datapath.registers.838[17] [30])
);

DFFPOSX1 _21076_ (
    .CLK(CLK_bF$buf120),
    .D(_4042_),
    .Q(\datapath.registers.838[17] [31])
);

DFFPOSX1 _21077_ (
    .CLK(CLK_bF$buf119),
    .D(_4402_),
    .Q(\datapath.registers.838[28] [0])
);

DFFPOSX1 _21078_ (
    .CLK(CLK_bF$buf118),
    .D(_4413_),
    .Q(\datapath.registers.838[28] [1])
);

DFFPOSX1 _21079_ (
    .CLK(CLK_bF$buf117),
    .D(_4424_),
    .Q(\datapath.registers.838[28] [2])
);

DFFPOSX1 _21080_ (
    .CLK(CLK_bF$buf116),
    .D(_4427_),
    .Q(\datapath.registers.838[28] [3])
);

DFFPOSX1 _21081_ (
    .CLK(CLK_bF$buf115),
    .D(_4428_),
    .Q(\datapath.registers.838[28] [4])
);

DFFPOSX1 _21082_ (
    .CLK(CLK_bF$buf114),
    .D(_4429_),
    .Q(\datapath.registers.838[28] [5])
);

DFFPOSX1 _21083_ (
    .CLK(CLK_bF$buf113),
    .D(_4430_),
    .Q(\datapath.registers.838[28] [6])
);

DFFPOSX1 _21084_ (
    .CLK(CLK_bF$buf112),
    .D(_4431_),
    .Q(\datapath.registers.838[28] [7])
);

DFFPOSX1 _21085_ (
    .CLK(CLK_bF$buf111),
    .D(_4432_),
    .Q(\datapath.registers.838[28] [8])
);

DFFPOSX1 _21086_ (
    .CLK(CLK_bF$buf110),
    .D(_4433_),
    .Q(\datapath.registers.838[28] [9])
);

DFFPOSX1 _21087_ (
    .CLK(CLK_bF$buf109),
    .D(_4403_),
    .Q(\datapath.registers.838[28] [10])
);

DFFPOSX1 _21088_ (
    .CLK(CLK_bF$buf108),
    .D(_4404_),
    .Q(\datapath.registers.838[28] [11])
);

DFFPOSX1 _21089_ (
    .CLK(CLK_bF$buf107),
    .D(_4405_),
    .Q(\datapath.registers.838[28] [12])
);

DFFPOSX1 _21090_ (
    .CLK(CLK_bF$buf106),
    .D(_4406_),
    .Q(\datapath.registers.838[28] [13])
);

DFFPOSX1 _21091_ (
    .CLK(CLK_bF$buf105),
    .D(_4407_),
    .Q(\datapath.registers.838[28] [14])
);

DFFPOSX1 _21092_ (
    .CLK(CLK_bF$buf104),
    .D(_4408_),
    .Q(\datapath.registers.838[28] [15])
);

DFFPOSX1 _21093_ (
    .CLK(CLK_bF$buf103),
    .D(_4409_),
    .Q(\datapath.registers.838[28] [16])
);

DFFPOSX1 _21094_ (
    .CLK(CLK_bF$buf102),
    .D(_4410_),
    .Q(\datapath.registers.838[28] [17])
);

DFFPOSX1 _21095_ (
    .CLK(CLK_bF$buf101),
    .D(_4411_),
    .Q(\datapath.registers.838[28] [18])
);

DFFPOSX1 _21096_ (
    .CLK(CLK_bF$buf100),
    .D(_4412_),
    .Q(\datapath.registers.838[28] [19])
);

DFFPOSX1 _21097_ (
    .CLK(CLK_bF$buf99),
    .D(_4414_),
    .Q(\datapath.registers.838[28] [20])
);

DFFPOSX1 _21098_ (
    .CLK(CLK_bF$buf98),
    .D(_4415_),
    .Q(\datapath.registers.838[28] [21])
);

DFFPOSX1 _21099_ (
    .CLK(CLK_bF$buf97),
    .D(_4416_),
    .Q(\datapath.registers.838[28] [22])
);

DFFPOSX1 _21100_ (
    .CLK(CLK_bF$buf96),
    .D(_4417_),
    .Q(\datapath.registers.838[28] [23])
);

DFFPOSX1 _21101_ (
    .CLK(CLK_bF$buf95),
    .D(_4418_),
    .Q(\datapath.registers.838[28] [24])
);

DFFPOSX1 _21102_ (
    .CLK(CLK_bF$buf94),
    .D(_4419_),
    .Q(\datapath.registers.838[28] [25])
);

DFFPOSX1 _21103_ (
    .CLK(CLK_bF$buf93),
    .D(_4420_),
    .Q(\datapath.registers.838[28] [26])
);

DFFPOSX1 _21104_ (
    .CLK(CLK_bF$buf92),
    .D(_4421_),
    .Q(\datapath.registers.838[28] [27])
);

DFFPOSX1 _21105_ (
    .CLK(CLK_bF$buf91),
    .D(_4422_),
    .Q(\datapath.registers.838[28] [28])
);

DFFPOSX1 _21106_ (
    .CLK(CLK_bF$buf90),
    .D(_4423_),
    .Q(\datapath.registers.838[28] [29])
);

DFFPOSX1 _21107_ (
    .CLK(CLK_bF$buf89),
    .D(_4425_),
    .Q(\datapath.registers.838[28] [30])
);

DFFPOSX1 _21108_ (
    .CLK(CLK_bF$buf88),
    .D(_4426_),
    .Q(\datapath.registers.838[28] [31])
);

BUFX2 _9191_ (
    .A(_0__0_bF$buf1),
    .Y(DMEM_ADDR[0])
);

BUFX2 _9192_ (
    .A(_0__1_bF$buf3),
    .Y(DMEM_ADDR[1])
);

BUFX2 _9193_ (
    .A(_0_[2]),
    .Y(DMEM_ADDR[2])
);

BUFX2 _9194_ (
    .A(_0_[3]),
    .Y(DMEM_ADDR[3])
);

BUFX2 _9195_ (
    .A(_0_[4]),
    .Y(DMEM_ADDR[4])
);

BUFX2 _9196_ (
    .A(_0_[5]),
    .Y(DMEM_ADDR[5])
);

BUFX2 _9197_ (
    .A(_0_[6]),
    .Y(DMEM_ADDR[6])
);

BUFX2 _9198_ (
    .A(_0_[7]),
    .Y(DMEM_ADDR[7])
);

BUFX2 _9199_ (
    .A(_0_[8]),
    .Y(DMEM_ADDR[8])
);

BUFX2 _9200_ (
    .A(_0_[9]),
    .Y(DMEM_ADDR[9])
);

BUFX2 _9201_ (
    .A(_0_[10]),
    .Y(DMEM_ADDR[10])
);

BUFX2 _9202_ (
    .A(_0_[11]),
    .Y(DMEM_ADDR[11])
);

BUFX2 _9203_ (
    .A(_0_[12]),
    .Y(DMEM_ADDR[12])
);

BUFX2 _9204_ (
    .A(_0_[13]),
    .Y(DMEM_ADDR[13])
);

BUFX2 _9205_ (
    .A(_0_[14]),
    .Y(DMEM_ADDR[14])
);

BUFX2 _9206_ (
    .A(_0_[15]),
    .Y(DMEM_ADDR[15])
);

BUFX2 _9207_ (
    .A(_0_[16]),
    .Y(DMEM_ADDR[16])
);

BUFX2 _9208_ (
    .A(_0_[17]),
    .Y(DMEM_ADDR[17])
);

BUFX2 _9209_ (
    .A(_0_[18]),
    .Y(DMEM_ADDR[18])
);

BUFX2 _9210_ (
    .A(_0_[19]),
    .Y(DMEM_ADDR[19])
);

BUFX2 _9211_ (
    .A(_0_[20]),
    .Y(DMEM_ADDR[20])
);

BUFX2 _9212_ (
    .A(_0_[21]),
    .Y(DMEM_ADDR[21])
);

BUFX2 _9213_ (
    .A(_0_[22]),
    .Y(DMEM_ADDR[22])
);

BUFX2 _9214_ (
    .A(_0_[23]),
    .Y(DMEM_ADDR[23])
);

BUFX2 _9215_ (
    .A(_0_[24]),
    .Y(DMEM_ADDR[24])
);

BUFX2 _9216_ (
    .A(_0_[25]),
    .Y(DMEM_ADDR[25])
);

BUFX2 _9217_ (
    .A(_0_[26]),
    .Y(DMEM_ADDR[26])
);

BUFX2 _9218_ (
    .A(_0_[27]),
    .Y(DMEM_ADDR[27])
);

BUFX2 _9219_ (
    .A(_0_[28]),
    .Y(DMEM_ADDR[28])
);

BUFX2 _9220_ (
    .A(_0_[29]),
    .Y(DMEM_ADDR[29])
);

BUFX2 _9221_ (
    .A(_0_[30]),
    .Y(DMEM_ADDR[30])
);

BUFX2 _9222_ (
    .A(_0_[31]),
    .Y(DMEM_ADDR[31])
);

BUFX2 _9223_ (
    .A(_1_[0]),
    .Y(DMEM_DATA_S[0])
);

BUFX2 _9224_ (
    .A(_1_[1]),
    .Y(DMEM_DATA_S[1])
);

BUFX2 _9225_ (
    .A(_1_[2]),
    .Y(DMEM_DATA_S[2])
);

BUFX2 _9226_ (
    .A(_1_[3]),
    .Y(DMEM_DATA_S[3])
);

BUFX2 _9227_ (
    .A(_1_[4]),
    .Y(DMEM_DATA_S[4])
);

BUFX2 _9228_ (
    .A(_1_[5]),
    .Y(DMEM_DATA_S[5])
);

BUFX2 _9229_ (
    .A(_1_[6]),
    .Y(DMEM_DATA_S[6])
);

BUFX2 _9230_ (
    .A(_1_[7]),
    .Y(DMEM_DATA_S[7])
);

BUFX2 _9231_ (
    .A(_1_[8]),
    .Y(DMEM_DATA_S[8])
);

BUFX2 _9232_ (
    .A(_1_[9]),
    .Y(DMEM_DATA_S[9])
);

BUFX2 _9233_ (
    .A(_1_[10]),
    .Y(DMEM_DATA_S[10])
);

BUFX2 _9234_ (
    .A(_1_[11]),
    .Y(DMEM_DATA_S[11])
);

BUFX2 _9235_ (
    .A(_1_[12]),
    .Y(DMEM_DATA_S[12])
);

BUFX2 _9236_ (
    .A(_1_[13]),
    .Y(DMEM_DATA_S[13])
);

BUFX2 _9237_ (
    .A(_1_[14]),
    .Y(DMEM_DATA_S[14])
);

BUFX2 _9238_ (
    .A(_1_[15]),
    .Y(DMEM_DATA_S[15])
);

BUFX2 _9239_ (
    .A(_1_[16]),
    .Y(DMEM_DATA_S[16])
);

BUFX2 _9240_ (
    .A(_1_[17]),
    .Y(DMEM_DATA_S[17])
);

BUFX2 _9241_ (
    .A(_1_[18]),
    .Y(DMEM_DATA_S[18])
);

BUFX2 _9242_ (
    .A(_1_[19]),
    .Y(DMEM_DATA_S[19])
);

BUFX2 _9243_ (
    .A(_1_[20]),
    .Y(DMEM_DATA_S[20])
);

BUFX2 _9244_ (
    .A(_1_[21]),
    .Y(DMEM_DATA_S[21])
);

BUFX2 _9245_ (
    .A(_1_[22]),
    .Y(DMEM_DATA_S[22])
);

BUFX2 _9246_ (
    .A(_1_[23]),
    .Y(DMEM_DATA_S[23])
);

BUFX2 _9247_ (
    .A(_1_[24]),
    .Y(DMEM_DATA_S[24])
);

BUFX2 _9248_ (
    .A(_1_[25]),
    .Y(DMEM_DATA_S[25])
);

BUFX2 _9249_ (
    .A(_1_[26]),
    .Y(DMEM_DATA_S[26])
);

BUFX2 _9250_ (
    .A(_1_[27]),
    .Y(DMEM_DATA_S[27])
);

BUFX2 _9251_ (
    .A(_1_[28]),
    .Y(DMEM_DATA_S[28])
);

BUFX2 _9252_ (
    .A(_1_[29]),
    .Y(DMEM_DATA_S[29])
);

BUFX2 _9253_ (
    .A(_1_[30]),
    .Y(DMEM_DATA_S[30])
);

BUFX2 _9254_ (
    .A(_1_[31]),
    .Y(DMEM_DATA_S[31])
);

BUFX2 _9255_ (
    .A(_2_),
    .Y(DMEM_WEN)
);

BUFX2 _9256_ (
    .A(\datapath.programcounter.pc [0]),
    .Y(IMEM_ADDR[0])
);

BUFX2 _9257_ (
    .A(\datapath.programcounter.pc [1]),
    .Y(IMEM_ADDR[1])
);

BUFX2 _9258_ (
    .A(\datapath.programcounter.pc [2]),
    .Y(IMEM_ADDR[2])
);

BUFX2 _9259_ (
    .A(\datapath.programcounter.pc [3]),
    .Y(IMEM_ADDR[3])
);

BUFX2 _9260_ (
    .A(\datapath.programcounter.pc [4]),
    .Y(IMEM_ADDR[4])
);

BUFX2 _9261_ (
    .A(\datapath.programcounter.pc [5]),
    .Y(IMEM_ADDR[5])
);

BUFX2 _9262_ (
    .A(\datapath.programcounter.pc [6]),
    .Y(IMEM_ADDR[6])
);

BUFX2 _9263_ (
    .A(\datapath.programcounter.pc [7]),
    .Y(IMEM_ADDR[7])
);

BUFX2 _9264_ (
    .A(\datapath.programcounter.pc [8]),
    .Y(IMEM_ADDR[8])
);

BUFX2 _9265_ (
    .A(\datapath.programcounter.pc [9]),
    .Y(IMEM_ADDR[9])
);

BUFX2 _9266_ (
    .A(\datapath.programcounter.pc [10]),
    .Y(IMEM_ADDR[10])
);

BUFX2 _9267_ (
    .A(\datapath.programcounter.pc [11]),
    .Y(IMEM_ADDR[11])
);

BUFX2 _9268_ (
    .A(\datapath.programcounter.pc [12]),
    .Y(IMEM_ADDR[12])
);

BUFX2 _9269_ (
    .A(\datapath.programcounter.pc [13]),
    .Y(IMEM_ADDR[13])
);

BUFX2 _9270_ (
    .A(\datapath.programcounter.pc [14]),
    .Y(IMEM_ADDR[14])
);

BUFX2 _9271_ (
    .A(\datapath.programcounter.pc [15]),
    .Y(IMEM_ADDR[15])
);

BUFX2 _9272_ (
    .A(\datapath.programcounter.pc [16]),
    .Y(IMEM_ADDR[16])
);

BUFX2 _9273_ (
    .A(\datapath.programcounter.pc [17]),
    .Y(IMEM_ADDR[17])
);

BUFX2 _9274_ (
    .A(\datapath.programcounter.pc [18]),
    .Y(IMEM_ADDR[18])
);

BUFX2 _9275_ (
    .A(\datapath.programcounter.pc [19]),
    .Y(IMEM_ADDR[19])
);

BUFX2 _9276_ (
    .A(\datapath.programcounter.pc [20]),
    .Y(IMEM_ADDR[20])
);

BUFX2 _9277_ (
    .A(\datapath.programcounter.pc [21]),
    .Y(IMEM_ADDR[21])
);

BUFX2 _9278_ (
    .A(\datapath.programcounter.pc [22]),
    .Y(IMEM_ADDR[22])
);

BUFX2 _9279_ (
    .A(\datapath.programcounter.pc [23]),
    .Y(IMEM_ADDR[23])
);

BUFX2 _9280_ (
    .A(\datapath.programcounter.pc [24]),
    .Y(IMEM_ADDR[24])
);

BUFX2 _9281_ (
    .A(\datapath.programcounter.pc [25]),
    .Y(IMEM_ADDR[25])
);

BUFX2 _9282_ (
    .A(\datapath.programcounter.pc [26]),
    .Y(IMEM_ADDR[26])
);

BUFX2 _9283_ (
    .A(\datapath.programcounter.pc [27]),
    .Y(IMEM_ADDR[27])
);

BUFX2 _9284_ (
    .A(\datapath.programcounter.pc [28]),
    .Y(IMEM_ADDR[28])
);

BUFX2 _9285_ (
    .A(\datapath.programcounter.pc [29]),
    .Y(IMEM_ADDR[29])
);

BUFX2 _9286_ (
    .A(\datapath.programcounter.pc [30]),
    .Y(IMEM_ADDR[30])
);

BUFX2 _9287_ (
    .A(\datapath.programcounter.pc [31]),
    .Y(IMEM_ADDR[31])
);

NAND2X1 _9288_ (
    .A(\datapath.idinstr [1]),
    .B(\datapath.idinstr [0]),
    .Y(_79_)
);

NOR3X1 _9289_ (
    .A(\datapath.idinstr [2]),
    .B(\datapath.idinstr [3]),
    .C(_79_),
    .Y(_80_)
);

NOR2X1 _9290_ (
    .A(\datapath.idinstr [4]),
    .B(\datapath.idinstr [6]),
    .Y(_81_)
);

NAND3X1 _9291_ (
    .A(\datapath.idinstr [5]),
    .B(_81_),
    .C(_80_),
    .Y(_4_)
);

NOR2X1 _9292_ (
    .A(\datapath.meminstr [3]),
    .B(\datapath.meminstr [2]),
    .Y(_82_)
);

NAND3X1 _9293_ (
    .A(\datapath.meminstr [1]),
    .B(\datapath.meminstr [0]),
    .C(_82_),
    .Y(_83_)
);

INVX1 _9294_ (
    .A(\datapath.meminstr [6]),
    .Y(_84_)
);

NOR2X1 _9295_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf2 ),
    .B(\datapath.meminstr [4]),
    .Y(_85_)
);

NAND3X1 _9296_ (
    .A(\datapath.meminstr [5]),
    .B(_84_),
    .C(_85_),
    .Y(_86_)
);

NOR2X1 _9297_ (
    .A(_83_),
    .B(_86_),
    .Y(_2_)
);

OR2X2 _9298_ (
    .A(\datapath.meminstr [13]),
    .B(\datapath.meminstr [14]),
    .Y(_87_)
);

NOR2X1 _9299_ (
    .A(\datapath.meminstr [12]),
    .B(_87_),
    .Y(_88_)
);

INVX1 _9300_ (
    .A(\controlunit.csrfile_trap_wen_bF$buf1 ),
    .Y(_89_)
);

AND2X2 _9301_ (
    .A(\datapath.meminstr [5]),
    .B(\datapath.meminstr [6]),
    .Y(_90_)
);

NAND3X1 _9302_ (
    .A(_89_),
    .B(\datapath.meminstr [4]),
    .C(_90_),
    .Y(_91_)
);

OR2X2 _9303_ (
    .A(_91_),
    .B(_83_),
    .Y(_92_)
);

NOR2X1 _9304_ (
    .A(_88_),
    .B(_92_),
    .Y(\controlunit.csrfile_wen )
);

INVX1 _9305_ (
    .A(\datapath.meminstr [21]),
    .Y(_93_)
);

NOR2X1 _9306_ (
    .A(\datapath.meminstr [20]),
    .B(_93_),
    .Y(_94_)
);

NAND3X1 _9307_ (
    .A(\datapath.meminstr [29]),
    .B(_94_),
    .C(_88_),
    .Y(_95_)
);

NOR2X1 _9308_ (
    .A(_95_),
    .B(_92_),
    .Y(\controlunit.mret )
);

INVX1 _9309_ (
    .A(\datapath.wbinstr [2]),
    .Y(_96_)
);

NAND2X1 _9310_ (
    .A(\datapath.wbinstr [1]),
    .B(\datapath.wbinstr [0]),
    .Y(_97_)
);

NOR2X1 _9311_ (
    .A(\datapath.wbinstr [3]),
    .B(_97_),
    .Y(_98_)
);

NAND2X1 _9312_ (
    .A(_96_),
    .B(_98_),
    .Y(_99_)
);

INVX1 _9313_ (
    .A(\datapath.wbinstr [4]),
    .Y(_100_)
);

NAND2X1 _9314_ (
    .A(\datapath.wbinstr [6]),
    .B(\datapath.wbinstr [5]),
    .Y(_101_)
);

OR2X2 _9315_ (
    .A(_101_),
    .B(_100_),
    .Y(_102_)
);

NOR2X1 _9316_ (
    .A(_102_),
    .B(_99_),
    .Y(_103_)
);

OR2X2 _9317_ (
    .A(\datapath.wbinstr [14]),
    .B(\datapath.wbinstr [12]),
    .Y(_104_)
);

OAI21X1 _9318_ (
    .A(\datapath.wbinstr [13]),
    .B(_104_),
    .C(_103_),
    .Y(_5_)
);

OR2X2 _9319_ (
    .A(_97_),
    .B(_96_),
    .Y(_6_)
);

NOR2X1 _9320_ (
    .A(_101_),
    .B(_6_),
    .Y(_7_)
);

INVX1 _9321_ (
    .A(_98_),
    .Y(_8_)
);

INVX1 _9322_ (
    .A(\datapath.wbinstr [6]),
    .Y(_9_)
);

NAND2X1 _9323_ (
    .A(\datapath.wbinstr [4]),
    .B(_9_),
    .Y(_10_)
);

NOR2X1 _9324_ (
    .A(\datapath.wbinstr [5]),
    .B(\datapath.wbinstr [4]),
    .Y(_11_)
);

NAND3X1 _9325_ (
    .A(_96_),
    .B(_9_),
    .C(_11_),
    .Y(_12_)
);

AOI21X1 _9326_ (
    .A(_12_),
    .B(_10_),
    .C(_8_),
    .Y(_13_)
);

AOI21X1 _9327_ (
    .A(_100_),
    .B(_7_),
    .C(_13_),
    .Y(_14_)
);

AOI21X1 _9328_ (
    .A(_5_),
    .B(_14_),
    .C(\datapath.regwbtrap ),
    .Y(\controlunit.regfile_wen )
);

INVX1 _9329_ (
    .A(\datapath.aluinstr [4]),
    .Y(_15_)
);

NAND3X1 _9330_ (
    .A(\datapath.aluinstr [5]),
    .B(\datapath.aluinstr [6]),
    .C(_15_),
    .Y(_16_)
);

NAND3X1 _9331_ (
    .A(\datapath.aluinstr [1]),
    .B(\datapath.aluinstr [0]),
    .C(\datapath.aluinstr [2]),
    .Y(_17_)
);

INVX1 _9332_ (
    .A(_17_),
    .Y(_18_)
);

NAND2X1 _9333_ (
    .A(\datapath.aluinstr [3]),
    .B(_18_),
    .Y(_19_)
);

NOR2X1 _9334_ (
    .A(_16_),
    .B(_19_),
    .Y(\controlunit.pc_sel [0])
);

OR2X2 _9335_ (
    .A(_17_),
    .B(\datapath.aluinstr [3]),
    .Y(_20_)
);

NOR2X1 _9336_ (
    .A(_16_),
    .B(_20_),
    .Y(\controlunit.pc_sel [1])
);

INVX1 _9337_ (
    .A(\datapath.idinstr [13]),
    .Y(_21_)
);

INVX1 _9338_ (
    .A(\datapath.idinstr [5]),
    .Y(_22_)
);

INVX1 _9339_ (
    .A(\datapath.idinstr [6]),
    .Y(_23_)
);

NOR3X1 _9340_ (
    .A(\datapath.idinstr [4]),
    .B(_22_),
    .C(_23_),
    .Y(_24_)
);

NAND2X1 _9341_ (
    .A(_80_),
    .B(_24_),
    .Y(_25_)
);

AND2X2 _9342_ (
    .A(_23_),
    .B(\datapath.idinstr [4]),
    .Y(_26_)
);

NAND3X1 _9343_ (
    .A(\datapath.idinstr [4]),
    .B(\datapath.idinstr [5]),
    .C(\datapath.idinstr [6]),
    .Y(_27_)
);

INVX1 _9344_ (
    .A(_27_),
    .Y(_28_)
);

OAI21X1 _9345_ (
    .A(_26_),
    .B(_28_),
    .C(_80_),
    .Y(_29_)
);

NOR2X1 _9346_ (
    .A(\datapath.idinstr [2]),
    .B(\datapath.idinstr [3]),
    .Y(_30_)
);

NAND3X1 _9347_ (
    .A(\datapath.idinstr [1]),
    .B(\datapath.idinstr [0]),
    .C(_30_),
    .Y(_31_)
);

NAND2X1 _9348_ (
    .A(\datapath.idinstr [4]),
    .B(_23_),
    .Y(_32_)
);

NOR2X1 _9349_ (
    .A(_32_),
    .B(_31_),
    .Y(_33_)
);

OAI21X1 _9350_ (
    .A(\datapath.idinstr [13]),
    .B(_33_),
    .C(\datapath.idinstr [12]),
    .Y(_34_)
);

OAI22X1 _9351_ (
    .A(_21_),
    .B(_25_),
    .C(_29_),
    .D(_34_),
    .Y(_3_[0])
);

INVX1 _9352_ (
    .A(\datapath.idinstr [3]),
    .Y(_35_)
);

NAND2X1 _9353_ (
    .A(\datapath.idinstr [2]),
    .B(_35_),
    .Y(_36_)
);

NOR2X1 _9354_ (
    .A(_79_),
    .B(_36_),
    .Y(_37_)
);

OAI21X1 _9355_ (
    .A(_80_),
    .B(_37_),
    .C(_24_),
    .Y(_38_)
);

NOR2X1 _9356_ (
    .A(\datapath.idinstr [5]),
    .B(_32_),
    .Y(_39_)
);

AND2X2 _9357_ (
    .A(_81_),
    .B(_22_),
    .Y(_40_)
);

AOI22X1 _9358_ (
    .A(_80_),
    .B(_40_),
    .C(_39_),
    .D(_37_),
    .Y(_41_)
);

NAND3X1 _9359_ (
    .A(_29_),
    .B(_41_),
    .C(_38_),
    .Y(_42_)
);

INVX1 _9360_ (
    .A(\datapath.idinstr [14]),
    .Y(_43_)
);

NAND2X1 _9361_ (
    .A(_21_),
    .B(_43_),
    .Y(_44_)
);

NAND2X1 _9362_ (
    .A(_28_),
    .B(_80_),
    .Y(_45_)
);

NAND3X1 _9363_ (
    .A(\datapath.idinstr [13]),
    .B(_26_),
    .C(_80_),
    .Y(_46_)
);

NAND3X1 _9364_ (
    .A(\datapath.idinstr [14]),
    .B(_80_),
    .C(_24_),
    .Y(_47_)
);

NAND3X1 _9365_ (
    .A(_45_),
    .B(_46_),
    .C(_47_),
    .Y(_48_)
);

NAND2X1 _9366_ (
    .A(_44_),
    .B(_48_),
    .Y(_49_)
);

NAND2X1 _9367_ (
    .A(_42_),
    .B(_49_),
    .Y(_3_[1])
);

NOR2X1 _9368_ (
    .A(_27_),
    .B(_31_),
    .Y(_50_)
);

AOI21X1 _9369_ (
    .A(_33_),
    .B(\datapath.idinstr [14]),
    .C(_50_),
    .Y(_51_)
);

NAND2X1 _9370_ (
    .A(_51_),
    .B(_42_),
    .Y(_3_[2])
);

INVX1 _9371_ (
    .A(\datapath.idinstr [12]),
    .Y(_52_)
);

NAND2X1 _9372_ (
    .A(\datapath.idinstr [14]),
    .B(_21_),
    .Y(_53_)
);

OAI21X1 _9373_ (
    .A(_52_),
    .B(_53_),
    .C(_22_),
    .Y(_54_)
);

NAND3X1 _9374_ (
    .A(\datapath.idinstr [30]),
    .B(_54_),
    .C(_33_),
    .Y(_55_)
);

NAND2X1 _9375_ (
    .A(\datapath.idinstr [13]),
    .B(_52_),
    .Y(_56_)
);

AOI22X1 _9376_ (
    .A(_80_),
    .B(_24_),
    .C(_56_),
    .D(_50_),
    .Y(_57_)
);

NAND3X1 _9377_ (
    .A(_55_),
    .B(_57_),
    .C(_42_),
    .Y(_3_[3])
);

OAI21X1 _9378_ (
    .A(_81_),
    .B(_39_),
    .C(_80_),
    .Y(_58_)
);

NAND2X1 _9379_ (
    .A(\datapath.idinstr [2]),
    .B(\datapath.idinstr [3]),
    .Y(_59_)
);

NOR2X1 _9380_ (
    .A(_79_),
    .B(_59_),
    .Y(_60_)
);

AOI22X1 _9381_ (
    .A(_80_),
    .B(_28_),
    .C(_24_),
    .D(_60_),
    .Y(_61_)
);

NAND3X1 _9382_ (
    .A(_61_),
    .B(_38_),
    .C(_58_),
    .Y(_62_)
);

NAND3X1 _9383_ (
    .A(_4_),
    .B(_45_),
    .C(_62_),
    .Y(\controlunit.imm_sel [0])
);

NAND2X1 _9384_ (
    .A(_25_),
    .B(_62_),
    .Y(\controlunit.imm_sel [1])
);

INVX4 _9385_ (
    .A(_61_),
    .Y(\controlunit.imm_sel [2])
);

OAI21X1 _9386_ (
    .A(\datapath.idinstr [4]),
    .B(\datapath.idinstr [6]),
    .C(\datapath.idinstr [5]),
    .Y(_63_)
);

NOR2X1 _9387_ (
    .A(_63_),
    .B(_31_),
    .Y(_64_)
);

OAI21X1 _9388_ (
    .A(_43_),
    .B(_45_),
    .C(_64_),
    .Y(bsel[0])
);

NOR2X1 _9389_ (
    .A(\datapath.idinstr [14]),
    .B(_45_),
    .Y(bsel[1])
);

OAI22X1 _9390_ (
    .A(_8_),
    .B(_12_),
    .C(_102_),
    .D(_99_),
    .Y(\controlunit.wb_sel [0])
);

INVX1 _9391_ (
    .A(_13_),
    .Y(\controlunit.wb_sel [1])
);

NAND2X1 _9392_ (
    .A(_29_),
    .B(_38_),
    .Y(_65_)
);

OAI21X1 _9393_ (
    .A(_24_),
    .B(_40_),
    .C(_60_),
    .Y(_66_)
);

AOI22X1 _9394_ (
    .A(_80_),
    .B(_81_),
    .C(_26_),
    .D(_37_),
    .Y(_67_)
);

NAND2X1 _9395_ (
    .A(_66_),
    .B(_67_),
    .Y(_68_)
);

INVX1 _9396_ (
    .A(\datapath.idinstr_20_bF$buf29 ),
    .Y(_69_)
);

NAND3X1 _9397_ (
    .A(\datapath.idinstr_21_bF$buf42 ),
    .B(\datapath.idinstr [29]),
    .C(_69_),
    .Y(_70_)
);

NOR2X1 _9398_ (
    .A(\datapath.idinstr [12]),
    .B(_44_),
    .Y(_71_)
);

NOR2X1 _9399_ (
    .A(\datapath.idinstr_21_bF$buf41 ),
    .B(\datapath.idinstr [29]),
    .Y(_72_)
);

INVX1 _9400_ (
    .A(_72_),
    .Y(_73_)
);

NAND3X1 _9401_ (
    .A(_73_),
    .B(_70_),
    .C(_71_),
    .Y(_74_)
);

OAI22X1 _9402_ (
    .A(_45_),
    .B(_74_),
    .C(_68_),
    .D(_65_),
    .Y(\controlunit.ill_op )
);

OAI21X1 _9403_ (
    .A(\datapath.idinstr [6]),
    .B(_31_),
    .C(_38_),
    .Y(_75_)
);

NOR2X1 _9404_ (
    .A(_50_),
    .B(_75_),
    .Y(asel[0])
);

NOR2X1 _9405_ (
    .A(_43_),
    .B(_45_),
    .Y(asel[1])
);

NAND2X1 _9406_ (
    .A(_72_),
    .B(_71_),
    .Y(_76_)
);

NAND2X1 _9407_ (
    .A(\datapath.idinstr_20_bF$buf28 ),
    .B(_50_),
    .Y(_77_)
);

NOR2X1 _9408_ (
    .A(_76_),
    .B(_77_),
    .Y(\controlunit.ebreak )
);

NAND2X1 _9409_ (
    .A(_69_),
    .B(_50_),
    .Y(_78_)
);

NOR2X1 _9410_ (
    .A(_76_),
    .B(_78_),
    .Y(\controlunit.ecall )
);

\$_DLATCH_P_  _9411_ (
    .D(_3_[0]),
    .E(_4_),
    .Q(alusel[0])
);

\$_DLATCH_P_  _9412_ (
    .D(_3_[1]),
    .E(_4_),
    .Q(alusel[1])
);

\$_DLATCH_P_  _9413_ (
    .D(_3_[2]),
    .E(_4_),
    .Q(alusel[2])
);

\$_DLATCH_P_  _9414_ (
    .D(_3_[3]),
    .E(_4_),
    .Q(alusel[3])
);

INVX1 _9415_ (
    .A(\datapath.programcounter.pc [0]),
    .Y(_729_)
);

NAND2X1 _9416_ (
    .A(\datapath.idpc [0]),
    .B(1'h0),
    .Y(_730_)
);

OAI21X1 _9417_ (
    .A(1'h0),
    .B(_729_),
    .C(_730_),
    .Y(\datapath._03_ [0])
);

INVX1 _9418_ (
    .A(\datapath.programcounter.pc [1]),
    .Y(_731_)
);

NAND2X1 _9419_ (
    .A(1'h0),
    .B(\datapath.idpc [1]),
    .Y(_732_)
);

OAI21X1 _9420_ (
    .A(1'h0),
    .B(_731_),
    .C(_732_),
    .Y(\datapath._03_ [1])
);

INVX1 _9421_ (
    .A(\datapath.programcounter.pc [2]),
    .Y(_733_)
);

NAND2X1 _9422_ (
    .A(1'h0),
    .B(\datapath.idpc [2]),
    .Y(_734_)
);

OAI21X1 _9423_ (
    .A(1'h0),
    .B(_733_),
    .C(_734_),
    .Y(\datapath._03_ [2])
);

INVX1 _9424_ (
    .A(\datapath.programcounter.pc [3]),
    .Y(_735_)
);

NAND2X1 _9425_ (
    .A(1'h0),
    .B(\datapath.idpc [3]),
    .Y(_736_)
);

OAI21X1 _9426_ (
    .A(1'h0),
    .B(_735_),
    .C(_736_),
    .Y(\datapath._03_ [3])
);

INVX1 _9427_ (
    .A(\datapath.programcounter.pc [4]),
    .Y(_737_)
);

NAND2X1 _9428_ (
    .A(1'h0),
    .B(\datapath.idpc [4]),
    .Y(_738_)
);

OAI21X1 _9429_ (
    .A(1'h0),
    .B(_737_),
    .C(_738_),
    .Y(\datapath._03_ [4])
);

INVX1 _9430_ (
    .A(\datapath.programcounter.pc [5]),
    .Y(_739_)
);

NAND2X1 _9431_ (
    .A(1'h0),
    .B(\datapath.idpc [5]),
    .Y(_740_)
);

OAI21X1 _9432_ (
    .A(1'h0),
    .B(_739_),
    .C(_740_),
    .Y(\datapath._03_ [5])
);

INVX1 _9433_ (
    .A(\datapath.programcounter.pc [6]),
    .Y(_741_)
);

NAND2X1 _9434_ (
    .A(1'h0),
    .B(\datapath.idpc [6]),
    .Y(_742_)
);

OAI21X1 _9435_ (
    .A(1'h0),
    .B(_741_),
    .C(_742_),
    .Y(\datapath._03_ [6])
);

INVX1 _9436_ (
    .A(\datapath.programcounter.pc [7]),
    .Y(_743_)
);

NAND2X1 _9437_ (
    .A(1'h0),
    .B(\datapath.idpc [7]),
    .Y(_744_)
);

OAI21X1 _9438_ (
    .A(1'h0),
    .B(_743_),
    .C(_744_),
    .Y(\datapath._03_ [7])
);

INVX1 _9439_ (
    .A(\datapath.programcounter.pc [8]),
    .Y(_745_)
);

NAND2X1 _9440_ (
    .A(1'h0),
    .B(\datapath.idpc [8]),
    .Y(_746_)
);

OAI21X1 _9441_ (
    .A(1'h0),
    .B(_745_),
    .C(_746_),
    .Y(\datapath._03_ [8])
);

INVX1 _9442_ (
    .A(\datapath.programcounter.pc [9]),
    .Y(_747_)
);

NAND2X1 _9443_ (
    .A(1'h0),
    .B(\datapath.idpc [9]),
    .Y(_748_)
);

OAI21X1 _9444_ (
    .A(1'h0),
    .B(_747_),
    .C(_748_),
    .Y(\datapath._03_ [9])
);

INVX1 _9445_ (
    .A(\datapath.programcounter.pc [10]),
    .Y(_749_)
);

NAND2X1 _9446_ (
    .A(1'h0),
    .B(\datapath.idpc [10]),
    .Y(_750_)
);

OAI21X1 _9447_ (
    .A(1'h0),
    .B(_749_),
    .C(_750_),
    .Y(\datapath._03_ [10])
);

INVX1 _9448_ (
    .A(\datapath.programcounter.pc [11]),
    .Y(_751_)
);

NAND2X1 _9449_ (
    .A(1'h0),
    .B(\datapath.idpc [11]),
    .Y(_752_)
);

OAI21X1 _9450_ (
    .A(1'h0),
    .B(_751_),
    .C(_752_),
    .Y(\datapath._03_ [11])
);

INVX1 _9451_ (
    .A(\datapath.programcounter.pc [12]),
    .Y(_753_)
);

NAND2X1 _9452_ (
    .A(1'h0),
    .B(\datapath.idpc [12]),
    .Y(_754_)
);

OAI21X1 _9453_ (
    .A(1'h0),
    .B(_753_),
    .C(_754_),
    .Y(\datapath._03_ [12])
);

INVX1 _9454_ (
    .A(\datapath.programcounter.pc [13]),
    .Y(_755_)
);

NAND2X1 _9455_ (
    .A(1'h0),
    .B(\datapath.idpc [13]),
    .Y(_756_)
);

OAI21X1 _9456_ (
    .A(1'h0),
    .B(_755_),
    .C(_756_),
    .Y(\datapath._03_ [13])
);

INVX1 _9457_ (
    .A(\datapath.programcounter.pc [14]),
    .Y(_757_)
);

NAND2X1 _9458_ (
    .A(1'h0),
    .B(\datapath.idpc [14]),
    .Y(_758_)
);

OAI21X1 _9459_ (
    .A(1'h0),
    .B(_757_),
    .C(_758_),
    .Y(\datapath._03_ [14])
);

INVX1 _9460_ (
    .A(\datapath.programcounter.pc [15]),
    .Y(_759_)
);

NAND2X1 _9461_ (
    .A(1'h0),
    .B(\datapath.idpc [15]),
    .Y(_760_)
);

OAI21X1 _9462_ (
    .A(1'h0),
    .B(_759_),
    .C(_760_),
    .Y(\datapath._03_ [15])
);

INVX1 _9463_ (
    .A(\datapath.programcounter.pc [16]),
    .Y(_761_)
);

NAND2X1 _9464_ (
    .A(1'h0),
    .B(\datapath.idpc [16]),
    .Y(_762_)
);

OAI21X1 _9465_ (
    .A(1'h0),
    .B(_761_),
    .C(_762_),
    .Y(\datapath._03_ [16])
);

INVX1 _9466_ (
    .A(\datapath.programcounter.pc [17]),
    .Y(_763_)
);

NAND2X1 _9467_ (
    .A(1'h0),
    .B(\datapath.idpc [17]),
    .Y(_764_)
);

OAI21X1 _9468_ (
    .A(1'h0),
    .B(_763_),
    .C(_764_),
    .Y(\datapath._03_ [17])
);

INVX1 _9469_ (
    .A(\datapath.programcounter.pc [18]),
    .Y(_765_)
);

NAND2X1 _9470_ (
    .A(1'h0),
    .B(\datapath.idpc [18]),
    .Y(_766_)
);

OAI21X1 _9471_ (
    .A(1'h0),
    .B(_765_),
    .C(_766_),
    .Y(\datapath._03_ [18])
);

INVX1 _9472_ (
    .A(\datapath.programcounter.pc [19]),
    .Y(_767_)
);

NAND2X1 _9473_ (
    .A(1'h0),
    .B(\datapath.idpc [19]),
    .Y(_768_)
);

OAI21X1 _9474_ (
    .A(1'h0),
    .B(_767_),
    .C(_768_),
    .Y(\datapath._03_ [19])
);

INVX1 _9475_ (
    .A(\datapath.programcounter.pc [20]),
    .Y(_769_)
);

NAND2X1 _9476_ (
    .A(1'h0),
    .B(\datapath.idpc [20]),
    .Y(_770_)
);

OAI21X1 _9477_ (
    .A(1'h0),
    .B(_769_),
    .C(_770_),
    .Y(\datapath._03_ [20])
);

INVX1 _9478_ (
    .A(\datapath.programcounter.pc [21]),
    .Y(_771_)
);

NAND2X1 _9479_ (
    .A(1'h0),
    .B(\datapath.idpc [21]),
    .Y(_772_)
);

OAI21X1 _9480_ (
    .A(1'h0),
    .B(_771_),
    .C(_772_),
    .Y(\datapath._03_ [21])
);

INVX1 _9481_ (
    .A(\datapath.programcounter.pc [22]),
    .Y(_773_)
);

NAND2X1 _9482_ (
    .A(1'h0),
    .B(\datapath.idpc [22]),
    .Y(_774_)
);

OAI21X1 _9483_ (
    .A(1'h0),
    .B(_773_),
    .C(_774_),
    .Y(\datapath._03_ [22])
);

INVX1 _9484_ (
    .A(\datapath.programcounter.pc [23]),
    .Y(_775_)
);

NAND2X1 _9485_ (
    .A(1'h0),
    .B(\datapath.idpc [23]),
    .Y(_776_)
);

OAI21X1 _9486_ (
    .A(1'h0),
    .B(_775_),
    .C(_776_),
    .Y(\datapath._03_ [23])
);

INVX1 _9487_ (
    .A(\datapath.programcounter.pc [24]),
    .Y(_777_)
);

NAND2X1 _9488_ (
    .A(1'h0),
    .B(\datapath.idpc [24]),
    .Y(_778_)
);

OAI21X1 _9489_ (
    .A(1'h0),
    .B(_777_),
    .C(_778_),
    .Y(\datapath._03_ [24])
);

INVX1 _9490_ (
    .A(\datapath.programcounter.pc [25]),
    .Y(_779_)
);

NAND2X1 _9491_ (
    .A(1'h0),
    .B(\datapath.idpc [25]),
    .Y(_780_)
);

OAI21X1 _9492_ (
    .A(1'h0),
    .B(_779_),
    .C(_780_),
    .Y(\datapath._03_ [25])
);

INVX1 _9493_ (
    .A(\datapath.programcounter.pc [26]),
    .Y(_781_)
);

NAND2X1 _9494_ (
    .A(1'h0),
    .B(\datapath.idpc [26]),
    .Y(_782_)
);

OAI21X1 _9495_ (
    .A(1'h0),
    .B(_781_),
    .C(_782_),
    .Y(\datapath._03_ [26])
);

INVX1 _9496_ (
    .A(\datapath.programcounter.pc [27]),
    .Y(_783_)
);

NAND2X1 _9497_ (
    .A(1'h0),
    .B(\datapath.idpc [27]),
    .Y(_784_)
);

OAI21X1 _9498_ (
    .A(1'h0),
    .B(_783_),
    .C(_784_),
    .Y(\datapath._03_ [27])
);

INVX1 _9499_ (
    .A(\datapath.programcounter.pc [28]),
    .Y(_785_)
);

NAND2X1 _9500_ (
    .A(1'h0),
    .B(\datapath.idpc [28]),
    .Y(_786_)
);

OAI21X1 _9501_ (
    .A(1'h0),
    .B(_785_),
    .C(_786_),
    .Y(\datapath._03_ [28])
);

INVX1 _9502_ (
    .A(\datapath.programcounter.pc [29]),
    .Y(_787_)
);

NAND2X1 _9503_ (
    .A(1'h0),
    .B(\datapath.idpc [29]),
    .Y(_788_)
);

OAI21X1 _9504_ (
    .A(1'h0),
    .B(_787_),
    .C(_788_),
    .Y(\datapath._03_ [29])
);

INVX1 _9505_ (
    .A(\datapath.programcounter.pc [30]),
    .Y(_789_)
);

NAND2X1 _9506_ (
    .A(1'h0),
    .B(\datapath.idpc [30]),
    .Y(_790_)
);

OAI21X1 _9507_ (
    .A(1'h0),
    .B(_789_),
    .C(_790_),
    .Y(\datapath._03_ [30])
);

INVX1 _9508_ (
    .A(\datapath.programcounter.pc [31]),
    .Y(_791_)
);

NAND2X1 _9509_ (
    .A(1'h0),
    .B(\datapath.idpc [31]),
    .Y(_792_)
);

OAI21X1 _9510_ (
    .A(1'h0),
    .B(_791_),
    .C(_792_),
    .Y(\datapath._03_ [31])
);

INVX1 _9511_ (
    .A(\datapath.programcounter.pc [0]),
    .Y(_793_)
);

NAND2X1 _9512_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [0]),
    .Y(_794_)
);

OAI21X1 _9513_ (
    .A(1'h0),
    .B(_793_),
    .C(_794_),
    .Y(\datapath._04_ [0])
);

INVX1 _9514_ (
    .A(\datapath.programcounter.pc [1]),
    .Y(_795_)
);

NAND2X1 _9515_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [1]),
    .Y(_796_)
);

OAI21X1 _9516_ (
    .A(1'h0),
    .B(_795_),
    .C(_796_),
    .Y(\datapath._04_ [1])
);

INVX1 _9517_ (
    .A(\datapath.nextpc [2]),
    .Y(_797_)
);

NAND2X1 _9518_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [2]),
    .Y(_798_)
);

OAI21X1 _9519_ (
    .A(1'h0),
    .B(_797_),
    .C(_798_),
    .Y(\datapath._04_ [2])
);

INVX1 _9520_ (
    .A(\datapath.nextpc [3]),
    .Y(_799_)
);

NAND2X1 _9521_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [3]),
    .Y(_800_)
);

OAI21X1 _9522_ (
    .A(1'h0),
    .B(_799_),
    .C(_800_),
    .Y(\datapath._04_ [3])
);

INVX1 _9523_ (
    .A(\datapath.nextpc [4]),
    .Y(_801_)
);

NAND2X1 _9524_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [4]),
    .Y(_802_)
);

OAI21X1 _9525_ (
    .A(1'h0),
    .B(_801_),
    .C(_802_),
    .Y(\datapath._04_ [4])
);

INVX1 _9526_ (
    .A(\datapath.nextpc [5]),
    .Y(_803_)
);

NAND2X1 _9527_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [5]),
    .Y(_804_)
);

OAI21X1 _9528_ (
    .A(1'h0),
    .B(_803_),
    .C(_804_),
    .Y(\datapath._04_ [5])
);

INVX1 _9529_ (
    .A(\datapath.nextpc [6]),
    .Y(_805_)
);

NAND2X1 _9530_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [6]),
    .Y(_806_)
);

OAI21X1 _9531_ (
    .A(1'h0),
    .B(_805_),
    .C(_806_),
    .Y(\datapath._04_ [6])
);

INVX1 _9532_ (
    .A(\datapath.nextpc [7]),
    .Y(_807_)
);

NAND2X1 _9533_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [7]),
    .Y(_808_)
);

OAI21X1 _9534_ (
    .A(1'h0),
    .B(_807_),
    .C(_808_),
    .Y(\datapath._04_ [7])
);

INVX1 _9535_ (
    .A(\datapath.nextpc [8]),
    .Y(_809_)
);

NAND2X1 _9536_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [8]),
    .Y(_810_)
);

OAI21X1 _9537_ (
    .A(1'h0),
    .B(_809_),
    .C(_810_),
    .Y(\datapath._04_ [8])
);

INVX1 _9538_ (
    .A(\datapath.nextpc [9]),
    .Y(_811_)
);

NAND2X1 _9539_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [9]),
    .Y(_812_)
);

OAI21X1 _9540_ (
    .A(1'h0),
    .B(_811_),
    .C(_812_),
    .Y(\datapath._04_ [9])
);

INVX1 _9541_ (
    .A(\datapath.nextpc [10]),
    .Y(_813_)
);

NAND2X1 _9542_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [10]),
    .Y(_814_)
);

OAI21X1 _9543_ (
    .A(1'h0),
    .B(_813_),
    .C(_814_),
    .Y(\datapath._04_ [10])
);

INVX1 _9544_ (
    .A(\datapath.nextpc [11]),
    .Y(_815_)
);

NAND2X1 _9545_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [11]),
    .Y(_816_)
);

OAI21X1 _9546_ (
    .A(1'h0),
    .B(_815_),
    .C(_816_),
    .Y(\datapath._04_ [11])
);

INVX1 _9547_ (
    .A(\datapath.nextpc [12]),
    .Y(_817_)
);

NAND2X1 _9548_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [12]),
    .Y(_818_)
);

OAI21X1 _9549_ (
    .A(1'h0),
    .B(_817_),
    .C(_818_),
    .Y(\datapath._04_ [12])
);

INVX1 _9550_ (
    .A(\datapath.nextpc [13]),
    .Y(_819_)
);

NAND2X1 _9551_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [13]),
    .Y(_820_)
);

OAI21X1 _9552_ (
    .A(1'h0),
    .B(_819_),
    .C(_820_),
    .Y(\datapath._04_ [13])
);

INVX1 _9553_ (
    .A(\datapath.nextpc [14]),
    .Y(_821_)
);

NAND2X1 _9554_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [14]),
    .Y(_822_)
);

OAI21X1 _9555_ (
    .A(1'h0),
    .B(_821_),
    .C(_822_),
    .Y(\datapath._04_ [14])
);

INVX1 _9556_ (
    .A(\datapath.nextpc [15]),
    .Y(_823_)
);

NAND2X1 _9557_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [15]),
    .Y(_824_)
);

OAI21X1 _9558_ (
    .A(1'h0),
    .B(_823_),
    .C(_824_),
    .Y(\datapath._04_ [15])
);

INVX1 _9559_ (
    .A(\datapath.nextpc [16]),
    .Y(_825_)
);

NAND2X1 _9560_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [16]),
    .Y(_826_)
);

OAI21X1 _9561_ (
    .A(1'h0),
    .B(_825_),
    .C(_826_),
    .Y(\datapath._04_ [16])
);

INVX1 _9562_ (
    .A(\datapath.nextpc [17]),
    .Y(_827_)
);

NAND2X1 _9563_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [17]),
    .Y(_828_)
);

OAI21X1 _9564_ (
    .A(1'h0),
    .B(_827_),
    .C(_828_),
    .Y(\datapath._04_ [17])
);

INVX1 _9565_ (
    .A(\datapath.nextpc [18]),
    .Y(_829_)
);

NAND2X1 _9566_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [18]),
    .Y(_830_)
);

OAI21X1 _9567_ (
    .A(1'h0),
    .B(_829_),
    .C(_830_),
    .Y(\datapath._04_ [18])
);

INVX1 _9568_ (
    .A(\datapath.nextpc [19]),
    .Y(_831_)
);

NAND2X1 _9569_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [19]),
    .Y(_832_)
);

OAI21X1 _9570_ (
    .A(1'h0),
    .B(_831_),
    .C(_832_),
    .Y(\datapath._04_ [19])
);

INVX1 _9571_ (
    .A(\datapath.nextpc [20]),
    .Y(_833_)
);

NAND2X1 _9572_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [20]),
    .Y(_834_)
);

OAI21X1 _9573_ (
    .A(1'h0),
    .B(_833_),
    .C(_834_),
    .Y(\datapath._04_ [20])
);

INVX1 _9574_ (
    .A(\datapath.nextpc [21]),
    .Y(_835_)
);

NAND2X1 _9575_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [21]),
    .Y(_836_)
);

OAI21X1 _9576_ (
    .A(1'h0),
    .B(_835_),
    .C(_836_),
    .Y(\datapath._04_ [21])
);

INVX1 _9577_ (
    .A(\datapath.nextpc [22]),
    .Y(_837_)
);

NAND2X1 _9578_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [22]),
    .Y(_838_)
);

OAI21X1 _9579_ (
    .A(1'h0),
    .B(_837_),
    .C(_838_),
    .Y(\datapath._04_ [22])
);

INVX1 _9580_ (
    .A(\datapath.nextpc [23]),
    .Y(_839_)
);

NAND2X1 _9581_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [23]),
    .Y(_840_)
);

OAI21X1 _9582_ (
    .A(1'h0),
    .B(_839_),
    .C(_840_),
    .Y(\datapath._04_ [23])
);

INVX1 _9583_ (
    .A(\datapath.nextpc [24]),
    .Y(_841_)
);

NAND2X1 _9584_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [24]),
    .Y(_842_)
);

OAI21X1 _9585_ (
    .A(1'h0),
    .B(_841_),
    .C(_842_),
    .Y(\datapath._04_ [24])
);

INVX1 _9586_ (
    .A(\datapath.nextpc [25]),
    .Y(_843_)
);

NAND2X1 _9587_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [25]),
    .Y(_844_)
);

OAI21X1 _9588_ (
    .A(1'h0),
    .B(_843_),
    .C(_844_),
    .Y(\datapath._04_ [25])
);

INVX1 _9589_ (
    .A(\datapath.nextpc [26]),
    .Y(_845_)
);

NAND2X1 _9590_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [26]),
    .Y(_846_)
);

OAI21X1 _9591_ (
    .A(1'h0),
    .B(_845_),
    .C(_846_),
    .Y(\datapath._04_ [26])
);

INVX1 _9592_ (
    .A(\datapath.nextpc [27]),
    .Y(_847_)
);

NAND2X1 _9593_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [27]),
    .Y(_848_)
);

OAI21X1 _9594_ (
    .A(1'h0),
    .B(_847_),
    .C(_848_),
    .Y(\datapath._04_ [27])
);

INVX1 _9595_ (
    .A(\datapath.nextpc [28]),
    .Y(_849_)
);

NAND2X1 _9596_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [28]),
    .Y(_850_)
);

OAI21X1 _9597_ (
    .A(1'h0),
    .B(_849_),
    .C(_850_),
    .Y(\datapath._04_ [28])
);

INVX1 _9598_ (
    .A(\datapath.nextpc [29]),
    .Y(_851_)
);

NAND2X1 _9599_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [29]),
    .Y(_852_)
);

OAI21X1 _9600_ (
    .A(1'h0),
    .B(_851_),
    .C(_852_),
    .Y(\datapath._04_ [29])
);

INVX1 _9601_ (
    .A(\datapath.nextpc [30]),
    .Y(_853_)
);

NAND2X1 _9602_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [30]),
    .Y(_854_)
);

OAI21X1 _9603_ (
    .A(1'h0),
    .B(_853_),
    .C(_854_),
    .Y(\datapath._04_ [30])
);

INVX1 _9604_ (
    .A(\datapath.nextpc [31]),
    .Y(_855_)
);

NAND2X1 _9605_ (
    .A(1'h0),
    .B(\datapath.idpc_4 [31]),
    .Y(_856_)
);

OAI21X1 _9606_ (
    .A(1'h0),
    .B(_855_),
    .C(_856_),
    .Y(\datapath._04_ [31])
);

INVX1 _9607_ (
    .A(IMEM_DATA[0]),
    .Y(_857_)
);

NAND2X1 _9608_ (
    .A(1'h0),
    .B(\datapath.idinstr [0]),
    .Y(_858_)
);

OAI21X1 _9609_ (
    .A(1'h0),
    .B(_857_),
    .C(_858_),
    .Y(\datapath._05_ [0])
);

INVX1 _9610_ (
    .A(IMEM_DATA[1]),
    .Y(_859_)
);

NAND2X1 _9611_ (
    .A(1'h0),
    .B(\datapath.idinstr [1]),
    .Y(_860_)
);

OAI21X1 _9612_ (
    .A(1'h0),
    .B(_859_),
    .C(_860_),
    .Y(\datapath._05_ [1])
);

INVX1 _9613_ (
    .A(IMEM_DATA[2]),
    .Y(_861_)
);

NAND2X1 _9614_ (
    .A(1'h0),
    .B(\datapath.idinstr [2]),
    .Y(_862_)
);

OAI21X1 _9615_ (
    .A(1'h0),
    .B(_861_),
    .C(_862_),
    .Y(\datapath._05_ [2])
);

INVX1 _9616_ (
    .A(IMEM_DATA[3]),
    .Y(_863_)
);

NAND2X1 _9617_ (
    .A(1'h0),
    .B(\datapath.idinstr [3]),
    .Y(_864_)
);

OAI21X1 _9618_ (
    .A(1'h0),
    .B(_863_),
    .C(_864_),
    .Y(\datapath._05_ [3])
);

INVX1 _9619_ (
    .A(IMEM_DATA[4]),
    .Y(_865_)
);

NAND2X1 _9620_ (
    .A(1'h0),
    .B(\datapath.idinstr [4]),
    .Y(_866_)
);

OAI21X1 _9621_ (
    .A(1'h0),
    .B(_865_),
    .C(_866_),
    .Y(\datapath._05_ [4])
);

INVX1 _9622_ (
    .A(IMEM_DATA[5]),
    .Y(_867_)
);

NAND2X1 _9623_ (
    .A(1'h0),
    .B(\datapath.idinstr [5]),
    .Y(_868_)
);

OAI21X1 _9624_ (
    .A(1'h0),
    .B(_867_),
    .C(_868_),
    .Y(\datapath._05_ [5])
);

INVX1 _9625_ (
    .A(IMEM_DATA[6]),
    .Y(_869_)
);

NAND2X1 _9626_ (
    .A(1'h0),
    .B(\datapath.idinstr [6]),
    .Y(_870_)
);

OAI21X1 _9627_ (
    .A(1'h0),
    .B(_869_),
    .C(_870_),
    .Y(\datapath._05_ [6])
);

INVX1 _9628_ (
    .A(IMEM_DATA[7]),
    .Y(_871_)
);

NAND2X1 _9629_ (
    .A(1'h0),
    .B(\datapath.idinstr [7]),
    .Y(_872_)
);

OAI21X1 _9630_ (
    .A(1'h0),
    .B(_871_),
    .C(_872_),
    .Y(\datapath._05_ [7])
);

INVX1 _9631_ (
    .A(IMEM_DATA[8]),
    .Y(_105_)
);

NAND2X1 _9632_ (
    .A(1'h0),
    .B(\datapath.idinstr [8]),
    .Y(_106_)
);

OAI21X1 _9633_ (
    .A(1'h0),
    .B(_105_),
    .C(_106_),
    .Y(\datapath._05_ [8])
);

INVX1 _9634_ (
    .A(IMEM_DATA[9]),
    .Y(_107_)
);

NAND2X1 _9635_ (
    .A(1'h0),
    .B(\datapath.idinstr [9]),
    .Y(_108_)
);

OAI21X1 _9636_ (
    .A(1'h0),
    .B(_107_),
    .C(_108_),
    .Y(\datapath._05_ [9])
);

INVX1 _9637_ (
    .A(IMEM_DATA[10]),
    .Y(_109_)
);

NAND2X1 _9638_ (
    .A(1'h0),
    .B(\datapath.idinstr [10]),
    .Y(_110_)
);

OAI21X1 _9639_ (
    .A(1'h0),
    .B(_109_),
    .C(_110_),
    .Y(\datapath._05_ [10])
);

INVX1 _9640_ (
    .A(IMEM_DATA[11]),
    .Y(_111_)
);

NAND2X1 _9641_ (
    .A(1'h0),
    .B(\datapath.idinstr [11]),
    .Y(_112_)
);

OAI21X1 _9642_ (
    .A(1'h0),
    .B(_111_),
    .C(_112_),
    .Y(\datapath._05_ [11])
);

INVX1 _9643_ (
    .A(IMEM_DATA[12]),
    .Y(_113_)
);

NAND2X1 _9644_ (
    .A(1'h0),
    .B(\datapath.idinstr [12]),
    .Y(_114_)
);

OAI21X1 _9645_ (
    .A(1'h0),
    .B(_113_),
    .C(_114_),
    .Y(\datapath._05_ [12])
);

INVX1 _9646_ (
    .A(IMEM_DATA[13]),
    .Y(_115_)
);

NAND2X1 _9647_ (
    .A(1'h0),
    .B(\datapath.idinstr [13]),
    .Y(_116_)
);

OAI21X1 _9648_ (
    .A(1'h0),
    .B(_115_),
    .C(_116_),
    .Y(\datapath._05_ [13])
);

INVX1 _9649_ (
    .A(IMEM_DATA[14]),
    .Y(_117_)
);

NAND2X1 _9650_ (
    .A(1'h0),
    .B(\datapath.idinstr [14]),
    .Y(_118_)
);

OAI21X1 _9651_ (
    .A(1'h0),
    .B(_117_),
    .C(_118_),
    .Y(\datapath._05_ [14])
);

INVX1 _9652_ (
    .A(IMEM_DATA[15]),
    .Y(_119_)
);

NAND2X1 _9653_ (
    .A(1'h0),
    .B(\datapath.idinstr_15_bF$buf24 ),
    .Y(_120_)
);

OAI21X1 _9654_ (
    .A(1'h0),
    .B(_119_),
    .C(_120_),
    .Y(\datapath._05_ [15])
);

INVX1 _9655_ (
    .A(IMEM_DATA[16]),
    .Y(_121_)
);

NAND2X1 _9656_ (
    .A(1'h0),
    .B(\datapath.idinstr_16_bF$buf39 ),
    .Y(_122_)
);

OAI21X1 _9657_ (
    .A(1'h0),
    .B(_121_),
    .C(_122_),
    .Y(\datapath._05_ [16])
);

INVX1 _9658_ (
    .A(IMEM_DATA[17]),
    .Y(_123_)
);

NAND2X1 _9659_ (
    .A(1'h0),
    .B(\datapath.idinstr_17_bF$buf5 ),
    .Y(_124_)
);

OAI21X1 _9660_ (
    .A(1'h0),
    .B(_123_),
    .C(_124_),
    .Y(\datapath._05_ [17])
);

INVX1 _9661_ (
    .A(IMEM_DATA[18]),
    .Y(_125_)
);

NAND2X1 _9662_ (
    .A(1'h0),
    .B(\datapath.idinstr_18_bF$buf2 ),
    .Y(_126_)
);

OAI21X1 _9663_ (
    .A(1'h0),
    .B(_125_),
    .C(_126_),
    .Y(\datapath._05_ [18])
);

INVX1 _9664_ (
    .A(IMEM_DATA[19]),
    .Y(_127_)
);

NAND2X1 _9665_ (
    .A(1'h0),
    .B(\datapath.idinstr_19_bF$buf4 ),
    .Y(_128_)
);

OAI21X1 _9666_ (
    .A(1'h0),
    .B(_127_),
    .C(_128_),
    .Y(\datapath._05_ [19])
);

INVX1 _9667_ (
    .A(IMEM_DATA[20]),
    .Y(_129_)
);

NAND2X1 _9668_ (
    .A(1'h0),
    .B(\datapath.idinstr_20_bF$buf27 ),
    .Y(_130_)
);

OAI21X1 _9669_ (
    .A(1'h0),
    .B(_129_),
    .C(_130_),
    .Y(\datapath._05_ [20])
);

INVX1 _9670_ (
    .A(IMEM_DATA[21]),
    .Y(_131_)
);

NAND2X1 _9671_ (
    .A(1'h0),
    .B(\datapath.idinstr_21_bF$buf40 ),
    .Y(_132_)
);

OAI21X1 _9672_ (
    .A(1'h0),
    .B(_131_),
    .C(_132_),
    .Y(\datapath._05_ [21])
);

INVX1 _9673_ (
    .A(IMEM_DATA[22]),
    .Y(_133_)
);

NAND2X1 _9674_ (
    .A(1'h0),
    .B(\datapath.idinstr_22_bF$buf15 ),
    .Y(_134_)
);

OAI21X1 _9675_ (
    .A(1'h0),
    .B(_133_),
    .C(_134_),
    .Y(\datapath._05_ [22])
);

INVX1 _9676_ (
    .A(IMEM_DATA[23]),
    .Y(_135_)
);

NAND2X1 _9677_ (
    .A(1'h0),
    .B(\datapath.idinstr_23_bF$buf3 ),
    .Y(_136_)
);

OAI21X1 _9678_ (
    .A(1'h0),
    .B(_135_),
    .C(_136_),
    .Y(\datapath._05_ [23])
);

INVX1 _9679_ (
    .A(IMEM_DATA[24]),
    .Y(_137_)
);

NAND2X1 _9680_ (
    .A(1'h0),
    .B(\datapath.idinstr_24_bF$buf3 ),
    .Y(_138_)
);

OAI21X1 _9681_ (
    .A(1'h0),
    .B(_137_),
    .C(_138_),
    .Y(\datapath._05_ [24])
);

INVX1 _9682_ (
    .A(IMEM_DATA[25]),
    .Y(_139_)
);

NAND2X1 _9683_ (
    .A(1'h0),
    .B(\datapath.idinstr [25]),
    .Y(_140_)
);

OAI21X1 _9684_ (
    .A(1'h0),
    .B(_139_),
    .C(_140_),
    .Y(\datapath._05_ [25])
);

INVX1 _9685_ (
    .A(IMEM_DATA[26]),
    .Y(_141_)
);

NAND2X1 _9686_ (
    .A(1'h0),
    .B(\datapath.idinstr [26]),
    .Y(_142_)
);

OAI21X1 _9687_ (
    .A(1'h0),
    .B(_141_),
    .C(_142_),
    .Y(\datapath._05_ [26])
);

INVX1 _9688_ (
    .A(IMEM_DATA[27]),
    .Y(_143_)
);

NAND2X1 _9689_ (
    .A(1'h0),
    .B(\datapath.idinstr [27]),
    .Y(_144_)
);

OAI21X1 _9690_ (
    .A(1'h0),
    .B(_143_),
    .C(_144_),
    .Y(\datapath._05_ [27])
);

INVX1 _9691_ (
    .A(IMEM_DATA[28]),
    .Y(_145_)
);

NAND2X1 _9692_ (
    .A(1'h0),
    .B(\datapath.idinstr [28]),
    .Y(_146_)
);

OAI21X1 _9693_ (
    .A(1'h0),
    .B(_145_),
    .C(_146_),
    .Y(\datapath._05_ [28])
);

INVX1 _9694_ (
    .A(IMEM_DATA[29]),
    .Y(_147_)
);

NAND2X1 _9695_ (
    .A(1'h0),
    .B(\datapath.idinstr [29]),
    .Y(_148_)
);

OAI21X1 _9696_ (
    .A(1'h0),
    .B(_147_),
    .C(_148_),
    .Y(\datapath._05_ [29])
);

INVX1 _9697_ (
    .A(IMEM_DATA[30]),
    .Y(_149_)
);

NAND2X1 _9698_ (
    .A(1'h0),
    .B(\datapath.idinstr [30]),
    .Y(_150_)
);

OAI21X1 _9699_ (
    .A(1'h0),
    .B(_149_),
    .C(_150_),
    .Y(\datapath._05_ [30])
);

INVX1 _9700_ (
    .A(IMEM_DATA[31]),
    .Y(_151_)
);

NAND2X1 _9701_ (
    .A(1'h0),
    .B(\datapath.idinstr [31]),
    .Y(_152_)
);

OAI21X1 _9702_ (
    .A(1'h0),
    .B(_151_),
    .C(_152_),
    .Y(\datapath._05_ [31])
);

INVX1 _9703_ (
    .A(\datapath.memexecptions [0]),
    .Y(_153_)
);

INVX1 _9704_ (
    .A(\datapath.meminstr [5]),
    .Y(_154_)
);

NOR2X1 _9705_ (
    .A(\datapath.meminstr [4]),
    .B(_154_),
    .Y(_155_)
);

NAND2X1 _9706_ (
    .A(\datapath.meminstr [6]),
    .B(_155_),
    .Y(_156_)
);

NAND2X1 _9707_ (
    .A(\datapath.meminstr [1]),
    .B(\datapath.meminstr [0]),
    .Y(_157_)
);

INVX1 _9708_ (
    .A(_156_),
    .Y(_158_)
);

OR2X2 _9709_ (
    .A(\datapath.meminstr [3]),
    .B(\datapath.meminstr [2]),
    .Y(_159_)
);

NOR2X1 _9710_ (
    .A(_157_),
    .B(_159_),
    .Y(_160_)
);

NAND3X1 _9711_ (
    .A(\datapath.tkbranch ),
    .B(_160_),
    .C(_158_),
    .Y(_161_)
);

NAND3X1 _9712_ (
    .A(\datapath.meminstr [3]),
    .B(\datapath.meminstr [2]),
    .C(_158_),
    .Y(_162_)
);

OAI21X1 _9713_ (
    .A(_157_),
    .B(_162_),
    .C(_161_),
    .Y(_163_)
);

OAI21X1 _9714_ (
    .A(\datapath.programcounter.jumps [1]),
    .B(\datapath.programcounter.jumps [0]),
    .C(_163_),
    .Y(_164_)
);

AND2X2 _9715_ (
    .A(_0__1_bF$buf2),
    .B(\datapath.meminstr [2]),
    .Y(_165_)
);

NOR2X1 _9716_ (
    .A(\datapath.meminstr [3]),
    .B(_157_),
    .Y(_166_)
);

NAND2X1 _9717_ (
    .A(_165_),
    .B(_166_),
    .Y(_167_)
);

OAI21X1 _9718_ (
    .A(_156_),
    .B(_167_),
    .C(_164_),
    .Y(_168_)
);

INVX1 _9719_ (
    .A(_168_),
    .Y(_169_)
);

NAND3X1 _9720_ (
    .A(_153_),
    .B(\datapath.memexecptions [2]),
    .C(_169_),
    .Y(_170_)
);

NOR2X1 _9721_ (
    .A(\datapath.memexecptions [1]),
    .B(\datapath.csr.csr_irq ),
    .Y(_171_)
);

NAND2X1 _9722_ (
    .A(_171_),
    .B(_170_),
    .Y(\datapath.csr.csr_mcause [0])
);

NOR2X1 _9723_ (
    .A(\datapath.memexecptions [0]),
    .B(\datapath.memexecptions [2]),
    .Y(_172_)
);

NAND2X1 _9724_ (
    .A(_171_),
    .B(_172_),
    .Y(_173_)
);

INVX1 _9725_ (
    .A(_173_),
    .Y(_174_)
);

NOR2X1 _9726_ (
    .A(\datapath.meminstr [4]),
    .B(\datapath.meminstr [6]),
    .Y(_175_)
);

NAND2X1 _9727_ (
    .A(_0__1_bF$buf1),
    .B(\datapath.meminstr [12]),
    .Y(_176_)
);

OAI21X1 _9728_ (
    .A(_0__1_bF$buf0),
    .B(_0__0_bF$buf0),
    .C(\datapath.meminstr [13]),
    .Y(_177_)
);

NAND2X1 _9729_ (
    .A(_176_),
    .B(_177_),
    .Y(_178_)
);

NAND3X1 _9730_ (
    .A(_175_),
    .B(_178_),
    .C(_160_),
    .Y(_179_)
);

OR2X2 _9731_ (
    .A(_179_),
    .B(_154_),
    .Y(_180_)
);

AOI22X1 _9732_ (
    .A(_174_),
    .B(_180_),
    .C(_171_),
    .D(_168_),
    .Y(\datapath.csr.csr_mcause [1])
);

NOR2X1 _9733_ (
    .A(_173_),
    .B(_168_),
    .Y(\datapath.csr.csr_mcause [2])
);

INVX1 _9734_ (
    .A(\datapath.csr.csr_irq ),
    .Y(_181_)
);

OAI21X1 _9735_ (
    .A(\datapath.memexecptions [1]),
    .B(_170_),
    .C(_181_),
    .Y(\datapath.csr.csr_mcause [3])
);

NOR2X1 _9736_ (
    .A(\controlunit.wb_sel [0]),
    .B(\controlunit.wb_sel [1]),
    .Y(_182_)
);

INVX1 _9737_ (
    .A(\controlunit.wb_sel [1]),
    .Y(_183_)
);

NOR2X1 _9738_ (
    .A(\controlunit.wb_sel [0]),
    .B(_183_),
    .Y(_184_)
);

AOI22X1 _9739_ (
    .A(\datapath.regcwb [0]),
    .B(_182__bF$buf4),
    .C(\datapath.wbpc_4 [0]),
    .D(_184__bF$buf4),
    .Y(_185_)
);

INVX1 _9740_ (
    .A(\controlunit.wb_sel [0]),
    .Y(_186_)
);

NOR2X1 _9741_ (
    .A(\controlunit.wb_sel [1]),
    .B(_186_),
    .Y(_187_)
);

NAND2X1 _9742_ (
    .A(\datapath.regloadwb [0]),
    .B(_187__bF$buf4),
    .Y(_188_)
);

NOR2X1 _9743_ (
    .A(_186_),
    .B(_183_),
    .Y(_189_)
);

NAND2X1 _9744_ (
    .A(\datapath.regcsrwb [0]),
    .B(_189__bF$buf4),
    .Y(_190_)
);

NAND3X1 _9745_ (
    .A(_188_),
    .B(_190_),
    .C(_185_),
    .Y(\datapath.rd [0])
);

AOI22X1 _9746_ (
    .A(_184__bF$buf3),
    .B(\datapath.wbpc_4 [1]),
    .C(\datapath.regcsrwb [1]),
    .D(_189__bF$buf3),
    .Y(_191_)
);

NAND2X1 _9747_ (
    .A(\datapath.regcwb [1]),
    .B(_182__bF$buf3),
    .Y(_192_)
);

NAND2X1 _9748_ (
    .A(\datapath.regloadwb [1]),
    .B(_187__bF$buf3),
    .Y(_193_)
);

NAND3X1 _9749_ (
    .A(_192_),
    .B(_193_),
    .C(_191_),
    .Y(\datapath.rd [1])
);

AOI22X1 _9750_ (
    .A(_184__bF$buf2),
    .B(\datapath.wbpc_4 [2]),
    .C(\datapath.regcsrwb [2]),
    .D(_189__bF$buf2),
    .Y(_194_)
);

NAND2X1 _9751_ (
    .A(\datapath.regcwb [2]),
    .B(_182__bF$buf2),
    .Y(_195_)
);

NAND2X1 _9752_ (
    .A(\datapath.regloadwb [2]),
    .B(_187__bF$buf2),
    .Y(_196_)
);

NAND3X1 _9753_ (
    .A(_195_),
    .B(_196_),
    .C(_194_),
    .Y(\datapath.rd [2])
);

AOI22X1 _9754_ (
    .A(_184__bF$buf1),
    .B(\datapath.wbpc_4 [3]),
    .C(\datapath.regcsrwb [3]),
    .D(_189__bF$buf1),
    .Y(_197_)
);

NAND2X1 _9755_ (
    .A(\datapath.regcwb [3]),
    .B(_182__bF$buf1),
    .Y(_198_)
);

NAND2X1 _9756_ (
    .A(\datapath.regloadwb [3]),
    .B(_187__bF$buf1),
    .Y(_199_)
);

NAND3X1 _9757_ (
    .A(_198_),
    .B(_199_),
    .C(_197_),
    .Y(\datapath.rd [3])
);

AOI22X1 _9758_ (
    .A(_184__bF$buf0),
    .B(\datapath.wbpc_4 [4]),
    .C(\datapath.regcsrwb [4]),
    .D(_189__bF$buf0),
    .Y(_200_)
);

NAND2X1 _9759_ (
    .A(\datapath.regcwb [4]),
    .B(_182__bF$buf0),
    .Y(_201_)
);

NAND2X1 _9760_ (
    .A(\datapath.regloadwb [4]),
    .B(_187__bF$buf0),
    .Y(_202_)
);

NAND3X1 _9761_ (
    .A(_201_),
    .B(_202_),
    .C(_200_),
    .Y(\datapath.rd [4])
);

AOI22X1 _9762_ (
    .A(_184__bF$buf4),
    .B(\datapath.wbpc_4 [5]),
    .C(\datapath.regcsrwb [5]),
    .D(_189__bF$buf4),
    .Y(_203_)
);

NAND2X1 _9763_ (
    .A(\datapath.regcwb [5]),
    .B(_182__bF$buf4),
    .Y(_204_)
);

NAND2X1 _9764_ (
    .A(\datapath.regloadwb [5]),
    .B(_187__bF$buf4),
    .Y(_205_)
);

NAND3X1 _9765_ (
    .A(_204_),
    .B(_205_),
    .C(_203_),
    .Y(\datapath.rd [5])
);

NAND2X1 _9766_ (
    .A(\datapath.regloadwb [6]),
    .B(_187__bF$buf3),
    .Y(_206_)
);

NAND2X1 _9767_ (
    .A(\datapath.regcsrwb [6]),
    .B(_189__bF$buf3),
    .Y(_207_)
);

AOI22X1 _9768_ (
    .A(\datapath.regcwb [6]),
    .B(_182__bF$buf3),
    .C(\datapath.wbpc_4 [6]),
    .D(_184__bF$buf3),
    .Y(_208_)
);

NAND3X1 _9769_ (
    .A(_206_),
    .B(_207_),
    .C(_208_),
    .Y(\datapath.rd [6])
);

AOI22X1 _9770_ (
    .A(_184__bF$buf2),
    .B(\datapath.wbpc_4 [7]),
    .C(\datapath.regcsrwb [7]),
    .D(_189__bF$buf2),
    .Y(_209_)
);

NAND2X1 _9771_ (
    .A(\datapath.regcwb [7]),
    .B(_182__bF$buf2),
    .Y(_210_)
);

NAND2X1 _9772_ (
    .A(\datapath.regloadwb [7]),
    .B(_187__bF$buf2),
    .Y(_211_)
);

NAND3X1 _9773_ (
    .A(_210_),
    .B(_211_),
    .C(_209_),
    .Y(\datapath.rd [7])
);

AOI22X1 _9774_ (
    .A(_184__bF$buf1),
    .B(\datapath.wbpc_4 [8]),
    .C(\datapath.regcsrwb [8]),
    .D(_189__bF$buf1),
    .Y(_212_)
);

NAND2X1 _9775_ (
    .A(\datapath.regcwb [8]),
    .B(_182__bF$buf1),
    .Y(_213_)
);

NAND2X1 _9776_ (
    .A(\datapath.regloadwb [8]),
    .B(_187__bF$buf1),
    .Y(_214_)
);

NAND3X1 _9777_ (
    .A(_213_),
    .B(_214_),
    .C(_212_),
    .Y(\datapath.rd [8])
);

AOI22X1 _9778_ (
    .A(_184__bF$buf0),
    .B(\datapath.wbpc_4 [9]),
    .C(\datapath.regcsrwb [9]),
    .D(_189__bF$buf0),
    .Y(_215_)
);

NAND2X1 _9779_ (
    .A(\datapath.regcwb [9]),
    .B(_182__bF$buf0),
    .Y(_216_)
);

NAND2X1 _9780_ (
    .A(\datapath.regloadwb [9]),
    .B(_187__bF$buf0),
    .Y(_217_)
);

NAND3X1 _9781_ (
    .A(_216_),
    .B(_217_),
    .C(_215_),
    .Y(\datapath.rd [9])
);

AOI22X1 _9782_ (
    .A(_184__bF$buf4),
    .B(\datapath.wbpc_4 [10]),
    .C(\datapath.regcsrwb [10]),
    .D(_189__bF$buf4),
    .Y(_218_)
);

NAND2X1 _9783_ (
    .A(\datapath.regcwb [10]),
    .B(_182__bF$buf4),
    .Y(_219_)
);

NAND2X1 _9784_ (
    .A(\datapath.regloadwb [10]),
    .B(_187__bF$buf4),
    .Y(_220_)
);

NAND3X1 _9785_ (
    .A(_219_),
    .B(_220_),
    .C(_218_),
    .Y(\datapath.rd [10])
);

AOI22X1 _9786_ (
    .A(_184__bF$buf3),
    .B(\datapath.wbpc_4 [11]),
    .C(\datapath.regcsrwb [11]),
    .D(_189__bF$buf3),
    .Y(_221_)
);

NAND2X1 _9787_ (
    .A(\datapath.regcwb [11]),
    .B(_182__bF$buf3),
    .Y(_222_)
);

NAND2X1 _9788_ (
    .A(\datapath.regloadwb [11]),
    .B(_187__bF$buf3),
    .Y(_223_)
);

NAND3X1 _9789_ (
    .A(_222_),
    .B(_223_),
    .C(_221_),
    .Y(\datapath.rd [11])
);

AOI22X1 _9790_ (
    .A(_184__bF$buf2),
    .B(\datapath.wbpc_4 [12]),
    .C(\datapath.regcsrwb [12]),
    .D(_189__bF$buf2),
    .Y(_224_)
);

NAND2X1 _9791_ (
    .A(\datapath.regcwb [12]),
    .B(_182__bF$buf2),
    .Y(_225_)
);

NAND2X1 _9792_ (
    .A(\datapath.regloadwb [12]),
    .B(_187__bF$buf2),
    .Y(_226_)
);

NAND3X1 _9793_ (
    .A(_225_),
    .B(_226_),
    .C(_224_),
    .Y(\datapath.rd [12])
);

AOI22X1 _9794_ (
    .A(_184__bF$buf1),
    .B(\datapath.wbpc_4 [13]),
    .C(\datapath.regcsrwb [13]),
    .D(_189__bF$buf1),
    .Y(_227_)
);

NAND2X1 _9795_ (
    .A(\datapath.regcwb [13]),
    .B(_182__bF$buf1),
    .Y(_228_)
);

NAND2X1 _9796_ (
    .A(\datapath.regloadwb [13]),
    .B(_187__bF$buf1),
    .Y(_229_)
);

NAND3X1 _9797_ (
    .A(_228_),
    .B(_229_),
    .C(_227_),
    .Y(\datapath.rd [13])
);

NAND2X1 _9798_ (
    .A(\datapath.regloadwb [14]),
    .B(_187__bF$buf0),
    .Y(_230_)
);

NAND2X1 _9799_ (
    .A(\datapath.regcsrwb [14]),
    .B(_189__bF$buf0),
    .Y(_231_)
);

AOI22X1 _9800_ (
    .A(\datapath.regcwb [14]),
    .B(_182__bF$buf0),
    .C(\datapath.wbpc_4 [14]),
    .D(_184__bF$buf0),
    .Y(_232_)
);

NAND3X1 _9801_ (
    .A(_230_),
    .B(_231_),
    .C(_232_),
    .Y(\datapath.rd [14])
);

AOI22X1 _9802_ (
    .A(_184__bF$buf4),
    .B(\datapath.wbpc_4 [15]),
    .C(\datapath.regcsrwb [15]),
    .D(_189__bF$buf4),
    .Y(_233_)
);

NAND2X1 _9803_ (
    .A(\datapath.regcwb [15]),
    .B(_182__bF$buf4),
    .Y(_234_)
);

NAND2X1 _9804_ (
    .A(\datapath.regloadwb [15]),
    .B(_187__bF$buf4),
    .Y(_235_)
);

NAND3X1 _9805_ (
    .A(_234_),
    .B(_235_),
    .C(_233_),
    .Y(\datapath.rd [15])
);

AOI22X1 _9806_ (
    .A(_184__bF$buf3),
    .B(\datapath.wbpc_4 [16]),
    .C(\datapath.regcsrwb [16]),
    .D(_189__bF$buf3),
    .Y(_236_)
);

NAND2X1 _9807_ (
    .A(\datapath.regcwb [16]),
    .B(_182__bF$buf3),
    .Y(_237_)
);

NAND2X1 _9808_ (
    .A(\datapath.regloadwb [16]),
    .B(_187__bF$buf3),
    .Y(_238_)
);

NAND3X1 _9809_ (
    .A(_237_),
    .B(_238_),
    .C(_236_),
    .Y(\datapath.rd [16])
);

AOI22X1 _9810_ (
    .A(_184__bF$buf2),
    .B(\datapath.wbpc_4 [17]),
    .C(\datapath.regcsrwb [17]),
    .D(_189__bF$buf2),
    .Y(_239_)
);

NAND2X1 _9811_ (
    .A(\datapath.regcwb [17]),
    .B(_182__bF$buf2),
    .Y(_240_)
);

NAND2X1 _9812_ (
    .A(\datapath.regloadwb [17]),
    .B(_187__bF$buf2),
    .Y(_241_)
);

NAND3X1 _9813_ (
    .A(_240_),
    .B(_241_),
    .C(_239_),
    .Y(\datapath.rd [17])
);

AOI22X1 _9814_ (
    .A(_184__bF$buf1),
    .B(\datapath.wbpc_4 [18]),
    .C(\datapath.regcsrwb [18]),
    .D(_189__bF$buf1),
    .Y(_242_)
);

NAND2X1 _9815_ (
    .A(\datapath.regcwb [18]),
    .B(_182__bF$buf1),
    .Y(_243_)
);

NAND2X1 _9816_ (
    .A(\datapath.regloadwb [18]),
    .B(_187__bF$buf1),
    .Y(_244_)
);

NAND3X1 _9817_ (
    .A(_243_),
    .B(_244_),
    .C(_242_),
    .Y(\datapath.rd [18])
);

AOI22X1 _9818_ (
    .A(_184__bF$buf0),
    .B(\datapath.wbpc_4 [19]),
    .C(\datapath.regcsrwb [19]),
    .D(_189__bF$buf0),
    .Y(_245_)
);

NAND2X1 _9819_ (
    .A(\datapath.regcwb [19]),
    .B(_182__bF$buf0),
    .Y(_246_)
);

NAND2X1 _9820_ (
    .A(\datapath.regloadwb [19]),
    .B(_187__bF$buf0),
    .Y(_247_)
);

NAND3X1 _9821_ (
    .A(_246_),
    .B(_247_),
    .C(_245_),
    .Y(\datapath.rd [19])
);

AOI22X1 _9822_ (
    .A(_184__bF$buf4),
    .B(\datapath.wbpc_4 [20]),
    .C(\datapath.regcsrwb [20]),
    .D(_189__bF$buf4),
    .Y(_248_)
);

NAND2X1 _9823_ (
    .A(\datapath.regcwb [20]),
    .B(_182__bF$buf4),
    .Y(_249_)
);

NAND2X1 _9824_ (
    .A(\datapath.regloadwb [20]),
    .B(_187__bF$buf4),
    .Y(_250_)
);

NAND3X1 _9825_ (
    .A(_249_),
    .B(_250_),
    .C(_248_),
    .Y(\datapath.rd [20])
);

AOI22X1 _9826_ (
    .A(_184__bF$buf3),
    .B(\datapath.wbpc_4 [21]),
    .C(\datapath.regcsrwb [21]),
    .D(_189__bF$buf3),
    .Y(_251_)
);

NAND2X1 _9827_ (
    .A(\datapath.regcwb [21]),
    .B(_182__bF$buf3),
    .Y(_252_)
);

NAND2X1 _9828_ (
    .A(\datapath.regloadwb [21]),
    .B(_187__bF$buf3),
    .Y(_253_)
);

NAND3X1 _9829_ (
    .A(_252_),
    .B(_253_),
    .C(_251_),
    .Y(\datapath.rd [21])
);

NAND2X1 _9830_ (
    .A(\datapath.regloadwb [22]),
    .B(_187__bF$buf2),
    .Y(_254_)
);

NAND2X1 _9831_ (
    .A(\datapath.regcsrwb [22]),
    .B(_189__bF$buf2),
    .Y(_255_)
);

AOI22X1 _9832_ (
    .A(\datapath.regcwb [22]),
    .B(_182__bF$buf2),
    .C(\datapath.wbpc_4 [22]),
    .D(_184__bF$buf2),
    .Y(_256_)
);

NAND3X1 _9833_ (
    .A(_254_),
    .B(_255_),
    .C(_256_),
    .Y(\datapath.rd [22])
);

AOI22X1 _9834_ (
    .A(_184__bF$buf1),
    .B(\datapath.wbpc_4 [23]),
    .C(\datapath.regcsrwb [23]),
    .D(_189__bF$buf1),
    .Y(_257_)
);

NAND2X1 _9835_ (
    .A(\datapath.regcwb [23]),
    .B(_182__bF$buf1),
    .Y(_258_)
);

NAND2X1 _9836_ (
    .A(\datapath.regloadwb [23]),
    .B(_187__bF$buf1),
    .Y(_259_)
);

NAND3X1 _9837_ (
    .A(_258_),
    .B(_259_),
    .C(_257_),
    .Y(\datapath.rd [23])
);

AOI22X1 _9838_ (
    .A(_184__bF$buf0),
    .B(\datapath.wbpc_4 [24]),
    .C(\datapath.regcsrwb [24]),
    .D(_189__bF$buf0),
    .Y(_260_)
);

NAND2X1 _9839_ (
    .A(\datapath.regcwb [24]),
    .B(_182__bF$buf0),
    .Y(_261_)
);

NAND2X1 _9840_ (
    .A(\datapath.regloadwb [24]),
    .B(_187__bF$buf0),
    .Y(_262_)
);

NAND3X1 _9841_ (
    .A(_261_),
    .B(_262_),
    .C(_260_),
    .Y(\datapath.rd [24])
);

AOI22X1 _9842_ (
    .A(_184__bF$buf4),
    .B(\datapath.wbpc_4 [25]),
    .C(\datapath.regcsrwb [25]),
    .D(_189__bF$buf4),
    .Y(_263_)
);

NAND2X1 _9843_ (
    .A(\datapath.regcwb [25]),
    .B(_182__bF$buf4),
    .Y(_264_)
);

NAND2X1 _9844_ (
    .A(\datapath.regloadwb [25]),
    .B(_187__bF$buf4),
    .Y(_265_)
);

NAND3X1 _9845_ (
    .A(_264_),
    .B(_265_),
    .C(_263_),
    .Y(\datapath.rd [25])
);

AOI22X1 _9846_ (
    .A(_184__bF$buf3),
    .B(\datapath.wbpc_4 [26]),
    .C(\datapath.regcsrwb [26]),
    .D(_189__bF$buf3),
    .Y(_266_)
);

NAND2X1 _9847_ (
    .A(\datapath.regcwb [26]),
    .B(_182__bF$buf3),
    .Y(_267_)
);

NAND2X1 _9848_ (
    .A(\datapath.regloadwb [26]),
    .B(_187__bF$buf3),
    .Y(_268_)
);

NAND3X1 _9849_ (
    .A(_267_),
    .B(_268_),
    .C(_266_),
    .Y(\datapath.rd [26])
);

AOI22X1 _9850_ (
    .A(_184__bF$buf2),
    .B(\datapath.wbpc_4 [27]),
    .C(\datapath.regcsrwb [27]),
    .D(_189__bF$buf2),
    .Y(_269_)
);

NAND2X1 _9851_ (
    .A(\datapath.regcwb [27]),
    .B(_182__bF$buf2),
    .Y(_270_)
);

NAND2X1 _9852_ (
    .A(\datapath.regloadwb [27]),
    .B(_187__bF$buf2),
    .Y(_271_)
);

NAND3X1 _9853_ (
    .A(_270_),
    .B(_271_),
    .C(_269_),
    .Y(\datapath.rd [27])
);

AOI22X1 _9854_ (
    .A(_184__bF$buf1),
    .B(\datapath.wbpc_4 [28]),
    .C(\datapath.regcsrwb [28]),
    .D(_189__bF$buf1),
    .Y(_272_)
);

NAND2X1 _9855_ (
    .A(\datapath.regcwb [28]),
    .B(_182__bF$buf1),
    .Y(_273_)
);

NAND2X1 _9856_ (
    .A(\datapath.regloadwb [28]),
    .B(_187__bF$buf1),
    .Y(_274_)
);

NAND3X1 _9857_ (
    .A(_273_),
    .B(_274_),
    .C(_272_),
    .Y(\datapath.rd [28])
);

AOI22X1 _9858_ (
    .A(_184__bF$buf0),
    .B(\datapath.wbpc_4 [29]),
    .C(\datapath.regcsrwb [29]),
    .D(_189__bF$buf0),
    .Y(_275_)
);

NAND2X1 _9859_ (
    .A(\datapath.regcwb [29]),
    .B(_182__bF$buf0),
    .Y(_276_)
);

NAND2X1 _9860_ (
    .A(\datapath.regloadwb [29]),
    .B(_187__bF$buf0),
    .Y(_277_)
);

NAND3X1 _9861_ (
    .A(_276_),
    .B(_277_),
    .C(_275_),
    .Y(\datapath.rd [29])
);

NAND2X1 _9862_ (
    .A(\datapath.regloadwb [30]),
    .B(_187__bF$buf4),
    .Y(_278_)
);

NAND2X1 _9863_ (
    .A(\datapath.regcsrwb [30]),
    .B(_189__bF$buf4),
    .Y(_279_)
);

AOI22X1 _9864_ (
    .A(\datapath.regcwb [30]),
    .B(_182__bF$buf4),
    .C(\datapath.wbpc_4 [30]),
    .D(_184__bF$buf4),
    .Y(_280_)
);

NAND3X1 _9865_ (
    .A(_278_),
    .B(_279_),
    .C(_280_),
    .Y(\datapath.rd [30])
);

AOI22X1 _9866_ (
    .A(_184__bF$buf3),
    .B(\datapath.wbpc_4 [31]),
    .C(\datapath.regcsrwb [31]),
    .D(_189__bF$buf3),
    .Y(_281_)
);

NAND2X1 _9867_ (
    .A(\datapath.regcwb [31]),
    .B(_182__bF$buf3),
    .Y(_282_)
);

NAND2X1 _9868_ (
    .A(\datapath.regloadwb [31]),
    .B(_187__bF$buf3),
    .Y(_283_)
);

NAND3X1 _9869_ (
    .A(_282_),
    .B(_283_),
    .C(_281_),
    .Y(\datapath.rd [31])
);

MUX2X1 _9870_ (
    .A(\datapath.regcondt ),
    .B(\datapath.regz ),
    .S(\datapath.meminstr [14]),
    .Y(_284_)
);

XNOR2X1 _9871_ (
    .A(_284_),
    .B(\datapath.meminstr [12]),
    .Y(\datapath.tkbranch )
);

INVX1 _9872_ (
    .A(bsel[1]),
    .Y(_285_)
);

AND2X2 _9873_ (
    .A(_285_),
    .B(bsel[0]),
    .Y(_286_)
);

NOR2X1 _9874_ (
    .A(bsel[0]),
    .B(_285_),
    .Y(_287_)
);

NOR2X1 _9875_ (
    .A(_287__bF$buf3),
    .B(_286__bF$buf3),
    .Y(_288_)
);

NAND2X1 _9876_ (
    .A(\datapath.registers.regb_data [0]),
    .B(_288__bF$buf3),
    .Y(_289_)
);

NAND2X1 _9877_ (
    .A(\datapath.immediatedecoder._06_ ),
    .B(_286__bF$buf2),
    .Y(_290_)
);

NAND2X1 _9878_ (
    .A(\datapath.csr.csr_data [0]),
    .B(_287__bF$buf2),
    .Y(_291_)
);

NAND3X1 _9879_ (
    .A(_290_),
    .B(_291_),
    .C(_289_),
    .Y(\datapath.muxbval [0])
);

NAND2X1 _9880_ (
    .A(\datapath.registers.regb_data [1]),
    .B(_288__bF$buf2),
    .Y(_292_)
);

NAND2X1 _9881_ (
    .A(\datapath.imm [1]),
    .B(_286__bF$buf1),
    .Y(_293_)
);

NAND2X1 _9882_ (
    .A(\datapath.csr.csr_data [1]),
    .B(_287__bF$buf1),
    .Y(_294_)
);

NAND3X1 _9883_ (
    .A(_293_),
    .B(_294_),
    .C(_292_),
    .Y(\datapath.muxbval [1])
);

NAND2X1 _9884_ (
    .A(\datapath.registers.regb_data [2]),
    .B(_288__bF$buf1),
    .Y(_295_)
);

NAND2X1 _9885_ (
    .A(\datapath.imm [2]),
    .B(_286__bF$buf0),
    .Y(_296_)
);

NAND2X1 _9886_ (
    .A(\datapath.csr.csr_data [2]),
    .B(_287__bF$buf0),
    .Y(_297_)
);

NAND3X1 _9887_ (
    .A(_296_),
    .B(_297_),
    .C(_295_),
    .Y(\datapath.muxbval [2])
);

NAND2X1 _9888_ (
    .A(\datapath.registers.regb_data [3]),
    .B(_288__bF$buf0),
    .Y(_298_)
);

NAND2X1 _9889_ (
    .A(\datapath.imm [3]),
    .B(_286__bF$buf4),
    .Y(_299_)
);

NAND2X1 _9890_ (
    .A(\datapath.csr.csr_data [3]),
    .B(_287__bF$buf4),
    .Y(_300_)
);

NAND3X1 _9891_ (
    .A(_299_),
    .B(_300_),
    .C(_298_),
    .Y(\datapath.muxbval [3])
);

NAND2X1 _9892_ (
    .A(\datapath.registers.regb_data [4]),
    .B(_288__bF$buf4),
    .Y(_301_)
);

NAND2X1 _9893_ (
    .A(\datapath.imm [4]),
    .B(_286__bF$buf3),
    .Y(_302_)
);

NAND2X1 _9894_ (
    .A(\datapath.csr.csr_data [4]),
    .B(_287__bF$buf3),
    .Y(_303_)
);

NAND3X1 _9895_ (
    .A(_302_),
    .B(_303_),
    .C(_301_),
    .Y(\datapath.muxbval [4])
);

NAND2X1 _9896_ (
    .A(\datapath.registers.regb_data [5]),
    .B(_288__bF$buf3),
    .Y(_304_)
);

NAND2X1 _9897_ (
    .A(\datapath.imm [5]),
    .B(_286__bF$buf2),
    .Y(_305_)
);

NAND2X1 _9898_ (
    .A(\datapath.csr.csr_data [5]),
    .B(_287__bF$buf2),
    .Y(_306_)
);

NAND3X1 _9899_ (
    .A(_305_),
    .B(_306_),
    .C(_304_),
    .Y(\datapath.muxbval [5])
);

NAND2X1 _9900_ (
    .A(\datapath.registers.regb_data [6]),
    .B(_288__bF$buf2),
    .Y(_307_)
);

NAND2X1 _9901_ (
    .A(\datapath.imm [6]),
    .B(_286__bF$buf1),
    .Y(_308_)
);

NAND2X1 _9902_ (
    .A(\datapath.csr.csr_data [6]),
    .B(_287__bF$buf1),
    .Y(_309_)
);

NAND3X1 _9903_ (
    .A(_308_),
    .B(_309_),
    .C(_307_),
    .Y(\datapath.muxbval [6])
);

NAND2X1 _9904_ (
    .A(\datapath.registers.regb_data [7]),
    .B(_288__bF$buf1),
    .Y(_310_)
);

NAND2X1 _9905_ (
    .A(\datapath.imm [7]),
    .B(_286__bF$buf0),
    .Y(_311_)
);

NAND2X1 _9906_ (
    .A(\datapath.csr.csr_data [7]),
    .B(_287__bF$buf0),
    .Y(_312_)
);

NAND3X1 _9907_ (
    .A(_311_),
    .B(_312_),
    .C(_310_),
    .Y(\datapath.muxbval [7])
);

NAND2X1 _9908_ (
    .A(\datapath.registers.regb_data [8]),
    .B(_288__bF$buf0),
    .Y(_313_)
);

NAND2X1 _9909_ (
    .A(\datapath.imm [8]),
    .B(_286__bF$buf4),
    .Y(_314_)
);

NAND2X1 _9910_ (
    .A(\datapath.csr.csr_data [8]),
    .B(_287__bF$buf4),
    .Y(_315_)
);

NAND3X1 _9911_ (
    .A(_314_),
    .B(_315_),
    .C(_313_),
    .Y(\datapath.muxbval [8])
);

NAND2X1 _9912_ (
    .A(\datapath.registers.regb_data [9]),
    .B(_288__bF$buf4),
    .Y(_316_)
);

NAND2X1 _9913_ (
    .A(\datapath.imm [9]),
    .B(_286__bF$buf3),
    .Y(_317_)
);

NAND2X1 _9914_ (
    .A(\datapath.csr.csr_data [9]),
    .B(_287__bF$buf3),
    .Y(_318_)
);

NAND3X1 _9915_ (
    .A(_317_),
    .B(_318_),
    .C(_316_),
    .Y(\datapath.muxbval [9])
);

NAND2X1 _9916_ (
    .A(\datapath.registers.regb_data [10]),
    .B(_288__bF$buf3),
    .Y(_319_)
);

NAND2X1 _9917_ (
    .A(\datapath.imm [10]),
    .B(_286__bF$buf2),
    .Y(_320_)
);

NAND2X1 _9918_ (
    .A(\datapath.csr.csr_data [10]),
    .B(_287__bF$buf2),
    .Y(_321_)
);

NAND3X1 _9919_ (
    .A(_320_),
    .B(_321_),
    .C(_319_),
    .Y(\datapath.muxbval [10])
);

NAND2X1 _9920_ (
    .A(\datapath.registers.regb_data [11]),
    .B(_288__bF$buf2),
    .Y(_322_)
);

NAND2X1 _9921_ (
    .A(\datapath.immediatedecoder._09_ ),
    .B(_286__bF$buf1),
    .Y(_323_)
);

NAND2X1 _9922_ (
    .A(\datapath.csr.csr_data [11]),
    .B(_287__bF$buf1),
    .Y(_324_)
);

NAND3X1 _9923_ (
    .A(_323_),
    .B(_324_),
    .C(_322_),
    .Y(\datapath.muxbval [11])
);

NAND2X1 _9924_ (
    .A(\datapath.registers.regb_data [12]),
    .B(_288__bF$buf1),
    .Y(_325_)
);

NAND2X1 _9925_ (
    .A(\datapath.imm [12]),
    .B(_286__bF$buf0),
    .Y(_326_)
);

NAND2X1 _9926_ (
    .A(\datapath.csr.csr_data [12]),
    .B(_287__bF$buf0),
    .Y(_327_)
);

NAND3X1 _9927_ (
    .A(_326_),
    .B(_327_),
    .C(_325_),
    .Y(\datapath.muxbval [12])
);

NAND2X1 _9928_ (
    .A(\datapath.registers.regb_data [13]),
    .B(_288__bF$buf0),
    .Y(_328_)
);

NAND2X1 _9929_ (
    .A(\datapath.imm [13]),
    .B(_286__bF$buf4),
    .Y(_329_)
);

NAND2X1 _9930_ (
    .A(\datapath.csr.csr_data [13]),
    .B(_287__bF$buf4),
    .Y(_330_)
);

NAND3X1 _9931_ (
    .A(_329_),
    .B(_330_),
    .C(_328_),
    .Y(\datapath.muxbval [13])
);

NAND2X1 _9932_ (
    .A(\datapath.registers.regb_data [14]),
    .B(_288__bF$buf4),
    .Y(_331_)
);

NAND2X1 _9933_ (
    .A(\datapath.imm [14]),
    .B(_286__bF$buf3),
    .Y(_332_)
);

NAND2X1 _9934_ (
    .A(\datapath.csr.csr_data [14]),
    .B(_287__bF$buf3),
    .Y(_333_)
);

NAND3X1 _9935_ (
    .A(_332_),
    .B(_333_),
    .C(_331_),
    .Y(\datapath.muxbval [14])
);

NAND2X1 _9936_ (
    .A(\datapath.registers.regb_data [15]),
    .B(_288__bF$buf3),
    .Y(_334_)
);

NAND2X1 _9937_ (
    .A(\datapath.imm [15]),
    .B(_286__bF$buf2),
    .Y(_335_)
);

NAND2X1 _9938_ (
    .A(\datapath.csr.csr_data [15]),
    .B(_287__bF$buf2),
    .Y(_336_)
);

NAND3X1 _9939_ (
    .A(_335_),
    .B(_336_),
    .C(_334_),
    .Y(\datapath.muxbval [15])
);

NAND2X1 _9940_ (
    .A(\datapath.registers.regb_data [16]),
    .B(_288__bF$buf2),
    .Y(_337_)
);

NAND2X1 _9941_ (
    .A(\datapath.imm [16]),
    .B(_286__bF$buf1),
    .Y(_338_)
);

NAND2X1 _9942_ (
    .A(\datapath.csr.csr_data [16]),
    .B(_287__bF$buf1),
    .Y(_339_)
);

NAND3X1 _9943_ (
    .A(_338_),
    .B(_339_),
    .C(_337_),
    .Y(\datapath.muxbval [16])
);

NAND2X1 _9944_ (
    .A(\datapath.registers.regb_data [17]),
    .B(_288__bF$buf1),
    .Y(_340_)
);

NAND2X1 _9945_ (
    .A(\datapath.imm [17]),
    .B(_286__bF$buf0),
    .Y(_341_)
);

NAND2X1 _9946_ (
    .A(\datapath.csr.csr_data [17]),
    .B(_287__bF$buf0),
    .Y(_342_)
);

NAND3X1 _9947_ (
    .A(_341_),
    .B(_342_),
    .C(_340_),
    .Y(\datapath.muxbval [17])
);

NAND2X1 _9948_ (
    .A(\datapath.registers.regb_data [18]),
    .B(_288__bF$buf0),
    .Y(_343_)
);

NAND2X1 _9949_ (
    .A(\datapath.imm [18]),
    .B(_286__bF$buf4),
    .Y(_344_)
);

NAND2X1 _9950_ (
    .A(\datapath.csr.csr_data [18]),
    .B(_287__bF$buf4),
    .Y(_345_)
);

NAND3X1 _9951_ (
    .A(_344_),
    .B(_345_),
    .C(_343_),
    .Y(\datapath.muxbval [18])
);

NAND2X1 _9952_ (
    .A(\datapath.registers.regb_data [19]),
    .B(_288__bF$buf4),
    .Y(_346_)
);

NAND2X1 _9953_ (
    .A(\datapath.imm [19]),
    .B(_286__bF$buf3),
    .Y(_347_)
);

NAND2X1 _9954_ (
    .A(\datapath.csr.csr_data [19]),
    .B(_287__bF$buf3),
    .Y(_348_)
);

NAND3X1 _9955_ (
    .A(_347_),
    .B(_348_),
    .C(_346_),
    .Y(\datapath.muxbval [19])
);

NAND2X1 _9956_ (
    .A(\datapath.registers.regb_data [20]),
    .B(_288__bF$buf3),
    .Y(_349_)
);

NAND2X1 _9957_ (
    .A(\datapath.imm [20]),
    .B(_286__bF$buf2),
    .Y(_350_)
);

NAND2X1 _9958_ (
    .A(\datapath.csr.csr_data [20]),
    .B(_287__bF$buf2),
    .Y(_351_)
);

NAND3X1 _9959_ (
    .A(_350_),
    .B(_351_),
    .C(_349_),
    .Y(\datapath.muxbval [20])
);

NAND2X1 _9960_ (
    .A(\datapath.registers.regb_data [21]),
    .B(_288__bF$buf2),
    .Y(_352_)
);

NAND2X1 _9961_ (
    .A(\datapath.imm [21]),
    .B(_286__bF$buf1),
    .Y(_353_)
);

NAND2X1 _9962_ (
    .A(\datapath.csr.csr_data [21]),
    .B(_287__bF$buf1),
    .Y(_354_)
);

NAND3X1 _9963_ (
    .A(_353_),
    .B(_354_),
    .C(_352_),
    .Y(\datapath.muxbval [21])
);

NAND2X1 _9964_ (
    .A(\datapath.registers.regb_data [22]),
    .B(_288__bF$buf1),
    .Y(_355_)
);

NAND2X1 _9965_ (
    .A(\datapath.imm [22]),
    .B(_286__bF$buf0),
    .Y(_356_)
);

NAND2X1 _9966_ (
    .A(\datapath.csr.csr_data [22]),
    .B(_287__bF$buf0),
    .Y(_357_)
);

NAND3X1 _9967_ (
    .A(_356_),
    .B(_357_),
    .C(_355_),
    .Y(\datapath.muxbval [22])
);

NAND2X1 _9968_ (
    .A(\datapath.registers.regb_data [23]),
    .B(_288__bF$buf0),
    .Y(_358_)
);

NAND2X1 _9969_ (
    .A(\datapath.imm [23]),
    .B(_286__bF$buf4),
    .Y(_359_)
);

NAND2X1 _9970_ (
    .A(\datapath.csr.csr_data [23]),
    .B(_287__bF$buf4),
    .Y(_360_)
);

NAND3X1 _9971_ (
    .A(_359_),
    .B(_360_),
    .C(_358_),
    .Y(\datapath.muxbval [23])
);

NAND2X1 _9972_ (
    .A(\datapath.registers.regb_data [24]),
    .B(_288__bF$buf4),
    .Y(_361_)
);

NAND2X1 _9973_ (
    .A(\datapath.imm [24]),
    .B(_286__bF$buf3),
    .Y(_362_)
);

NAND2X1 _9974_ (
    .A(\datapath.csr.csr_data [24]),
    .B(_287__bF$buf3),
    .Y(_363_)
);

NAND3X1 _9975_ (
    .A(_362_),
    .B(_363_),
    .C(_361_),
    .Y(\datapath.muxbval [24])
);

NAND2X1 _9976_ (
    .A(\datapath.registers.regb_data [25]),
    .B(_288__bF$buf3),
    .Y(_364_)
);

NAND2X1 _9977_ (
    .A(\datapath.imm [25]),
    .B(_286__bF$buf2),
    .Y(_365_)
);

NAND2X1 _9978_ (
    .A(\datapath.csr.csr_data [25]),
    .B(_287__bF$buf2),
    .Y(_366_)
);

NAND3X1 _9979_ (
    .A(_365_),
    .B(_366_),
    .C(_364_),
    .Y(\datapath.muxbval [25])
);

NAND2X1 _9980_ (
    .A(\datapath.registers.regb_data [26]),
    .B(_288__bF$buf2),
    .Y(_367_)
);

NAND2X1 _9981_ (
    .A(\datapath.imm [26]),
    .B(_286__bF$buf1),
    .Y(_368_)
);

NAND2X1 _9982_ (
    .A(\datapath.csr.csr_data [26]),
    .B(_287__bF$buf1),
    .Y(_369_)
);

NAND3X1 _9983_ (
    .A(_368_),
    .B(_369_),
    .C(_367_),
    .Y(\datapath.muxbval [26])
);

NAND2X1 _9984_ (
    .A(\datapath.registers.regb_data [27]),
    .B(_288__bF$buf1),
    .Y(_370_)
);

NAND2X1 _9985_ (
    .A(\datapath.imm [27]),
    .B(_286__bF$buf0),
    .Y(_371_)
);

NAND2X1 _9986_ (
    .A(\datapath.csr.csr_data [27]),
    .B(_287__bF$buf0),
    .Y(_372_)
);

NAND3X1 _9987_ (
    .A(_371_),
    .B(_372_),
    .C(_370_),
    .Y(\datapath.muxbval [27])
);

NAND2X1 _9988_ (
    .A(\datapath.registers.regb_data [28]),
    .B(_288__bF$buf0),
    .Y(_373_)
);

NAND2X1 _9989_ (
    .A(\datapath.imm [28]),
    .B(_286__bF$buf4),
    .Y(_374_)
);

NAND2X1 _9990_ (
    .A(\datapath.csr.csr_data [28]),
    .B(_287__bF$buf4),
    .Y(_375_)
);

NAND3X1 _9991_ (
    .A(_374_),
    .B(_375_),
    .C(_373_),
    .Y(\datapath.muxbval [28])
);

NAND2X1 _9992_ (
    .A(\datapath.registers.regb_data [29]),
    .B(_288__bF$buf4),
    .Y(_376_)
);

NAND2X1 _9993_ (
    .A(\datapath.imm [29]),
    .B(_286__bF$buf3),
    .Y(_377_)
);

NAND2X1 _9994_ (
    .A(\datapath.csr.csr_data [29]),
    .B(_287__bF$buf3),
    .Y(_378_)
);

NAND3X1 _9995_ (
    .A(_377_),
    .B(_378_),
    .C(_376_),
    .Y(\datapath.muxbval [29])
);

NAND2X1 _9996_ (
    .A(\datapath.registers.regb_data [30]),
    .B(_288__bF$buf3),
    .Y(_379_)
);

NAND2X1 _9997_ (
    .A(\datapath.imm [30]),
    .B(_286__bF$buf2),
    .Y(_380_)
);

NAND2X1 _9998_ (
    .A(\datapath.csr.csr_data [30]),
    .B(_287__bF$buf2),
    .Y(_381_)
);

NAND3X1 _9999_ (
    .A(_380_),
    .B(_381_),
    .C(_379_),
    .Y(\datapath.muxbval [30])
);

endmodule
