/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */

module RISCV32I(
    inout vdd,
    inout gnd,
    input CLK,
    output [31:0] DMEM_ADDR,
    input [31:0] DMEM_DATA_L,
    output [31:0] DMEM_DATA_S,
    output DMEM_WEN,
    output [31:0] IMEM_ADDR,
    input [31:0] IMEM_DATA,
    input IRQ
);

wire _9417_ ;
wire _4972_ ;
wire _4552_ ;
wire _4132_ ;
wire _5757_ ;
wire _5337_ ;
wire _9170_ ;
wire _5488__bF$buf0 ;
wire _5488__bF$buf1 ;
wire _5488__bF$buf2 ;
wire _5488__bF$buf3 ;
wire _5488__bF$buf4 ;
wire _1677_ ;
wire _1257_ ;
wire _7903_ ;
wire _5090_ ;
wire _588_ ;
wire _168_ ;
wire _3823_ ;
wire _3403_ ;
wire _6295_ ;
wire _4608_ ;
wire _8861_ ;
wire _8441_ ;
wire _8021_ ;
wire \datapath.alu.b_4_bF$buf1  ;
wire _9226_ ;
wire _4781_ ;
wire _4361_ ;
wire _800_ ;
wire _5986_ ;
wire _5566_ ;
wire _5146_ ;
wire _60_ ;
wire _1486_ ;
wire _1066_ ;
wire _7712_ ;
wire _397_ ;
wire _8917_ ;
wire _3632_ ;
wire _3212_ ;
wire _4837_ ;
wire _4417_ ;
wire _8670_ ;
wire _8250_ ;
wire \datapath.immediatedecoder._06_  ;
wire _9035_ ;
wire _4590_ ;
wire _4170_ ;
wire _2903_ ;
wire _5795_ ;
wire _5375_ ;
wire _2708__bF$buf0 ;
wire _2708__bF$buf1 ;
wire _2708__bF$buf2 ;
wire _2708__bF$buf3 ;
wire _1295_ ;
wire _7941_ ;
wire _7521_ ;
wire _7101_ ;
wire _8726_ ;
wire _8306_ ;
wire _3861_ ;
wire _3441_ ;
wire _3021_ ;
wire _4646_ ;
wire _4226_ ;
wire CLK_bF$buf50 ;
wire CLK_bF$buf51 ;
wire CLK_bF$buf52 ;
wire CLK_bF$buf53 ;
wire CLK_bF$buf54 ;
wire CLK_bF$buf55 ;
wire CLK_bF$buf56 ;
wire CLK_bF$buf57 ;
wire CLK_bF$buf58 ;
wire CLK_bF$buf59 ;
wire _9264_ ;
wire _2712_ ;
wire _5184_ ;
wire _3917_ ;
wire _6389_ ;
wire _7750_ ;
wire _7330_ ;
wire _4193__bF$buf0 ;
wire _4193__bF$buf1 ;
wire _4193__bF$buf2 ;
wire _4193__bF$buf3 ;
wire _4193__bF$buf4 ;
wire _8955_ ;
wire _8535_ ;
wire _8115_ ;
wire _3670_ ;
wire _3250_ ;
wire _4875_ ;
wire _4455_ ;
wire _4035_ ;
wire [31:0] \datapath.memoryinterface.byte_size_store.storebyte  ;
wire _6601_ ;
wire _9073_ ;
wire _7806_ ;
wire _2941_ ;
wire _2521_ ;
wire _2101_ ;
wire [31:0] \datapath.registers.1226[22]  ;
wire _3726_ ;
wire _3306_ ;
wire _6198_ ;
wire _8764_ ;
wire _8344_ ;
wire _9129_ ;
wire _4684_ ;
wire _4264_ ;
wire _703_ ;
wire _5889_ ;
wire _5469_ ;
wire _5049_ ;
wire _6830_ ;
wire _6410_ ;
wire _1389_ ;
wire _7615_ ;
wire _2750_ ;
wire _2330_ ;
wire _3955_ ;
wire _3535_ ;
wire _3115_ ;
wire _8993_ ;
wire _8573_ ;
wire _8153_ ;
wire _19_ ;
wire _1601_ ;
wire _9358_ ;
wire _4493_ ;
wire _4073_ ;
wire \datapath.idinstr_20_bF$buf12  ;
wire _932_ ;
wire _512_ ;
wire _2806_ ;
wire _5698_ ;
wire _5278_ ;
wire [1:0] asel ;
wire _1198_ ;
wire _7844_ ;
wire _7424_ ;
wire _7004_ ;
wire _8629_ ;
wire _8209_ ;
wire _3764_ ;
wire _3344_ ;
wire _4969_ ;
wire _4549_ ;
wire \datapath.idinstr_21_bF$buf21  ;
wire _4129_ ;
wire _5910_ ;
wire _8382_ ;
wire _1830_ ;
wire _1410_ ;
wire _9167_ ;
wire _741_ ;
wire _321_ ;
wire _2615_ ;
wire _5087_ ;
wire \datapath.idinstr_15_bF$buf26  ;
wire \datapath.idinstr_22_bF$buf30  ;
wire _7653_ ;
wire _7233_ ;
wire _8858_ ;
wire _8438_ ;
wire _8018_ ;
wire _3993_ ;
wire _3573_ ;
wire _3153_ ;
wire \bypassandflushunit.stall_bF$buf0  ;
wire _4778_ ;
wire _4358_ ;
wire _8191_ ;
wire \datapath.idinstr_16_bF$buf35  ;
wire _57_ ;
wire _6924_ ;
wire _6504_ ;
wire _9396_ ;
wire \datapath.idinstr_20_bF$buf50  ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _7709_ ;
wire _2844_ ;
wire _2424_ ;
wire _2004_ ;
wire _3629_ ;
wire _3209_ ;
wire _7882_ ;
wire _7462_ ;
wire _7042_ ;
wire _8667_ ;
wire _8247_ ;
wire _3382_ ;
wire _4587_ ;
wire _4167_ ;
wire _606_ ;
wire _6733_ ;
wire _6313_ ;
wire _7938_ ;
wire _7518_ ;
wire _2653_ ;
wire _2233_ ;
wire _3858_ ;
wire _3438_ ;
wire _3018_ ;
wire _7691_ ;
wire _7271_ ;
wire _8896_ ;
wire _8476_ ;
wire _8056_ ;
wire _3191_ ;
wire _5436__bF$buf0 ;
wire _5436__bF$buf1 ;
wire _5436__bF$buf2 ;
wire _5436__bF$buf3 ;
wire _1924_ ;
wire _5436__bF$buf4 ;
wire _1504_ ;
wire _4396_ ;
wire _835_ ;
wire _415_ ;
wire _2709_ ;
wire _95_ ;
wire _6962_ ;
wire _6542_ ;
wire _6122_ ;
wire _7747_ ;
wire _7327_ ;
wire _2882_ ;
wire _2462_ ;
wire _2042_ ;
wire _3667_ ;
wire _3247_ ;
wire _7080_ ;
wire _5813_ ;
wire _8285_ ;
wire _5440__bF$buf0 ;
wire _5440__bF$buf1 ;
wire _5440__bF$buf2 ;
wire _5440__bF$buf3 ;
wire _5440__bF$buf4 ;
wire _1733_ ;
wire _1313_ ;
wire _1236__bF$buf0 ;
wire _1236__bF$buf1 ;
wire _1236__bF$buf2 ;
wire _1236__bF$buf3 ;
wire _644_ ;
wire _1236__bF$buf4 ;
wire _224_ ;
wire _2938_ ;
wire _2518_ ;
wire _6771_ ;
wire _6351_ ;
wire _7976_ ;
wire _7556_ ;
wire _7136_ ;
wire _2691_ ;
wire _2271_ ;
wire _3896_ ;
wire _3476_ ;
wire _3056_ ;
wire _5622_ ;
wire _5202_ ;
wire _8094_ ;
wire _6827_ ;
wire _6407_ ;
wire _1962_ ;
wire _1542_ ;
wire _1122_ ;
wire _9299_ ;
wire _1240__bF$buf0 ;
wire _1240__bF$buf1 ;
wire _1240__bF$buf2 ;
wire _1240__bF$buf3 ;
wire _1240__bF$buf4 ;
wire _873_ ;
wire _453_ ;
wire _2747_ ;
wire _2327_ ;
wire _6580_ ;
wire _6160_ ;
wire _7785_ ;
wire _7365_ ;
wire _2080_ ;
wire _3285_ ;
wire _5851_ ;
wire _5431_ ;
wire _5011_ ;
wire _929_ ;
wire _509_ ;
wire _6636_ ;
wire _6216_ ;
wire _1771_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _2976_ ;
wire _2556_ ;
wire _2136_ ;
wire _4702_ ;
wire _7594_ ;
wire _7174_ ;
wire \datapath.idinstr_21_bF$buf18  ;
wire _5907_ ;
wire _8799_ ;
wire _8379_ ;
wire _3094_ ;
wire _9320_ ;
wire _1827_ ;
wire _1407_ ;
wire _4299_ ;
wire _5660_ ;
wire _5240_ ;
wire _738_ ;
wire _318_ ;
wire \datapath.idinstr_17_bF$buf3  ;
wire _6865_ ;
wire _6445_ ;
wire _6025_ ;
wire _1580_ ;
wire _1160_ ;
wire _491_ ;
wire \datapath.idinstr_22_bF$buf27  ;
wire _2785_ ;
wire _2365_ ;
wire _9210__bF$buf0 ;
wire _9210__bF$buf1 ;
wire _9210__bF$buf2 ;
wire _9210__bF$buf3 ;
wire _9210__bF$buf4 ;
wire _4931_ ;
wire _4511_ ;
wire _5716_ ;
wire _2865__bF$buf0 ;
wire _2865__bF$buf1 ;
wire _2865__bF$buf2 ;
wire _2865__bF$buf3 ;
wire _8188_ ;
wire _1636_ ;
wire _1216_ ;
wire \datapath.idinstr_21_bF$buf3  ;
wire \datapath.idinstr_20_bF$buf47  ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _6674_ ;
wire _6254_ ;
wire _7879_ ;
wire _7459_ ;
wire _7039_ ;
wire _2594_ ;
wire _2174_ ;
wire _8820_ ;
wire _8400_ ;
wire _3799_ ;
wire _3379_ ;
wire _4740_ ;
wire _4320_ ;
wire _5945_ ;
wire _5525_ ;
wire _5105_ ;
wire _1865_ ;
wire _1445_ ;
wire _1025_ ;
wire _776_ ;
wire _356_ ;
wire _6483_ ;
wire _6063_ ;
wire _7688_ ;
wire _7268_ ;
wire _3188_ ;
wire _9414_ ;
wire _5754_ ;
wire _5334_ ;
wire _6959_ ;
wire _6539_ ;
wire _6119_ ;
wire _1674_ ;
wire _1254_ ;
wire _7900_ ;
wire _585_ ;
wire _165_ ;
wire _2879_ ;
wire _2459_ ;
wire _2039_ ;
wire _3820_ ;
wire _3400_ ;
wire _6292_ ;
wire _4605_ ;
wire _7497_ ;
wire _7077_ ;
wire _9223_ ;
wire _5983_ ;
wire _5563_ ;
wire _5143_ ;
wire _6768_ ;
wire _6348_ ;
wire _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _2688_ ;
wire _2268_ ;
wire _8914_ ;
wire _4834_ ;
wire _4414_ ;
wire _5619_ ;
wire _9032_ ;
wire \datapath.alu.b_2_bF$buf5  ;
wire _1959_ ;
wire _1539_ ;
wire _1119_ ;
wire _2900_ ;
wire _5792_ ;
wire _5372_ ;
wire _6997_ ;
wire _6577_ ;
wire _6157_ ;
wire _1292_ ;
wire _2497_ ;
wire _2077_ ;
wire _8723_ ;
wire _8303_ ;
wire _4643_ ;
wire _4223_ ;
wire CLK_bF$buf20 ;
wire CLK_bF$buf21 ;
wire CLK_bF$buf22 ;
wire CLK_bF$buf23 ;
wire CLK_bF$buf24 ;
wire CLK_bF$buf25 ;
wire CLK_bF$buf26 ;
wire CLK_bF$buf27 ;
wire CLK_bF$buf28 ;
wire CLK_bF$buf29 ;
wire _5848_ ;
wire _5428_ ;
wire _5008_ ;
wire _9261_ ;
wire _1768_ ;
wire _1348_ ;
wire _5181_ ;
wire _679_ ;
wire _259_ ;
wire _3914_ ;
wire _6386_ ;
wire _8952_ ;
wire _8532_ ;
wire _8112_ ;
wire _9317_ ;
wire _4872_ ;
wire _4452_ ;
wire _4032_ ;
wire _5657_ ;
wire _5237_ ;
wire _9070_ ;
wire _1997_ ;
wire _1577_ ;
wire _1157_ ;
wire _7803_ ;
wire _488_ ;
wire _3723_ ;
wire _3303_ ;
wire _6195_ ;
wire _4928_ ;
wire _4508_ ;
wire _8761_ ;
wire _8341_ ;
wire _9126_ ;
wire _4681_ ;
wire _4261_ ;
wire _700_ ;
wire _5886_ ;
wire _5466_ ;
wire _5046_ ;
wire _6107__bF$buf0 ;
wire _6107__bF$buf1 ;
wire _6107__bF$buf2 ;
wire _6107__bF$buf3 ;
wire _6107__bF$buf4 ;
wire _1386_ ;
wire _7612_ ;
wire _297_ ;
wire \datapath.idinstr_20_hier0_bF$buf4  ;
wire _8817_ ;
wire _3952_ ;
wire _3532_ ;
wire _3112_ ;
wire _4737_ ;
wire _4317_ ;
wire _8990_ ;
wire _8570_ ;
wire _8150_ ;
wire _16_ ;
wire _9355_ ;
wire _4490_ ;
wire _4070_ ;
wire _2803_ ;
wire _5695_ ;
wire _5275_ ;
wire _1195_ ;
wire _7841_ ;
wire _7421_ ;
wire _7001_ ;
wire [31:0] \datapath.regcwb  ;
wire _8626_ ;
wire _8206_ ;
wire _3761_ ;
wire _3341_ ;
wire _4966_ ;
wire _4546_ ;
wire _4126_ ;
wire _4196__bF$buf0 ;
wire _4196__bF$buf1 ;
wire _4196__bF$buf2 ;
wire _4196__bF$buf3 ;
wire _4196__bF$buf4 ;
wire _9164_ ;
wire _2612_ ;
wire _5084_ ;
wire \datapath.idinstr_15_bF$buf23  ;
wire _3817_ ;
wire _6289_ ;
wire _7650_ ;
wire _7230_ ;
wire _8855_ ;
wire _8435_ ;
wire _8015_ ;
wire _3990_ ;
wire _3570_ ;
wire _3150_ ;
wire _4775_ ;
wire _4355_ ;
wire [31:0] \datapath.csr.mvect  ;
wire \datapath.idinstr_16_bF$buf32  ;
wire _54_ ;
wire _6921_ ;
wire _6501_ ;
wire _9393_ ;
wire _7706_ ;
wire _2841_ ;
wire _2421_ ;
wire _2001_ ;
wire [31:0] \datapath.registers.1226[12]  ;
wire _3626_ ;
wire _3206_ ;
wire _6098_ ;
wire _8664_ ;
wire _8244_ ;
wire \datapath.idinstr_17_bF$buf41  ;
wire _9029_ ;
wire _4584_ ;
wire _4164_ ;
wire _603_ ;
wire _5789_ ;
wire _5369_ ;
wire _6730_ ;
wire _6310_ ;
wire _1289_ ;
wire _7935_ ;
wire _7515_ ;
wire _2650_ ;
wire _2230_ ;
wire _3855_ ;
wire _3435_ ;
wire _3015_ ;
wire _8893_ ;
wire _8473_ ;
wire _8053_ ;
wire _1921_ ;
wire _1501_ ;
wire _9258_ ;
wire _4393_ ;
wire _832_ ;
wire _412_ ;
wire _2706_ ;
wire _5598_ ;
wire _5178_ ;
wire _92_ ;
wire _1098_ ;
wire _7744_ ;
wire _7324_ ;
wire _8949_ ;
wire _8529_ ;
wire _8109_ ;
wire _3664_ ;
wire _3244_ ;
wire _4869_ ;
wire _4449_ ;
wire _4029_ ;
wire _5810_ ;
wire _8282_ ;
wire _1730_ ;
wire _1310_ ;
wire _9067_ ;
wire _641_ ;
wire _221_ ;
wire _2935_ ;
wire _2515_ ;
wire _7973_ ;
wire _7553_ ;
wire _7133_ ;
wire _8758_ ;
wire _8338_ ;
wire _3893_ ;
wire _3473_ ;
wire _3053_ ;
wire _4678_ ;
wire _4258_ ;
wire _8091_ ;
wire _6824_ ;
wire _6404_ ;
wire _9296_ ;
wire _870_ ;
wire _450_ ;
wire _7609_ ;
wire _2744_ ;
wire _2324_ ;
wire _3949_ ;
wire _3529_ ;
wire _3109_ ;
wire _7782_ ;
wire _7362_ ;
wire _8987_ ;
wire _8567_ ;
wire _8147_ ;
wire _3282_ ;
wire _4487_ ;
wire _4067_ ;
wire _926_ ;
wire _506_ ;
wire _6633_ ;
wire _6213_ ;
wire _7838_ ;
wire _7418_ ;
wire _2973_ ;
wire _2553_ ;
wire _2133_ ;
wire _3758_ ;
wire _3338_ ;
wire _7591_ ;
wire _7171_ ;
wire \datapath.idinstr_21_bF$buf15  ;
wire _5904_ ;
wire _8796_ ;
wire _8376_ ;
wire _3091_ ;
wire \datapath.regmret_bF$buf4  ;
wire _1824_ ;
wire _1404_ ;
wire _4296_ ;
wire _735_ ;
wire _315_ ;
wire \datapath.idinstr_17_bF$buf0  ;
wire _2609_ ;
wire _6862_ ;
wire _6442_ ;
wire _6022_ ;
wire \datapath.idinstr_22_bF$buf24  ;
wire _7647_ ;
wire _7227_ ;
wire _2782_ ;
wire _2362_ ;
wire _3987_ ;
wire _3567_ ;
wire _3147_ ;
wire _5713_ ;
wire _8185_ ;
wire \datapath.idinstr_16_bF$buf29  ;
wire _6918_ ;
wire _1633_ ;
wire _1213_ ;
wire \datapath.idinstr_21_bF$buf0  ;
wire \datapath.idinstr_20_bF$buf44  ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire _2838_ ;
wire \datapath.idinstr_15_bF$buf7  ;
wire _2418_ ;
wire _6671_ ;
wire _963__bF$buf0 ;
wire _6251_ ;
wire _963__bF$buf1 ;
wire \controlunit.mret  ;
wire _963__bF$buf2 ;
wire _963__bF$buf3 ;
wire _963__bF$buf4 ;
wire _7876_ ;
wire _7456_ ;
wire _7036_ ;
wire _2591_ ;
wire _2171_ ;
wire IRQ ;
wire [31:0] \datapath.registers.1226[29]  ;
wire _3796_ ;
wire _3376_ ;
wire \datapath.idinstr_17_bF$buf38  ;
wire _5942_ ;
wire _5522_ ;
wire _5102_ ;
wire _6727_ ;
wire _6307_ ;
wire _1862_ ;
wire _1442_ ;
wire _1022_ ;
wire _9199_ ;
wire _773_ ;
wire _353_ ;
wire _2647_ ;
wire _2227_ ;
wire _6480_ ;
wire _6060_ ;
wire _7685_ ;
wire _7265_ ;
wire _3185_ ;
wire _9411_ ;
wire _1918_ ;
wire _5751_ ;
wire _5331_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _6956_ ;
wire _6536_ ;
wire _6116_ ;
wire _1671_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _2876_ ;
wire _2456_ ;
wire _2036_ ;
wire _4602_ ;
wire _7494_ ;
wire _7074_ ;
wire _5807_ ;
wire _8699_ ;
wire _8279_ ;
wire _9220_ ;
wire _1727_ ;
wire _1307_ ;
wire _4199_ ;
wire _5980_ ;
wire _5560_ ;
wire _5140_ ;
wire _638_ ;
wire _218_ ;
wire _6765_ ;
wire _6345_ ;
wire _1480_ ;
wire _1060_ ;
wire _391_ ;
wire \datapath.idinstr_24_bF$buf3  ;
wire _2685_ ;
wire _2265_ ;
wire _8911_ ;
wire _4831_ ;
wire _4411_ ;
wire _5616_ ;
wire _8088_ ;
wire \datapath.alu.b_2_bF$buf2  ;
wire _1956_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire _6994_ ;
wire _6574_ ;
wire _6154_ ;
wire [2:0] \datapath._31_  ;
wire _7779_ ;
wire _7359_ ;
wire _2494_ ;
wire _2074_ ;
wire _8720_ ;
wire _8300_ ;
wire _3699_ ;
wire _3279_ ;
wire _4640_ ;
wire _4220_ ;
wire _2703__bF$buf0 ;
wire _2703__bF$buf1 ;
wire _2703__bF$buf2 ;
wire _5845_ ;
wire _2703__bF$buf3 ;
wire _5425_ ;
wire _5005_ ;
wire _1765_ ;
wire _1345_ ;
wire _676_ ;
wire _256_ ;
wire _3911_ ;
wire _6383_ ;
wire _7588_ ;
wire _7168_ ;
wire _3088_ ;
wire _9314_ ;
wire _5510__bF$buf0 ;
wire _5510__bF$buf1 ;
wire _5510__bF$buf2 ;
wire _5510__bF$buf3 ;
wire _5510__bF$buf4 ;
wire _5510__bF$buf5 ;
wire _5510__bF$buf6 ;
wire _5510__bF$buf7 ;
wire _5510__bF$buf8 ;
wire _5510__bF$buf9 ;
wire _5654_ ;
wire _5234_ ;
wire _6859_ ;
wire _6439_ ;
wire _6019_ ;
wire _1994_ ;
wire _1574_ ;
wire _1154_ ;
wire _7800_ ;
wire _485_ ;
wire _2779_ ;
wire _2359_ ;
wire _3720_ ;
wire _3300_ ;
wire _6192_ ;
wire _4925_ ;
wire _4505_ ;
wire _7397_ ;
wire _9123_ ;
wire _5883_ ;
wire _5463_ ;
wire _5043_ ;
wire _6668_ ;
wire _6248_ ;
wire _1383_ ;
wire _294_ ;
wire _2588_ ;
wire _2168_ ;
wire \datapath.idinstr_20_hier0_bF$buf1  ;
wire _8814_ ;
wire _4734_ ;
wire _4314_ ;
wire _5939_ ;
wire _5519_ ;
wire _13_ ;
wire _9352_ ;
wire _1859_ ;
wire _1439_ ;
wire _1019_ ;
wire _2800_ ;
wire _5692_ ;
wire _5272_ ;
wire _6897_ ;
wire _6477_ ;
wire _6057_ ;
wire _1192_ ;
wire _2397_ ;
wire _8623_ ;
wire _8203_ ;
wire _9408_ ;
wire _4963_ ;
wire _4543_ ;
wire _4123_ ;
wire _5748_ ;
wire _5328_ ;
wire \datapath.alu.condtrue  ;
wire _9161_ ;
wire _1668_ ;
wire _1248_ ;
wire _5081_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire \datapath.idinstr_15_bF$buf20  ;
wire _3814_ ;
wire _6286_ ;
wire _8852_ ;
wire _8432_ ;
wire _8012_ ;
wire _5498__bF$buf0 ;
wire _5498__bF$buf1 ;
wire _5498__bF$buf2 ;
wire _5498__bF$buf3 ;
wire _5498__bF$buf4 ;
wire _9217_ ;
wire _4772_ ;
wire _4352_ ;
wire _5977_ ;
wire _5557_ ;
wire _5137_ ;
wire _51_ ;
wire _9390_ ;
wire _1897_ ;
wire _1477_ ;
wire _1057_ ;
wire _7703_ ;
wire _388_ ;
wire _8908_ ;
wire _3623_ ;
wire _3203_ ;
wire _6095_ ;
wire _4828_ ;
wire _4408_ ;
wire _8661_ ;
wire _8241_ ;
wire _9026_ ;
wire _4581_ ;
wire _4161_ ;
wire _600_ ;
wire _5786_ ;
wire _5366_ ;
wire _1286_ ;
wire _7932_ ;
wire _7512_ ;
wire _197_ ;
wire _8717_ ;
wire _3852_ ;
wire _3432_ ;
wire _3012_ ;
wire _4637_ ;
wire _4217_ ;
wire [31:0] \datapath._06_  ;
wire _8890_ ;
wire _8470_ ;
wire _8050_ ;
wire _9255_ ;
wire _4390_ ;
wire _2703_ ;
wire _5595_ ;
wire _5175_ ;
wire _3908_ ;
wire _1095_ ;
wire _7741_ ;
wire _7321_ ;
wire _8946_ ;
wire _8526_ ;
wire _8106_ ;
wire _3661_ ;
wire _3241_ ;
wire _4866_ ;
wire _4446_ ;
wire _4026_ ;
wire _9064_ ;
wire _2932_ ;
wire _2512_ ;
wire _3717_ ;
wire _6189_ ;
wire _7970_ ;
wire _7550_ ;
wire _7130_ ;
wire _8755_ ;
wire _8335_ ;
wire _3890_ ;
wire _3470_ ;
wire _3050_ ;
wire _4675_ ;
wire _4255_ ;
wire _6821_ ;
wire _6401_ ;
wire _9293_ ;
wire _7606_ ;
wire _2741_ ;
wire _2321_ ;
wire _3946_ ;
wire _3526_ ;
wire _3106_ ;
wire _7_ ;
wire _8984_ ;
wire _8564_ ;
wire _8144_ ;
wire _9349_ ;
wire _4484_ ;
wire _4064_ ;
wire _923_ ;
wire _503_ ;
wire _5689_ ;
wire _5269_ ;
wire _6630_ ;
wire _6210_ ;
wire _1189_ ;
wire _7835_ ;
wire _7415_ ;
wire _2970_ ;
wire _2550_ ;
wire _2130_ ;
wire _3755_ ;
wire _3335_ ;
wire \datapath.idinstr_21_bF$buf12  ;
wire _5901_ ;
wire _8793_ ;
wire _8373_ ;
wire \datapath.regmret_bF$buf1  ;
wire _1821_ ;
wire _1401_ ;
wire _9158_ ;
wire _4293_ ;
wire _732_ ;
wire _312_ ;
wire _2606_ ;
wire _5498_ ;
wire _5078_ ;
wire \datapath.idinstr_15_bF$buf17  ;
wire \datapath.idinstr_15_hier0_bF$buf5  ;
wire \datapath.idinstr_22_bF$buf21  ;
wire _7644_ ;
wire _7224_ ;
wire [31:0] \datapath.registers.1226[3]  ;
wire _8849_ ;
wire _8429_ ;
wire _8009_ ;
wire _3984_ ;
wire _3564_ ;
wire _3144_ ;
wire _4769_ ;
wire _4349_ ;
wire _5710_ ;
wire _8182_ ;
wire \datapath.idinstr_16_bF$buf26  ;
wire _48_ ;
wire _6915_ ;
wire _1630_ ;
wire _1210_ ;
wire _9387_ ;
wire \datapath.idinstr_20_bF$buf41  ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _2835_ ;
wire \datapath.idinstr_15_bF$buf4  ;
wire _2415_ ;
wire _7873_ ;
wire _7453_ ;
wire _7033_ ;
wire _8658_ ;
wire _8238_ ;
wire _3793_ ;
wire _3373_ ;
wire \datapath.idinstr_17_bF$buf35  ;
wire _4998_ ;
wire _4578_ ;
wire _4158_ ;
wire _6724_ ;
wire _6304_ ;
wire _9196_ ;
wire _770_ ;
wire _350_ ;
wire _7929_ ;
wire _7509_ ;
wire _2644_ ;
wire _2224_ ;
wire _3849_ ;
wire _3429_ ;
wire _3009_ ;
wire _7682_ ;
wire _7262_ ;
wire _8887_ ;
wire _8467_ ;
wire _8047_ ;
wire _3182_ ;
wire _1915_ ;
wire _4387_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _6953_ ;
wire _6533_ ;
wire _6113_ ;
wire _7738_ ;
wire _7318_ ;
wire _2873_ ;
wire _2453_ ;
wire _2033_ ;
wire _3658_ ;
wire _3238_ ;
wire _2497__bF$buf0 ;
wire _2497__bF$buf1 ;
wire _2497__bF$buf2 ;
wire _5446__bF$buf0 ;
wire _2497__bF$buf3 ;
wire _5446__bF$buf1 ;
wire _2497__bF$buf4 ;
wire _5446__bF$buf2 ;
wire _2497__bF$buf5 ;
wire _5446__bF$buf3 ;
wire _2497__bF$buf6 ;
wire _5446__bF$buf4 ;
wire _7491_ ;
wire _7071_ ;
wire _5804_ ;
wire _8696_ ;
wire _8276_ ;
wire [31:0] \datapath.csr._32_  ;
wire _1724_ ;
wire _1304_ ;
wire _4196_ ;
wire _635_ ;
wire _215_ ;
wire _2929_ ;
wire _2509_ ;
wire _6762_ ;
wire _6342_ ;
wire _7967_ ;
wire _7547_ ;
wire _7127_ ;
wire \datapath.idinstr_24_bF$buf0  ;
wire _2682_ ;
wire _2262_ ;
wire \datapath.idinstr_18_bF$buf7  ;
wire _5450__bF$buf0 ;
wire _5450__bF$buf1 ;
wire _5450__bF$buf2 ;
wire _5450__bF$buf3 ;
wire _5450__bF$buf4 ;
wire _3887_ ;
wire _3467_ ;
wire _3047_ ;
wire _5613_ ;
wire _8085_ ;
wire \datapath.pcstall_bF$buf6  ;
wire _6818_ ;
wire _1953_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire _2738_ ;
wire _2318_ ;
wire _6991_ ;
wire _6571_ ;
wire _6151_ ;
wire _7776_ ;
wire _7356_ ;
wire _2491_ ;
wire _2071_ ;
wire \datapath.idinstr_22_bF$buf7  ;
wire _970__bF$buf0 ;
wire _970__bF$buf1 ;
wire _970__bF$buf2 ;
wire [31:0] \datapath.registers.1226[19]  ;
wire _970__bF$buf3 ;
wire _970__bF$buf4 ;
wire _3696_ ;
wire _3276_ ;
wire _5842_ ;
wire _5422_ ;
wire _5002_ ;
wire _6627_ ;
wire _6207_ ;
wire _1762_ ;
wire _1342_ ;
wire _9099_ ;
wire _673_ ;
wire _253_ ;
wire _2967_ ;
wire _2547_ ;
wire _2127_ ;
wire _6380_ ;
wire _7585_ ;
wire _7165_ ;
wire _3085_ ;
wire _9311_ ;
wire _1818_ ;
wire _5651_ ;
wire _5231_ ;
wire _729_ ;
wire _309_ ;
wire _6856_ ;
wire _6436_ ;
wire _6016_ ;
wire _1991_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire \datapath.idinstr_22_bF$buf18  ;
wire _2776_ ;
wire _2356_ ;
wire _4922_ ;
wire _4502_ ;
wire _7394_ ;
wire _5707_ ;
wire _8599_ ;
wire _8179_ ;
wire _9120_ ;
wire _1627_ ;
wire _1207_ ;
wire _4099_ ;
wire _5880_ ;
wire _5460_ ;
wire _5040_ ;
wire \datapath.idinstr_20_bF$buf38  ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _6665_ ;
wire _6245_ ;
wire _1380_ ;
wire _291_ ;
wire _2585_ ;
wire _2165_ ;
wire _8811_ ;
wire _4731_ ;
wire _4311_ ;
wire _5936_ ;
wire _5516_ ;
wire _10_ ;
wire \datapath.alu.b_0_bF$buf8  ;
wire _1856_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire _2706__bF$buf0 ;
wire _2706__bF$buf1 ;
wire _2706__bF$buf2 ;
wire _2706__bF$buf3 ;
wire _5509__bF$buf0 ;
wire _5509__bF$buf1 ;
wire _5509__bF$buf2 ;
wire _5509__bF$buf3 ;
wire _5509__bF$buf4 ;
wire _6894_ ;
wire _6474_ ;
wire _6054_ ;
wire _7679_ ;
wire _7259_ ;
wire _2394_ ;
wire _8620_ ;
wire _8200_ ;
wire _3599_ ;
wire _3179_ ;
wire _9405_ ;
wire _4960_ ;
wire _4540_ ;
wire _4120_ ;
wire _5745_ ;
wire _5325_ ;
wire _1665_ ;
wire _1245_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _3811_ ;
wire _6283_ ;
wire \datapath.csr.mie  ;
wire _7488_ ;
wire _7068_ ;
wire _9214_ ;
wire \datapath.idinstr_21_hier0_bF$buf3  ;
wire _5974_ ;
wire _5554_ ;
wire _5134_ ;
wire _6759_ ;
wire _6339_ ;
wire _1894_ ;
wire _1474_ ;
wire _1054_ ;
wire _7700_ ;
wire _385_ ;
wire _2679_ ;
wire _2259_ ;
wire _8905_ ;
wire _3620_ ;
wire _3200_ ;
wire _6092_ ;
wire _4825_ ;
wire _4405_ ;
wire _7297_ ;
wire _9023_ ;
wire _5783_ ;
wire _5363_ ;
wire _6988_ ;
wire _6568_ ;
wire _6148_ ;
wire _1283_ ;
wire _194_ ;
wire _2488_ ;
wire _2068_ ;
wire _8714_ ;
wire _4634_ ;
wire _4214_ ;
wire _5839_ ;
wire _5419_ ;
wire _9252_ ;
wire _1759_ ;
wire _1339_ ;
wire _2700_ ;
wire _5592_ ;
wire _5172_ ;
wire _3905_ ;
wire _6797_ ;
wire _6377_ ;
wire _1092_ ;
wire _2297_ ;
wire _8943_ ;
wire _8523_ ;
wire _8103_ ;
wire _9308_ ;
wire _4863_ ;
wire _4443_ ;
wire _4023_ ;
wire _5648_ ;
wire _5228_ ;
wire _9061_ ;
wire _1988_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire _3714_ ;
wire _6186_ ;
wire _4919_ ;
wire _8752_ ;
wire _8332_ ;
wire _9117_ ;
wire _4672_ ;
wire _4252_ ;
wire _5877_ ;
wire _5457_ ;
wire _5037_ ;
wire _9290_ ;
wire _1797_ ;
wire _1377_ ;
wire _7603_ ;
wire _288_ ;
wire _8808_ ;
wire _3943_ ;
wire _3523_ ;
wire _3103_ ;
wire _4_ ;
wire _4728_ ;
wire _4308_ ;
wire _8981_ ;
wire _8561_ ;
wire _8141_ ;
wire _9346_ ;
wire _4481_ ;
wire _4061_ ;
wire _920_ ;
wire _500_ ;
wire _5686_ ;
wire _5266_ ;
wire _1186_ ;
wire _7832_ ;
wire _7412_ ;
wire _8617_ ;
wire _3752_ ;
wire _3332_ ;
wire _4957_ ;
wire _4537_ ;
wire _4117_ ;
wire _8790_ ;
wire _8370_ ;
wire _9155_ ;
wire _4290_ ;
wire _2603_ ;
wire _5495_ ;
wire _5075_ ;
wire CLK_bF$buf140 ;
wire CLK_bF$buf141 ;
wire CLK_bF$buf142 ;
wire CLK_bF$buf143 ;
wire CLK_bF$buf144 ;
wire CLK_bF$buf145 ;
wire \datapath.idinstr_15_bF$buf14  ;
wire CLK_bF$buf146 ;
wire CLK_bF$buf147 ;
wire CLK_bF$buf148 ;
wire \datapath.csr.meta_irq  ;
wire _3808_ ;
wire CLK_bF$buf149 ;
wire \datapath.idinstr_15_hier0_bF$buf2  ;
wire _7641_ ;
wire _7221_ ;
wire _8846_ ;
wire _8426_ ;
wire _8006_ ;
wire _3981_ ;
wire _3561_ ;
wire _3141_ ;
wire _4766_ ;
wire _4346_ ;
wire \datapath.idinstr_16_bF$buf23  ;
wire _45_ ;
wire _6912_ ;
wire _9384_ ;
wire _2832_ ;
wire \datapath.idinstr_15_bF$buf1  ;
wire _2412_ ;
wire _3617_ ;
wire _6089_ ;
wire _7870_ ;
wire _7450_ ;
wire _7030_ ;
wire _8655_ ;
wire _8235_ ;
wire _3790_ ;
wire _3370_ ;
wire \datapath.idinstr_17_bF$buf32  ;
wire _4995_ ;
wire _4575_ ;
wire _4155_ ;
wire _6721_ ;
wire _6301_ ;
wire _9193_ ;
wire _7926_ ;
wire _7506_ ;
wire _2641_ ;
wire _2221_ ;
wire \datapath.idinstr_15_bF$buf52  ;
wire _3846_ ;
wire _3426_ ;
wire _3006_ ;
wire _3448__bF$buf0 ;
wire _3448__bF$buf1 ;
wire _3448__bF$buf2 ;
wire _3448__bF$buf3 ;
wire _3448__bF$buf4 ;
wire _8884_ ;
wire _8464_ ;
wire _8044_ ;
wire _1912_ ;
wire _9249_ ;
wire _4384_ ;
wire _823_ ;
wire _403_ ;
wire _5589_ ;
wire _5169_ ;
wire _83_ ;
wire _6950_ ;
wire _6530_ ;
wire _6110_ ;
wire _1089_ ;
wire _7735_ ;
wire _7315_ ;
wire _2870_ ;
wire _2450_ ;
wire _2030_ ;
wire _3655_ ;
wire _3235_ ;
wire _5801_ ;
wire _8693_ ;
wire _8273_ ;
wire _1721_ ;
wire _1301_ ;
wire _9058_ ;
wire _595__bF$buf0 ;
wire _4193_ ;
wire _595__bF$buf1 ;
wire _595__bF$buf2 ;
wire _595__bF$buf3 ;
wire _595__bF$buf4 ;
wire _632_ ;
wire _212_ ;
wire _2926_ ;
wire _2506_ ;
wire _5398_ ;
wire _7964_ ;
wire _7544_ ;
wire _7124_ ;
wire \datapath.idinstr_18_bF$buf4  ;
wire _8749_ ;
wire _8329_ ;
wire _3884_ ;
wire _3464_ ;
wire _3044_ ;
wire _4669_ ;
wire _4249_ ;
wire _5610_ ;
wire _8082_ ;
wire \datapath.pcstall_bF$buf3  ;
wire _6815_ ;
wire _1950_ ;
wire _1530_ ;
wire _1110_ ;
wire _9287_ ;
wire _861_ ;
wire _441_ ;
wire _2735_ ;
wire _2315_ ;
wire _7773_ ;
wire _7353_ ;
wire \datapath.idinstr_22_bF$buf4  ;
wire _8978_ ;
wire _8558_ ;
wire _8138_ ;
wire _3693_ ;
wire _3273_ ;
wire _4898_ ;
wire _4478_ ;
wire _4058_ ;
wire _917_ ;
wire _6624_ ;
wire _6204_ ;
wire _9096_ ;
wire _670_ ;
wire [31:0] _250_ ;
wire _7829_ ;
wire _7409_ ;
wire _2964_ ;
wire _2544_ ;
wire _2124_ ;
wire _3749_ ;
wire _3329_ ;
wire _7582_ ;
wire _7162_ ;
wire _8787_ ;
wire _8367_ ;
wire _3082_ ;
wire _1815_ ;
wire _4287_ ;
wire _726_ ;
wire _306_ ;
wire _6853_ ;
wire _6433_ ;
wire _6013_ ;
wire \datapath.idinstr_22_bF$buf15  ;
wire _7638_ ;
wire _7218_ ;
wire _2773_ ;
wire _2353_ ;
wire _3978_ ;
wire _3558_ ;
wire _3138_ ;
wire _7391_ ;
wire _5704_ ;
wire _8596_ ;
wire _8176_ ;
wire _6909_ ;
wire _1624_ ;
wire _1204_ ;
wire _4096_ ;
wire \datapath.idinstr_20_bF$buf35  ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _2829_ ;
wire _2409_ ;
wire _6662_ ;
wire _6242_ ;
wire _7867_ ;
wire _7447_ ;
wire _7027_ ;
wire _2582_ ;
wire _2162_ ;
wire _3787_ ;
wire _3367_ ;
wire \datapath.idinstr_17_bF$buf29  ;
wire \datapath.idinstr_21_bF$buf44  ;
wire _5933_ ;
wire _5513_ ;
wire _6718_ ;
wire \datapath.alu.b_0_bF$buf5  ;
wire _1853_ ;
wire _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _2638_ ;
wire _2218_ ;
wire _6891_ ;
wire _6471_ ;
wire _6051_ ;
wire \datapath.idinstr_15_bF$buf49  ;
wire _7676_ ;
wire _7256_ ;
wire _2391_ ;
wire _3596_ ;
wire _3176_ ;
wire _9402_ ;
wire _1909_ ;
wire _5742_ ;
wire _5322_ ;
wire _6947_ ;
wire _6527_ ;
wire _6107_ ;
wire _1662_ ;
wire _1242_ ;
wire _4060__bF$buf0 ;
wire _4060__bF$buf1 ;
wire _4060__bF$buf2 ;
wire _4060__bF$buf3 ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _2867_ ;
wire _2447_ ;
wire _2027_ ;
wire _6280_ ;
wire _7485_ ;
wire _7065_ ;
wire _9211_ ;
wire _1718_ ;
wire \datapath.idinstr_21_hier0_bF$buf0  ;
wire _5971_ ;
wire _5551_ ;
wire _5131_ ;
wire _629_ ;
wire _209_ ;
wire _6756_ ;
wire _6336_ ;
wire _1891_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _2676_ ;
wire _2256_ ;
wire _8902_ ;
wire _4822_ ;
wire _4402_ ;
wire _7294_ ;
wire _5607_ ;
wire _8499_ ;
wire _8079_ ;
wire _9440_ ;
wire _9020_ ;
wire _1947_ ;
wire _1527_ ;
wire _1107_ ;
wire _5780_ ;
wire _5360_ ;
wire _858_ ;
wire _438_ ;
wire _6985_ ;
wire _6565_ ;
wire _6145_ ;
wire _1280_ ;
wire _191_ ;
wire _2485_ ;
wire _2065_ ;
wire _8711_ ;
wire _4631_ ;
wire _4211_ ;
wire _5836_ ;
wire _5416_ ;
wire _1756_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _3902_ ;
wire _6794_ ;
wire _6374_ ;
wire _7999_ ;
wire _7579_ ;
wire _7159_ ;
wire _2294_ ;
wire _8940_ ;
wire _8520_ ;
wire _8100_ ;
wire _3499_ ;
wire _3079_ ;
wire _9305_ ;
wire _4860_ ;
wire _4440_ ;
wire _4020_ ;
wire _5645_ ;
wire _5225_ ;
wire _1985_ ;
wire _1565_ ;
wire _1145_ ;
wire _896_ ;
wire _476_ ;
wire [2:0] \datapath.memexecptions  ;
wire _3711_ ;
wire _6183_ ;
wire _4916_ ;
wire _7388_ ;
wire _9114_ ;
wire _5874_ ;
wire _5454_ ;
wire _5034_ ;
wire [31:0] \datapath.alupc_4  ;
wire _6659_ ;
wire _6239_ ;
wire _1794_ ;
wire _1374_ ;
wire _7600_ ;
wire _285_ ;
wire _2999_ ;
wire _2579_ ;
wire _2159_ ;
wire _8805_ ;
wire _3940_ ;
wire _3520_ ;
wire _3100_ ;
wire [31:0] _1_ ;
wire _4725_ ;
wire _4305_ ;
wire _7197_ ;
wire _9343_ ;
wire _5683_ ;
wire _5263_ ;
wire [2:0] bbpsel ;
wire _6888_ ;
wire _6468_ ;
wire _6048_ ;
wire _1183_ ;
wire _2388_ ;
wire _8614_ ;
wire _4954_ ;
wire _4534_ ;
wire _4114_ ;
wire _5739_ ;
wire _5319_ ;
wire _9152_ ;
wire _1659_ ;
wire _1239_ ;
wire _2600_ ;
wire _5492_ ;
wire _5072_ ;
wire CLK_bF$buf110 ;
wire CLK_bF$buf111 ;
wire CLK_bF$buf112 ;
wire CLK_bF$buf113 ;
wire CLK_bF$buf114 ;
wire CLK_bF$buf115 ;
wire \datapath.idinstr_15_bF$buf11  ;
wire CLK_bF$buf116 ;
wire CLK_bF$buf117 ;
wire CLK_bF$buf118 ;
wire _3805_ ;
wire CLK_bF$buf119 ;
wire _6697_ ;
wire _6277_ ;
wire _2197_ ;
wire _8843_ ;
wire _8423_ ;
wire _8003_ ;
wire _9208_ ;
wire _4763_ ;
wire _4343_ ;
wire _5968_ ;
wire _5548_ ;
wire _5128_ ;
wire \datapath.idinstr_16_bF$buf20  ;
wire _42_ ;
wire _9381_ ;
wire _1888_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _3614_ ;
wire _6086_ ;
wire _2799__bF$buf0 ;
wire _2799__bF$buf1 ;
wire _2799__bF$buf2 ;
wire _4819_ ;
wire _2799__bF$buf3 ;
wire _8652_ ;
wire _8232_ ;
wire _9437_ ;
wire _9017_ ;
wire _4992_ ;
wire _4572_ ;
wire _4152_ ;
wire _5777_ ;
wire _5357_ ;
wire _9190_ ;
wire _1697_ ;
wire _1277_ ;
wire _7923_ ;
wire _7503_ ;
wire _188_ ;
wire _8708_ ;
wire _3843_ ;
wire _3423_ ;
wire _3003_ ;
wire _4628_ ;
wire _4208_ ;
wire _8881_ ;
wire _8461_ ;
wire _8041_ ;
wire \datapath.idinstr_16_hier0_bF$buf4  ;
wire _9246_ ;
wire _4381_ ;
wire _820_ ;
wire _400_ ;
wire _5586_ ;
wire _5166_ ;
wire _80_ ;
wire _1086_ ;
wire _7732_ ;
wire _7312_ ;
wire _8937_ ;
wire _8517_ ;
wire _3652_ ;
wire _3232_ ;
wire _4857_ ;
wire _4437_ ;
wire _4017_ ;
wire [31:0] \datapath._28_  ;
wire _8690_ ;
wire _8270_ ;
wire _9055_ ;
wire _4190_ ;
wire _2923_ ;
wire _2503_ ;
wire _5395_ ;
wire _3708_ ;
wire _7961_ ;
wire _7541_ ;
wire _7121_ ;
wire \datapath.idinstr_18_bF$buf1  ;
wire _8746_ ;
wire _8326_ ;
wire _3881_ ;
wire _3461_ ;
wire _3041_ ;
wire _4666_ ;
wire _4246_ ;
wire \datapath.pcstall_bF$buf0  ;
wire _6812_ ;
wire _9284_ ;
wire _2732_ ;
wire _2312_ ;
wire _3937_ ;
wire _3517_ ;
wire _7770_ ;
wire _7350_ ;
wire \datapath.idinstr_22_bF$buf1  ;
wire \datapath.idinstr_16_bF$buf8  ;
wire _8975_ ;
wire _8555_ ;
wire _8135_ ;
wire _3690_ ;
wire _3270_ ;
wire _4895_ ;
wire _4475_ ;
wire _4055_ ;
wire _914_ ;
wire _6621_ ;
wire _6201_ ;
wire _9093_ ;
wire _7826_ ;
wire _7406_ ;
wire _2961_ ;
wire _2541_ ;
wire _2121_ ;
wire [31:0] \datapath.registers.1226[24]  ;
wire _3746_ ;
wire _3326_ ;
wire \datapath.idinstr_20_bF$buf8  ;
wire _8784_ ;
wire _8364_ ;
wire _1812_ ;
wire _9149_ ;
wire _4284_ ;
wire _723_ ;
wire _303_ ;
wire _5489_ ;
wire _5069_ ;
wire _6850_ ;
wire _6430_ ;
wire _6010_ ;
wire \datapath.idinstr_22_bF$buf12  ;
wire _7635_ ;
wire _7215_ ;
wire _2770_ ;
wire _2350_ ;
wire _3975_ ;
wire _3555_ ;
wire _3135_ ;
wire _5701_ ;
wire _8593_ ;
wire _8173_ ;
wire \datapath.idinstr_16_bF$buf17  ;
wire _39_ ;
wire _6906_ ;
wire _9211__bF$buf0 ;
wire _9211__bF$buf1 ;
wire _9211__bF$buf2 ;
wire _1621_ ;
wire _9211__bF$buf3 ;
wire _1201_ ;
wire _9211__bF$buf4 ;
wire _9211__bF$buf5 ;
wire _9211__bF$buf6 ;
wire _9378_ ;
wire _9211__bF$buf7 ;
wire _9211__bF$buf8 ;
wire _4093_ ;
wire \datapath.idinstr_20_bF$buf32  ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _2826_ ;
wire _2406_ ;
wire \controlunit.csrfile_wen  ;
wire _5298_ ;
wire [31:0] \datapath.regcsralu  ;
wire _7864_ ;
wire _7444_ ;
wire _7024_ ;
wire _8649_ ;
wire _8229_ ;
wire _3784_ ;
wire _3364_ ;
wire \datapath.idinstr_17_bF$buf26  ;
wire _4989_ ;
wire _4569_ ;
wire \datapath.idinstr_21_bF$buf41  ;
wire _4149_ ;
wire _5930_ ;
wire _5510_ ;
wire _6715_ ;
wire \datapath.alu.b_0_bF$buf2  ;
wire _1850_ ;
wire _1430_ ;
wire _1010_ ;
wire _9187_ ;
wire _761_ ;
wire _341_ ;
wire _2635_ ;
wire _2215_ ;
wire \datapath.idinstr_15_bF$buf46  ;
wire _7673_ ;
wire _7253_ ;
wire _8878_ ;
wire _8458_ ;
wire _8038_ ;
wire _3593_ ;
wire _3173_ ;
wire _1906_ ;
wire _4798_ ;
wire _4378_ ;
wire _817_ ;
wire _77_ ;
wire _6944_ ;
wire _6524_ ;
wire _6104_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _7729_ ;
wire _7309_ ;
wire _2864_ ;
wire _2444_ ;
wire _2024_ ;
wire _3649_ ;
wire _3229_ ;
wire _7482_ ;
wire _7062_ ;
wire _8687_ ;
wire _8267_ ;
wire _1715_ ;
wire _4187_ ;
wire _626_ ;
wire _206_ ;
wire _6753_ ;
wire _6333_ ;
wire _5456__bF$buf0 ;
wire _5456__bF$buf1 ;
wire _5456__bF$buf2 ;
wire _5456__bF$buf3 ;
wire _5456__bF$buf4 ;
wire _7958_ ;
wire _7538_ ;
wire _7118_ ;
wire _2673_ ;
wire _2253_ ;
wire _3878_ ;
wire _3458_ ;
wire _3038_ ;
wire _7291_ ;
wire _5604_ ;
wire _8496_ ;
wire _8076_ ;
wire \datapath.regcsrtrap_bF$buf6  ;
wire _6809_ ;
wire _1944_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire _2729_ ;
wire _2309_ ;
wire _5460__bF$buf0 ;
wire _5460__bF$buf1 ;
wire _5460__bF$buf2 ;
wire _5460__bF$buf3 ;
wire _5460__bF$buf4 ;
wire _6982_ ;
wire _6562_ ;
wire _6142_ ;
wire \datapath.alu.b_3_bF$buf5  ;
wire _7767_ ;
wire _7347_ ;
wire _2482_ ;
wire _2062_ ;
wire _3687_ ;
wire _3267_ ;
wire _5833_ ;
wire _5413_ ;
wire _6618_ ;
wire _1753_ ;
wire _1333_ ;
wire _664_ ;
wire _244_ ;
wire _2958_ ;
wire _2538_ ;
wire _2118_ ;
wire _6791_ ;
wire _6371_ ;
wire _7996_ ;
wire _7576_ ;
wire _7156_ ;
wire _2291_ ;
wire _3496_ ;
wire _3076_ ;
wire _9302_ ;
wire _1809_ ;
wire _5642_ ;
wire _5222_ ;
wire _6847_ ;
wire _6427_ ;
wire _6007_ ;
wire _1982_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _2767_ ;
wire _2347_ ;
wire _6180_ ;
wire _4913_ ;
wire _7385_ ;
wire _9111_ ;
wire _1618_ ;
wire _5871_ ;
wire _5451_ ;
wire _5031_ ;
wire \datapath.idinstr_20_bF$buf29  ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _6656_ ;
wire _6236_ ;
wire _1791_ ;
wire _1371_ ;
wire _282_ ;
wire _2996_ ;
wire _2576_ ;
wire _2156_ ;
wire _8802_ ;
wire _4722_ ;
wire _4302_ ;
wire _7194_ ;
wire \datapath.idinstr_21_bF$buf38  ;
wire _5927_ ;
wire _5507_ ;
wire _8399_ ;
wire _9340_ ;
wire _1847_ ;
wire _1427_ ;
wire _1007_ ;
wire _5680_ ;
wire _5260_ ;
wire _758_ ;
wire _338_ ;
wire _6885_ ;
wire _6465_ ;
wire _6045_ ;
wire _1180_ ;
wire \datapath.idinstr_22_hier0_bF$buf4  ;
wire _2385_ ;
wire _8611_ ;
wire _4951_ ;
wire _4531_ ;
wire _4111_ ;
wire _5736_ ;
wire _5316_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _3802_ ;
wire _6694_ ;
wire _6274_ ;
wire _7899_ ;
wire _7479_ ;
wire _7059_ ;
wire _2194_ ;
wire _8840_ ;
wire _8420_ ;
wire _8000_ ;
wire _3399_ ;
wire _9205_ ;
wire _4760_ ;
wire _4340_ ;
wire _5965_ ;
wire _5545_ ;
wire _5125_ ;
wire _1885_ ;
wire _1465_ ;
wire _1045_ ;
wire _796_ ;
wire _376_ ;
wire _3611_ ;
wire _6083_ ;
wire _4816_ ;
wire _7288_ ;
wire _9434_ ;
wire _9014_ ;
wire _5774_ ;
wire _5354_ ;
wire CLK_bF$buf0 ;
wire CLK_bF$buf1 ;
wire CLK_bF$buf2 ;
wire CLK_bF$buf3 ;
wire CLK_bF$buf4 ;
wire CLK_bF$buf5 ;
wire CLK_bF$buf6 ;
wire CLK_bF$buf7 ;
wire CLK_bF$buf8 ;
wire CLK_bF$buf9 ;
wire _6979_ ;
wire _6559_ ;
wire _6139_ ;
wire _1694_ ;
wire _1274_ ;
wire _7920_ ;
wire _7500_ ;
wire _185_ ;
wire _2899_ ;
wire _2479_ ;
wire _2059_ ;
wire _8705_ ;
wire _3840_ ;
wire _3420_ ;
wire _3000_ ;
wire _4625_ ;
wire _4205_ ;
wire _7097_ ;
wire \datapath.idinstr_16_hier0_bF$buf1  ;
wire _9243_ ;
wire _5583_ ;
wire _5163_ ;
wire _6788_ ;
wire _6368_ ;
wire _1083_ ;
wire _2288_ ;
wire _8934_ ;
wire _8514_ ;
wire _4854_ ;
wire _4434_ ;
wire _4014_ ;
wire _5639_ ;
wire _5219_ ;
wire _9052_ ;
wire _1979_ ;
wire _1559_ ;
wire _1139_ ;
wire _2920_ ;
wire _2500_ ;
wire _5392_ ;
wire _3705_ ;
wire _6597_ ;
wire _6177_ ;
wire _2097_ ;
wire _8743_ ;
wire _8323_ ;
wire _9108_ ;
wire _4663_ ;
wire _4243_ ;
wire _5868_ ;
wire _5448_ ;
wire _5028_ ;
wire _9281_ ;
wire _1788_ ;
wire _1368_ ;
wire _699_ ;
wire _279_ ;
wire _3934_ ;
wire _3514_ ;
wire _4719_ ;
wire \datapath.idinstr_16_bF$buf5  ;
wire _8972_ ;
wire _8552_ ;
wire _8132_ ;
wire _609__bF$buf0 ;
wire _609__bF$buf1 ;
wire _9337_ ;
wire _609__bF$buf2 ;
wire _609__bF$buf3 ;
wire _609__bF$buf4 ;
wire _4892_ ;
wire _4472_ ;
wire _4052_ ;
wire _911_ ;
wire _5677_ ;
wire _5257_ ;
wire _9090_ ;
wire _1597_ ;
wire _1177_ ;
wire _7823_ ;
wire _7403_ ;
wire _8608_ ;
wire _3743_ ;
wire _3323_ ;
wire _4948_ ;
wire \datapath.idinstr_20_bF$buf5  ;
wire _4528_ ;
wire _4108_ ;
wire _8781_ ;
wire _8361_ ;
wire _9146_ ;
wire _4281_ ;
wire _720_ ;
wire _300_ ;
wire _5486_ ;
wire _5066_ ;
wire _7632_ ;
wire _7212_ ;
wire _8837_ ;
wire _8417_ ;
wire _3972_ ;
wire _3552_ ;
wire _3132_ ;
wire _4757_ ;
wire _4337_ ;
wire _8590_ ;
wire _8170_ ;
wire \datapath.idinstr_16_bF$buf14  ;
wire _36_ ;
wire _6903_ ;
wire _9375_ ;
wire _4090_ ;
wire _2823_ ;
wire _2403_ ;
wire _5295_ ;
wire _3608_ ;
wire _7861_ ;
wire _7441_ ;
wire _7021_ ;
wire _8646_ ;
wire _8226_ ;
wire _3781_ ;
wire _3361_ ;
wire \datapath.idinstr_17_bF$buf23  ;
wire _964__bF$buf0 ;
wire _964__bF$buf1 ;
wire _964__bF$buf2 ;
wire _964__bF$buf3 ;
wire _964__bF$buf4 ;
wire _4986_ ;
wire _4566_ ;
wire _4146_ ;
wire _6712_ ;
wire _9184_ ;
wire _7917_ ;
wire _2632_ ;
wire _2212_ ;
wire \datapath.idinstr_15_bF$buf43  ;
wire _3837_ ;
wire _3417_ ;
wire _7670_ ;
wire _7250_ ;
wire _8875_ ;
wire _8455_ ;
wire _8035_ ;
wire _3590_ ;
wire _3170_ ;
wire _254__bF$buf0 ;
wire _254__bF$buf1 ;
wire _254__bF$buf2 ;
wire _254__bF$buf3 ;
wire _254__bF$buf4 ;
wire _1903_ ;
wire _4795_ ;
wire _4375_ ;
wire _814_ ;
wire _74_ ;
wire _6941_ ;
wire _6521_ ;
wire _6101_ ;
wire _7726_ ;
wire _7306_ ;
wire _2861_ ;
wire _2441_ ;
wire _2021_ ;
wire [31:0] \datapath.registers.1226[14]  ;
wire _3646_ ;
wire _3226_ ;
wire _5893__bF$buf0 ;
wire _5893__bF$buf1 ;
wire _5893__bF$buf2 ;
wire _5893__bF$buf3 ;
wire _5893__bF$buf4 ;
wire _8684_ ;
wire _8264_ ;
wire _1712_ ;
wire _9049_ ;
wire _4184_ ;
wire _623_ ;
wire _203_ ;
wire _2917_ ;
wire _5389_ ;
wire _6750_ ;
wire _6330_ ;
wire _7955_ ;
wire _7535_ ;
wire _7115_ ;
wire _2670_ ;
wire _2250_ ;
wire _3875_ ;
wire _3455_ ;
wire _2869__bF$buf0 ;
wire _3035_ ;
wire _2869__bF$buf1 ;
wire _2869__bF$buf2 ;
wire _2869__bF$buf3 ;
wire _5601_ ;
wire _8493_ ;
wire _8073_ ;
wire \datapath.regcsrtrap_bF$buf3  ;
wire _6806_ ;
wire _1941_ ;
wire _1521_ ;
wire _1101_ ;
wire _9278_ ;
wire _852_ ;
wire _432_ ;
wire _2726_ ;
wire _2306_ ;
wire _5198_ ;
wire \datapath.alu.b_3_bF$buf2  ;
wire _7764_ ;
wire _7344_ ;
wire _8969_ ;
wire _8549_ ;
wire _8129_ ;
wire _3684_ ;
wire _3264_ ;
wire _4889_ ;
wire _4469_ ;
wire _4049_ ;
wire _5830_ ;
wire _5410_ ;
wire _908_ ;
wire _6615_ ;
wire _1750_ ;
wire _1330_ ;
wire _9087_ ;
wire _661_ ;
wire _241_ ;
wire _2955_ ;
wire _2535_ ;
wire _2115_ ;
wire _7993_ ;
wire _7573_ ;
wire _7153_ ;
wire _8778_ ;
wire _8358_ ;
wire _3493_ ;
wire _3073_ ;
wire _1806_ ;
wire _4698_ ;
wire _4278_ ;
wire _717_ ;
wire _6844_ ;
wire _6424_ ;
wire _6004_ ;
wire _890_ ;
wire _470_ ;
wire _7629_ ;
wire _7209_ ;
wire _2764_ ;
wire _2344_ ;
wire _3969_ ;
wire _3549_ ;
wire _3129_ ;
wire _4910_ ;
wire _7382_ ;
wire _8587_ ;
wire _8167_ ;
wire _1615_ ;
wire _4087_ ;
wire \datapath.idinstr_20_bF$buf26  ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _6653_ ;
wire _6233_ ;
wire _7858_ ;
wire _7438_ ;
wire _7018_ ;
wire _2993_ ;
wire _2573_ ;
wire _2153_ ;
wire _3778_ ;
wire _3358_ ;
wire _979__bF$buf0 ;
wire _979__bF$buf1 ;
wire _979__bF$buf2 ;
wire _979__bF$buf3 ;
wire _979__bF$buf4 ;
wire _7191_ ;
wire \datapath.idinstr_21_bF$buf35  ;
wire _5924_ ;
wire _5504_ ;
wire _8396_ ;
wire _6709_ ;
wire _1844_ ;
wire _1424_ ;
wire _1004_ ;
wire _755_ ;
wire _335_ ;
wire _2629_ ;
wire _2209_ ;
wire _6882_ ;
wire _6462_ ;
wire _6042_ ;
wire \datapath.idinstr_22_hier0_bF$buf1  ;
wire _7667_ ;
wire _7247_ ;
wire _2382_ ;
wire _3587_ ;
wire _3167_ ;
wire _5733_ ;
wire _5313_ ;
wire _6938_ ;
wire _6518_ ;
wire _1653_ ;
wire _1233_ ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _2858_ ;
wire _2438_ ;
wire _2018_ ;
wire _6691_ ;
wire _6271_ ;
wire _7896_ ;
wire _7476_ ;
wire _7056_ ;
wire _2191_ ;
wire _3396_ ;
wire _9202_ ;
wire _1709_ ;
wire _5962_ ;
wire _5542_ ;
wire _5122_ ;
wire _6747_ ;
wire _6327_ ;
wire _1882_ ;
wire _1462_ ;
wire _1042_ ;
wire _793_ ;
wire _373_ ;
wire _2667_ ;
wire _2247_ ;
wire _6080_ ;
wire _4813_ ;
wire _7285_ ;
wire _9431_ ;
wire _9011_ ;
wire _1938_ ;
wire _1518_ ;
wire _5771_ ;
wire _5351_ ;
wire _849_ ;
wire _429_ ;
wire _6976_ ;
wire _6556_ ;
wire _6136_ ;
wire _1691_ ;
wire _1271_ ;
wire _182_ ;
wire _2896_ ;
wire _2476_ ;
wire _2056_ ;
wire _8702_ ;
wire _4622_ ;
wire _4202_ ;
wire _7094_ ;
wire _5827_ ;
wire _5407_ ;
wire _7610__bF$buf0 ;
wire _7610__bF$buf1 ;
wire _7610__bF$buf2 ;
wire _7610__bF$buf3 ;
wire _7610__bF$buf4 ;
wire _8299_ ;
wire _9240_ ;
wire _1747_ ;
wire _1327_ ;
wire _5580_ ;
wire _5160_ ;
wire _658_ ;
wire _238_ ;
wire _6785_ ;
wire _6365_ ;
wire _1080_ ;
wire _2285_ ;
wire _8931_ ;
wire _8511_ ;
wire _4851_ ;
wire _4431_ ;
wire _4011_ ;
wire _5636_ ;
wire _5216_ ;
wire _1976_ ;
wire _1556_ ;
wire _1136_ ;
wire _887_ ;
wire _467_ ;
wire _3702_ ;
wire _6594_ ;
wire _6174_ ;
wire _4907_ ;
wire _7799_ ;
wire _7379_ ;
wire _2094_ ;
wire _8740_ ;
wire _8320_ ;
wire _3299_ ;
wire _9105_ ;
wire _4660_ ;
wire _4240_ ;
wire _5865_ ;
wire _5445_ ;
wire _5025_ ;
wire [31:0] \datapath.idpc  ;
wire _1785_ ;
wire _1365_ ;
wire _696_ ;
wire _276_ ;
wire _3931_ ;
wire _3511_ ;
wire _4716_ ;
wire _7188_ ;
wire \datapath.idinstr_16_bF$buf2  ;
wire _9334_ ;
wire _5674_ ;
wire _5254_ ;
wire _6879_ ;
wire _6459_ ;
wire _6039_ ;
wire _1594_ ;
wire _1174_ ;
wire _7820_ ;
wire _7400_ ;
wire _2799_ ;
wire _2379_ ;
wire _8605_ ;
wire _3740_ ;
wire _3320_ ;
wire _4945_ ;
wire \datapath.idinstr_20_bF$buf2  ;
wire _4525_ ;
wire _4105_ ;
wire [1:0] \datapath.regpcsel  ;
wire _9143_ ;
wire _5483_ ;
wire _5063_ ;
wire _6688_ ;
wire _6268_ ;
wire _2188_ ;
wire _8834_ ;
wire _8414_ ;
wire _4754_ ;
wire _4334_ ;
wire _5959_ ;
wire _5539_ ;
wire _5119_ ;
wire \datapath.idinstr_16_bF$buf11  ;
wire _33_ ;
wire _6900_ ;
wire _9372_ ;
wire _1879_ ;
wire _1459_ ;
wire _1039_ ;
wire _2820_ ;
wire _2400_ ;
wire _5292_ ;
wire \datapath.idinstr_17_hier0_bF$buf5  ;
wire _3605_ ;
wire _6497_ ;
wire _6077_ ;
wire _8643_ ;
wire _8223_ ;
wire \datapath.idinstr_17_bF$buf20  ;
wire _9428_ ;
wire _9008_ ;
wire _4983_ ;
wire _4563_ ;
wire _4143_ ;
wire \datapath.idinstr_19_bF$buf5  ;
wire _5768_ ;
wire _5348_ ;
wire _9181_ ;
wire _1688_ ;
wire _1268_ ;
wire _7914_ ;
wire _599_ ;
wire _179_ ;
wire \datapath.idinstr_15_bF$buf40  ;
wire _3834_ ;
wire _3414_ ;
wire _4619_ ;
wire _8872_ ;
wire _8452_ ;
wire _8032_ ;
wire _1900_ ;
wire _9237_ ;
wire _4792_ ;
wire _4372_ ;
wire \datapath.idinstr_23_bF$buf5  ;
wire _811_ ;
wire _5997_ ;
wire _5577_ ;
wire _5157_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _7723_ ;
wire _7303_ ;
wire _8928_ ;
wire _8508_ ;
wire _3643_ ;
wire _3223_ ;
wire _4848_ ;
wire _4428_ ;
wire _4008_ ;
wire _8681_ ;
wire _8261_ ;
wire [31:0] \datapath.csr.csr_data  ;
wire _9046_ ;
wire _4181_ ;
wire _620_ ;
wire _200_ ;
wire _2914_ ;
wire _5386_ ;
wire _7952_ ;
wire _7532_ ;
wire _7112_ ;
wire _8737_ ;
wire _8317_ ;
wire _3872_ ;
wire _3452_ ;
wire _3032_ ;
wire _4657_ ;
wire _4237_ ;
wire _8490_ ;
wire _8070_ ;
wire \datapath.regcsrtrap_bF$buf0  ;
wire _6803_ ;
wire _9275_ ;
wire _5545__bF$buf0 ;
wire _5545__bF$buf1 ;
wire _5545__bF$buf2 ;
wire _5545__bF$buf3 ;
wire _5545__bF$buf4 ;
wire _2723_ ;
wire _2303_ ;
wire _5195_ ;
wire _3928_ ;
wire _3508_ ;
wire _7761_ ;
wire _7341_ ;
wire \bypassandflushunit.stall  ;
wire _8966_ ;
wire _8546_ ;
wire _8126_ ;
wire _3681_ ;
wire _3261_ ;
wire _4886_ ;
wire _4466_ ;
wire _4046_ ;
wire _905_ ;
wire _6612_ ;
wire _9084_ ;
wire _7817_ ;
wire _2952_ ;
wire _2532_ ;
wire _2112_ ;
wire _3737_ ;
wire _3317_ ;
wire \datapath.alu.b_1_bF$buf6  ;
wire _7990_ ;
wire _7570_ ;
wire _7150_ ;
wire _8775_ ;
wire _8355_ ;
wire _3490_ ;
wire _3070_ ;
wire _1803_ ;
wire _4695_ ;
wire _4275_ ;
wire _714_ ;
wire _6841_ ;
wire _6421_ ;
wire _6001_ ;
wire [31:0] \datapath.alu.c  ;
wire _7626_ ;
wire _7206_ ;
wire _2761_ ;
wire _2341_ ;
wire _3966_ ;
wire _3546_ ;
wire _3126_ ;
wire _8584_ ;
wire _8164_ ;
wire _1612_ ;
wire _9369_ ;
wire _4084_ ;
wire \datapath.idinstr_20_bF$buf23  ;
wire _943_ ;
wire _523_ ;
wire _103_ ;
wire _2817_ ;
wire _5289_ ;
wire _6650_ ;
wire _6230_ ;
wire _7855_ ;
wire _7435_ ;
wire _7015_ ;
wire _2990_ ;
wire _2570_ ;
wire _2150_ ;
wire _3775_ ;
wire _3355_ ;
wire \datapath.idinstr_17_bF$buf17  ;
wire _9075__bF$buf0 ;
wire _9075__bF$buf1 ;
wire _9075__bF$buf2 ;
wire _9075__bF$buf3 ;
wire _9075__bF$buf4 ;
wire \datapath.idinstr_21_bF$buf32  ;
wire _5921_ ;
wire _5501_ ;
wire _8393_ ;
wire _6706_ ;
wire _1841_ ;
wire _1421_ ;
wire _1001_ ;
wire _9178_ ;
wire _752_ ;
wire _332_ ;
wire _2626_ ;
wire _2206_ ;
wire _5098_ ;
wire \datapath.idinstr_15_bF$buf37  ;
wire \datapath.idinstr_22_bF$buf41  ;
wire _7664_ ;
wire _7244_ ;
wire [31:0] \datapath.registers.1226[5]  ;
wire _8869_ ;
wire _8449_ ;
wire _8029_ ;
wire _3584_ ;
wire _3164_ ;
wire _4789_ ;
wire _4369_ ;
wire _5730_ ;
wire _5310_ ;
wire _808_ ;
wire _68_ ;
wire _6935_ ;
wire _6515_ ;
wire _1650_ ;
wire _1230_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _2855_ ;
wire _2435_ ;
wire _2015_ ;
wire _7893_ ;
wire _7473_ ;
wire _7053_ ;
wire _8678_ ;
wire _8258_ ;
wire _3393_ ;
wire _1706_ ;
wire _4598_ ;
wire _4178_ ;
wire _617_ ;
wire _6744_ ;
wire _6324_ ;
wire _790_ ;
wire _370_ ;
wire _7949_ ;
wire _7529_ ;
wire _7109_ ;
wire _2664_ ;
wire _2244_ ;
wire _3869_ ;
wire _3449_ ;
wire _3029_ ;
wire _4810_ ;
wire _7282_ ;
wire _8487_ ;
wire _8067_ ;
wire _5466__bF$buf0 ;
wire _5466__bF$buf1 ;
wire _5466__bF$buf2 ;
wire _5466__bF$buf3 ;
wire _5466__bF$buf4 ;
wire _1935_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _6973_ ;
wire _6553_ ;
wire _6133_ ;
wire _7758_ ;
wire _7338_ ;
wire _2893_ ;
wire _2473_ ;
wire _2053_ ;
wire _3678_ ;
wire _3258_ ;
wire _7091_ ;
wire _5824_ ;
wire _5404_ ;
wire _8296_ ;
wire _5470__bF$buf0 ;
wire _5470__bF$buf1 ;
wire _5470__bF$buf2 ;
wire _5470__bF$buf3 ;
wire _5470__bF$buf4 ;
wire _6609_ ;
wire _1744_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _2949_ ;
wire _2529_ ;
wire _2109_ ;
wire _6782_ ;
wire _6362_ ;
wire _7987_ ;
wire _7567_ ;
wire _7147_ ;
wire _2282_ ;
wire _3487_ ;
wire _3067_ ;
wire _5633_ ;
wire _5213_ ;
wire _6838_ ;
wire _6418_ ;
wire _1973_ ;
wire _1553_ ;
wire _1133_ ;
wire _884_ ;
wire _464_ ;
wire _2758_ ;
wire _2338_ ;
wire _6591_ ;
wire _6171_ ;
wire _4904_ ;
wire _7796_ ;
wire _7376_ ;
wire _2091_ ;
wire \datapath.regz  ;
wire _3296_ ;
wire _9102_ ;
wire _1609_ ;
wire _5862_ ;
wire _5442_ ;
wire _5022_ ;
wire _6647_ ;
wire _6227_ ;
wire _1782_ ;
wire _1362_ ;
wire _693_ ;
wire _273_ ;
wire _2987_ ;
wire _9142__bF$buf0 ;
wire _2567_ ;
wire _9142__bF$buf1 ;
wire _2147_ ;
wire _9142__bF$buf2 ;
wire _9142__bF$buf3 ;
wire _9142__bF$buf4 ;
wire _4713_ ;
wire _7185_ ;
wire \datapath.idinstr_21_bF$buf29  ;
wire _5918_ ;
wire _9331_ ;
wire _1838_ ;
wire _1418_ ;
wire _5671_ ;
wire _5251_ ;
wire _749_ ;
wire _329_ ;
wire _6876_ ;
wire _6456_ ;
wire _6036_ ;
wire _1591_ ;
wire _1171_ ;
wire \datapath.idinstr_22_bF$buf38  ;
wire _2796_ ;
wire _2376_ ;
wire _8602_ ;
wire _604__bF$buf0 ;
wire _604__bF$buf1 ;
wire _604__bF$buf2 ;
wire _604__bF$buf3 ;
wire _604__bF$buf4 ;
wire _4942_ ;
wire _4522_ ;
wire _4102_ ;
wire \bypassandflushunit.stall_bF$buf8  ;
wire _5727_ ;
wire _5307_ ;
wire _8199_ ;
wire _9140_ ;
wire _1647_ ;
wire _1227_ ;
wire _5480_ ;
wire _5060_ ;
wire _978_ ;
wire _558_ ;
wire _138_ ;
wire _6685_ ;
wire _6265_ ;
wire _3267__bF$buf0 ;
wire _3267__bF$buf1 ;
wire _3267__bF$buf2 ;
wire _3267__bF$buf3 ;
wire _3267__bF$buf4 ;
wire _3267__bF$buf5 ;
wire _3267__bF$buf6 ;
wire _2185_ ;
wire _8831_ ;
wire _8411_ ;
wire _4751_ ;
wire _4331_ ;
wire _5956_ ;
wire _5536_ ;
wire _5116_ ;
wire _30_ ;
wire _1876_ ;
wire _1456_ ;
wire _1036_ ;
wire _787_ ;
wire _367_ ;
wire \datapath.idinstr_17_hier0_bF$buf2  ;
wire _3602_ ;
wire _6494_ ;
wire _6074_ ;
wire _6074__bF$buf0 ;
wire _6074__bF$buf1 ;
wire _6074__bF$buf2 ;
wire _6074__bF$buf3 ;
wire _6074__bF$buf4 ;
wire _4807_ ;
wire _7699_ ;
wire _7279_ ;
wire _8640_ ;
wire _8220_ ;
wire _3199_ ;
wire _9425_ ;
wire _9005_ ;
wire _4980_ ;
wire _4560_ ;
wire _4140_ ;
wire \datapath.idinstr_19_bF$buf2  ;
wire _5765_ ;
wire _5345_ ;
wire _1685_ ;
wire _1265_ ;
wire _7911_ ;
wire _596_ ;
wire _176_ ;
wire _3831_ ;
wire _3411_ ;
wire _4616_ ;
wire _7088_ ;
wire _9234_ ;
wire \datapath.idinstr_23_bF$buf2  ;
wire _5994_ ;
wire _5574_ ;
wire _5154_ ;
wire [31:0] \datapath.programcounter.pc_mux  ;
wire _6779_ ;
wire _6359_ ;
wire _1494_ ;
wire _1074_ ;
wire _7720_ ;
wire _7300_ ;
wire _2699_ ;
wire _2279_ ;
wire _8925_ ;
wire _8505_ ;
wire _3640_ ;
wire _3220_ ;
wire [31:0] \datapath.csr.csr_mepc  ;
wire _4845_ ;
wire _4425_ ;
wire _4005_ ;
wire _9043_ ;
wire _2911_ ;
wire _5383_ ;
wire _6588_ ;
wire _6168_ ;
wire _2088_ ;
wire _8734_ ;
wire _8314_ ;
wire _4654_ ;
wire _4234_ ;
wire _5859_ ;
wire _5439_ ;
wire _5019_ ;
wire _6800_ ;
wire _9272_ ;
wire _1779_ ;
wire _1359_ ;
wire _2720_ ;
wire _2300_ ;
wire _5192_ ;
wire _3925_ ;
wire _3505_ ;
wire _6397_ ;
wire _8963_ ;
wire _8543_ ;
wire _8123_ ;
wire _9328_ ;
wire _4883_ ;
wire _4463_ ;
wire _4043_ ;
wire _902_ ;
wire _5668_ ;
wire _5248_ ;
wire _9081_ ;
wire _1588_ ;
wire _1168_ ;
wire _7814_ ;
wire _499_ ;
wire _3734_ ;
wire _3314_ ;
wire \datapath.alu.b_1_bF$buf3  ;
wire _4939_ ;
wire _4519_ ;
wire _8772_ ;
wire _8352_ ;
wire _1800_ ;
wire _9137_ ;
wire _4692_ ;
wire _4272_ ;
wire _711_ ;
wire _5897_ ;
wire _5477_ ;
wire _5057_ ;
wire _1397_ ;
wire _7623_ ;
wire _7203_ ;
wire _8828_ ;
wire _8408_ ;
wire _3963_ ;
wire _3543_ ;
wire _3123_ ;
wire _4748_ ;
wire _4328_ ;
wire _8581_ ;
wire _8161_ ;
wire _27_ ;
wire _9366_ ;
wire _4081_ ;
wire \datapath.idinstr_20_bF$buf20  ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire _2814_ ;
wire _6141__bF$buf0 ;
wire _6141__bF$buf1 ;
wire _6141__bF$buf2 ;
wire _5286_ ;
wire _6141__bF$buf3 ;
wire _6141__bF$buf4 ;
wire _6141__bF$buf5 ;
wire _6141__bF$buf6 ;
wire _6141__bF$buf7 ;
wire _6141__bF$buf8 ;
wire _6141__bF$buf9 ;
wire _7852_ ;
wire _7432_ ;
wire _7012_ ;
wire _8637_ ;
wire _8217_ ;
wire _3772_ ;
wire _3352_ ;
wire \datapath.idinstr_17_bF$buf14  ;
wire _4977_ ;
wire _4557_ ;
wire _4137_ ;
wire _8390_ ;
wire _6703_ ;
wire _9175_ ;
wire _7908_ ;
wire _2623_ ;
wire _2203_ ;
wire _5095_ ;
wire \datapath.idinstr_15_bF$buf34  ;
wire _3828_ ;
wire _974__bF$buf0 ;
wire _3408_ ;
wire _974__bF$buf1 ;
wire _974__bF$buf2 ;
wire _974__bF$buf3 ;
wire _974__bF$buf4 ;
wire _7661_ ;
wire _7241_ ;
wire _8866_ ;
wire _8446_ ;
wire _8026_ ;
wire _3581_ ;
wire _3161_ ;
wire _4786_ ;
wire _4366_ ;
wire _805_ ;
wire \datapath.idinstr_16_bF$buf43  ;
wire _65_ ;
wire _6932_ ;
wire _6512_ ;
wire _7717_ ;
wire _2852_ ;
wire _2432_ ;
wire _2012_ ;
wire _3637_ ;
wire _3217_ ;
wire _7890_ ;
wire _7470_ ;
wire _7050_ ;
wire _8675_ ;
wire _8255_ ;
wire _3390_ ;
wire _1703_ ;
wire _4595_ ;
wire _4175_ ;
wire _614_ ;
wire _2908_ ;
wire _6741_ ;
wire _6321_ ;
wire _7946_ ;
wire _7526_ ;
wire _7106_ ;
wire _2661_ ;
wire _2241_ ;
wire _3866_ ;
wire _3446_ ;
wire _3026_ ;
wire _8484_ ;
wire _8064_ ;
wire _1932_ ;
wire _1512_ ;
wire _9269_ ;
wire _843_ ;
wire _423_ ;
wire _2717_ ;
wire _5189_ ;
wire _6970_ ;
wire _6550_ ;
wire _6130_ ;
wire _7755_ ;
wire _7335_ ;
wire _2890_ ;
wire _2470_ ;
wire _2050_ ;
wire _3675_ ;
wire _3255_ ;
wire _5821_ ;
wire _5401_ ;
wire _8293_ ;
wire _6606_ ;
wire _1741_ ;
wire _1321_ ;
wire _9078_ ;
wire _652_ ;
wire _232_ ;
wire _2946_ ;
wire _2526_ ;
wire _2106_ ;
wire _7984_ ;
wire _7564_ ;
wire _7144_ ;
wire _8769_ ;
wire _8349_ ;
wire _3484_ ;
wire _3064_ ;
wire _4689_ ;
wire _4269_ ;
wire _5630_ ;
wire _5210_ ;
wire _708_ ;
wire _6835_ ;
wire _6415_ ;
wire _1970_ ;
wire _1550_ ;
wire _1130_ ;
wire _881_ ;
wire _461_ ;
wire _2755_ ;
wire _2335_ ;
wire [3:0] alusel ;
wire _4901_ ;
wire _7793_ ;
wire _7373_ ;
wire _8998_ ;
wire _8578_ ;
wire _8158_ ;
wire _3293_ ;
wire _1606_ ;
wire _4498_ ;
wire _4078_ ;
wire \datapath.idinstr_20_bF$buf17  ;
wire _937_ ;
wire _517_ ;
wire _6644_ ;
wire _6224_ ;
wire _5615__bF$buf0 ;
wire _5615__bF$buf1 ;
wire _5615__bF$buf2 ;
wire _5615__bF$buf3 ;
wire _5615__bF$buf4 ;
wire _5615__bF$buf5 ;
wire _5615__bF$buf6 ;
wire _5615__bF$buf7 ;
wire _5615__bF$buf8 ;
wire _690_ ;
wire _270_ ;
wire _7849_ ;
wire _7429_ ;
wire _7009_ ;
wire _2984_ ;
wire _2564_ ;
wire _2144_ ;
wire _3769_ ;
wire _3349_ ;
wire _4710_ ;
wire _7182_ ;
wire \datapath.idinstr_21_bF$buf26  ;
wire _5915_ ;
wire _8387_ ;
wire _1835_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _6873_ ;
wire _6453_ ;
wire _6033_ ;
wire \datapath.idinstr_22_bF$buf35  ;
wire _7658_ ;
wire _7238_ ;
wire _2793_ ;
wire _2373_ ;
wire _3998_ ;
wire _3578_ ;
wire _3158_ ;
wire \bypassandflushunit.stall_bF$buf5  ;
wire _5724_ ;
wire _5304_ ;
wire _8196_ ;
wire _6929_ ;
wire _6509_ ;
wire _1644_ ;
wire _1224_ ;
wire \datapath.idinstr_20_bF$buf55  ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire _2849_ ;
wire _2429_ ;
wire _2009_ ;
wire _6682_ ;
wire _6262_ ;
wire _7887_ ;
wire _7467_ ;
wire _7047_ ;
wire _2182_ ;
wire _3387_ ;
wire _5953_ ;
wire _5533_ ;
wire _5113_ ;
wire DMEM_WEN ;
wire _6738_ ;
wire _6318_ ;
wire _1873_ ;
wire _1453_ ;
wire _1033_ ;
wire _784_ ;
wire _364_ ;
wire _2658_ ;
wire _2238_ ;
wire _6491_ ;
wire _6071_ ;
wire _4804_ ;
wire _7696_ ;
wire _7276_ ;
wire _3196_ ;
wire _9422_ ;
wire _9002_ ;
wire _1929_ ;
wire _1509_ ;
wire _5762_ ;
wire _5342_ ;
wire _6967_ ;
wire _6547_ ;
wire _6127_ ;
wire _1682_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _2887_ ;
wire _2467_ ;
wire _2047_ ;
wire _4613_ ;
wire _7085_ ;
wire _5818_ ;
wire _9231_ ;
wire _1738_ ;
wire _1318_ ;
wire _5991_ ;
wire _5571_ ;
wire _5151_ ;
wire _649_ ;
wire _229_ ;
wire _6776_ ;
wire _6356_ ;
wire _1491_ ;
wire _1071_ ;
wire _2696_ ;
wire _2276_ ;
wire _8922_ ;
wire _8502_ ;
wire _4842_ ;
wire _4422_ ;
wire _4002_ ;
wire _5627_ ;
wire _5207_ ;
wire _8099_ ;
wire _9040_ ;
wire _1967_ ;
wire _1547_ ;
wire _1127_ ;
wire _5380_ ;
wire _878_ ;
wire _458_ ;
wire _6585_ ;
wire _6165_ ;
wire _2085_ ;
wire _8731_ ;
wire _8311_ ;
wire _4651_ ;
wire _4231_ ;
wire _5856_ ;
wire _5436_ ;
wire _5016_ ;
wire _1776_ ;
wire _1356_ ;
wire _687_ ;
wire _267_ ;
wire _3922_ ;
wire _3502_ ;
wire _6394_ ;
wire _4707_ ;
wire _7599_ ;
wire _7179_ ;
wire _8960_ ;
wire _8540_ ;
wire _8120_ ;
wire _3099_ ;
wire _9325_ ;
wire _4880_ ;
wire _4460_ ;
wire _4040_ ;
wire _5665_ ;
wire _5245_ ;
wire \datapath.idinstr_17_bF$buf8  ;
wire _1585_ ;
wire _1165_ ;
wire _7811_ ;
wire _496_ ;
wire _3731_ ;
wire _3311_ ;
wire \datapath.alu.b_1_bF$buf0  ;
wire _4936_ ;
wire _4516_ ;
wire _9377__bF$buf0 ;
wire _9377__bF$buf1 ;
wire _9377__bF$buf2 ;
wire _9377__bF$buf3 ;
wire _9377__bF$buf4 ;
wire _9134_ ;
wire \datapath.idinstr_21_bF$buf8  ;
wire _5894_ ;
wire _5474_ ;
wire _5054_ ;
wire _5492__bF$buf0 ;
wire _5492__bF$buf1 ;
wire _5492__bF$buf2 ;
wire _5492__bF$buf3 ;
wire _5492__bF$buf4 ;
wire _6679_ ;
wire _6259_ ;
wire _1394_ ;
wire _7620_ ;
wire _7200_ ;
wire _2599_ ;
wire _2179_ ;
wire _8825_ ;
wire _8405_ ;
wire _3960_ ;
wire _3540_ ;
wire _3120_ ;
wire _4745_ ;
wire _4325_ ;
wire _24_ ;
wire _9363_ ;
wire _2811_ ;
wire _5283_ ;
wire [31:0] IMEM_DATA ;
wire _6488_ ;
wire _6068_ ;
wire _8634_ ;
wire _8214_ ;
wire \datapath.idinstr_17_bF$buf11  ;
wire _9419_ ;
wire _4974_ ;
wire _4554_ ;
wire _4134_ ;
wire [7:0] \datapath.memoryinterface.byte_size_load.byteval  ;
wire _5759_ ;
wire _5339_ ;
wire _6700_ ;
wire _9172_ ;
wire _1679_ ;
wire _1259_ ;
wire _7905_ ;
wire _2620_ ;
wire _2200_ ;
wire _5092_ ;
wire \datapath.idinstr_15_bF$buf31  ;
wire _3825_ ;
wire _3405_ ;
wire _6297_ ;
wire _9310__bF$buf0 ;
wire _9310__bF$buf1 ;
wire _9310__bF$buf2 ;
wire _9310__bF$buf3 ;
wire _9310__bF$buf4 ;
wire _9310__bF$buf5 ;
wire _9310__bF$buf6 ;
wire _9310__bF$buf7 ;
wire _8863_ ;
wire _8443_ ;
wire _8023_ ;
wire \datapath.alu.b_4_bF$buf3  ;
wire _9228_ ;
wire _4783_ ;
wire _4363_ ;
wire _802_ ;
wire _5988_ ;
wire _5568_ ;
wire _5148_ ;
wire \datapath.idinstr_16_bF$buf40  ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire _7714_ ;
wire _399_ ;
wire _8919_ ;
wire _3634_ ;
wire _3214_ ;
wire _4839_ ;
wire _4419_ ;
wire _8672_ ;
wire _8252_ ;
wire _1700_ ;
wire _9037_ ;
wire _4592_ ;
wire _4172_ ;
wire _611_ ;
wire _2905_ ;
wire _5797_ ;
wire _5377_ ;
wire _1297_ ;
wire _7943_ ;
wire _7523_ ;
wire _7103_ ;
wire _6144__bF$buf0 ;
wire _6144__bF$buf1 ;
wire _6144__bF$buf2 ;
wire _6144__bF$buf3 ;
wire _6144__bF$buf4 ;
wire _6144__bF$buf5 ;
wire _8728_ ;
wire _6144__bF$buf6 ;
wire _8308_ ;
wire _6144__bF$buf7 ;
wire _6144__bF$buf8 ;
wire _6144__bF$buf9 ;
wire _3863_ ;
wire _3443_ ;
wire _3023_ ;
wire _4648_ ;
wire _4228_ ;
wire _8481_ ;
wire CLK_bF$buf70 ;
wire _8061_ ;
wire CLK_bF$buf71 ;
wire CLK_bF$buf72 ;
wire CLK_bF$buf73 ;
wire CLK_bF$buf74 ;
wire CLK_bF$buf75 ;
wire CLK_bF$buf76 ;
wire CLK_bF$buf77 ;
wire CLK_bF$buf78 ;
wire CLK_bF$buf79 ;
wire _9266_ ;
wire _840_ ;
wire _420_ ;
wire _2714_ ;
wire _5186_ ;
wire _3919_ ;
wire _7752_ ;
wire _7332_ ;
wire _8957_ ;
wire _8537_ ;
wire _8117_ ;
wire _3672_ ;
wire _3252_ ;
wire _977__bF$buf0 ;
wire _977__bF$buf1 ;
wire _977__bF$buf2 ;
wire _977__bF$buf3 ;
wire _977__bF$buf4 ;
wire _4877_ ;
wire _4457_ ;
wire _4037_ ;
wire _8290_ ;
wire _6603_ ;
wire _9075_ ;
wire _7808_ ;
wire _2943_ ;
wire _2523_ ;
wire _2103_ ;
wire _3728_ ;
wire _3308_ ;
wire [2:0] \bypassandflushunit.rs2_bypass_sel  ;
wire _7981_ ;
wire _7561_ ;
wire _7141_ ;
wire _8766_ ;
wire _8346_ ;
wire _3481_ ;
wire _3061_ ;
wire _4686_ ;
wire _4266_ ;
wire _705_ ;
wire _6832_ ;
wire _6412_ ;
wire _7617_ ;
wire _2752_ ;
wire _2332_ ;
wire _3957_ ;
wire _3537_ ;
wire _3117_ ;
wire _7790_ ;
wire _7370_ ;
wire _8995_ ;
wire _8575_ ;
wire _8155_ ;
wire _3290_ ;
wire _1603_ ;
wire _4495_ ;
wire _4075_ ;
wire \datapath.idinstr_20_bF$buf14  ;
wire _934_ ;
wire _514_ ;
wire _2808_ ;
wire _6641_ ;
wire _6221_ ;
wire _7846_ ;
wire _7426_ ;
wire _7006_ ;
wire _2981_ ;
wire _2561_ ;
wire _2141_ ;
wire [31:0] \datapath.registers.1226[26]  ;
wire _3766_ ;
wire _3346_ ;
wire \datapath.idinstr_21_bF$buf23  ;
wire _5912_ ;
wire _8384_ ;
wire _1832_ ;
wire _1412_ ;
wire _9169_ ;
wire _743_ ;
wire _323_ ;
wire _2617_ ;
wire _5089_ ;
wire _6870_ ;
wire _6450_ ;
wire _6030_ ;
wire \datapath.idinstr_15_bF$buf28  ;
wire \datapath.csr.mip  ;
wire \datapath.idinstr_22_bF$buf32  ;
wire _7655_ ;
wire _7235_ ;
wire _2790_ ;
wire _2370_ ;
wire _3995_ ;
wire _3575_ ;
wire _3155_ ;
wire \bypassandflushunit.stall_bF$buf2  ;
wire _5721_ ;
wire _5301_ ;
wire _8193_ ;
wire branch ;
wire \datapath.idinstr_16_bF$buf37  ;
wire _59_ ;
wire _6926_ ;
wire _6506_ ;
wire _1641_ ;
wire _1221_ ;
wire _9398_ ;
wire \datapath.idinstr_20_bF$buf52  ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _2846_ ;
wire _2426_ ;
wire _2006_ ;
wire _7884_ ;
wire _7464_ ;
wire _7044_ ;
wire _8669_ ;
wire _8249_ ;
wire _3384_ ;
wire _4589_ ;
wire _4169_ ;
wire _5950_ ;
wire _5530_ ;
wire _5110_ ;
wire _608_ ;
wire _6735_ ;
wire _6315_ ;
wire _1870_ ;
wire _1450_ ;
wire _1030_ ;
wire _781_ ;
wire _361_ ;
wire _2655_ ;
wire _2235_ ;
wire _4801_ ;
wire _7693_ ;
wire _7273_ ;
wire _8898_ ;
wire _8478_ ;
wire _8058_ ;
wire _3193_ ;
wire _1926_ ;
wire _1506_ ;
wire _4398_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _6964_ ;
wire _6544_ ;
wire _6124_ ;
wire _590_ ;
wire _170_ ;
wire _7749_ ;
wire _7329_ ;
wire _2884_ ;
wire _2464_ ;
wire _2044_ ;
wire _5476__bF$buf0 ;
wire _5476__bF$buf1 ;
wire _5476__bF$buf2 ;
wire _3669_ ;
wire _5476__bF$buf3 ;
wire _3249_ ;
wire _5476__bF$buf4 ;
wire _4610_ ;
wire _7082_ ;
wire _5815_ ;
wire _8287_ ;
wire _1735_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire \datapath.alu.z  ;
wire _6773_ ;
wire _6353_ ;
wire _7978_ ;
wire _7558_ ;
wire _7138_ ;
wire _2693_ ;
wire _2273_ ;
wire _5480__bF$buf0 ;
wire _5480__bF$buf1 ;
wire _5480__bF$buf2 ;
wire _5480__bF$buf3 ;
wire _5480__bF$buf4 ;
wire _3898_ ;
wire _3478_ ;
wire _3058_ ;
wire _5624_ ;
wire _5204_ ;
wire _8096_ ;
wire _6829_ ;
wire _6409_ ;
wire _1964_ ;
wire _1544_ ;
wire _1124_ ;
wire _875_ ;
wire _455_ ;
wire _2749_ ;
wire _2329_ ;
wire _6582_ ;
wire _6162_ ;
wire _7787_ ;
wire _7367_ ;
wire _2082_ ;
wire _3287_ ;
wire _5853_ ;
wire _5433_ ;
wire _5013_ ;
wire _6638_ ;
wire _6218_ ;
wire _1773_ ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire _2978_ ;
wire _2558_ ;
wire _2138_ ;
wire _6391_ ;
wire _4704_ ;
wire _7596_ ;
wire _7176_ ;
wire _4008__bF$buf0 ;
wire _4008__bF$buf1 ;
wire _4008__bF$buf2 ;
wire _5909_ ;
wire _4008__bF$buf3 ;
wire _3096_ ;
wire _9322_ ;
wire _1829_ ;
wire _1409_ ;
wire _5662_ ;
wire _5242_ ;
wire \datapath.idinstr_17_bF$buf5  ;
wire _6867_ ;
wire _6447_ ;
wire _6027_ ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire \datapath.idinstr_22_bF$buf29  ;
wire _2787_ ;
wire _2367_ ;
wire _4933_ ;
wire _4513_ ;
wire _5718_ ;
wire _9131_ ;
wire _1638_ ;
wire _1218_ ;
wire \datapath.idinstr_21_bF$buf5  ;
wire _5891_ ;
wire _5471_ ;
wire _5051_ ;
wire \datapath.idinstr_20_bF$buf49  ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire _6676_ ;
wire _6256_ ;
wire _1391_ ;
wire _2596_ ;
wire _2176_ ;
wire _8822_ ;
wire _8402_ ;
wire _4742_ ;
wire _4322_ ;
wire _5947_ ;
wire _5527_ ;
wire _5107_ ;
wire _21_ ;
wire _9360_ ;
wire _1867_ ;
wire _1447_ ;
wire _1027_ ;
wire _5280_ ;
wire _778_ ;
wire _358_ ;
wire _6485_ ;
wire _6065_ ;
wire _8631_ ;
wire _8211_ ;
wire _9416_ ;
wire _4971_ ;
wire _4551_ ;
wire _4131_ ;
wire _5756_ ;
wire _5336_ ;
wire _1676_ ;
wire _1256_ ;
wire _7902_ ;
wire _587_ ;
wire _167_ ;
wire _3822_ ;
wire _3402_ ;
wire _2688__bF$buf0 ;
wire _2688__bF$buf1 ;
wire _2688__bF$buf2 ;
wire _2688__bF$buf3 ;
wire _6294_ ;
wire _4607_ ;
wire [31:0] \datapath._03_  ;
wire _7499_ ;
wire _7079_ ;
wire _8860_ ;
wire _8440_ ;
wire _8020_ ;
wire \datapath.alu.b_4_bF$buf0  ;
wire _9225_ ;
wire _4780_ ;
wire _4360_ ;
wire _5985_ ;
wire _5565_ ;
wire _5145_ ;
wire _1485_ ;
wire _1065_ ;
wire _7711_ ;
wire _396_ ;
wire _8916_ ;
wire _3631_ ;
wire _3211_ ;
wire _4836_ ;
wire _4416_ ;
wire _9034_ ;
wire \datapath.alu.b_2_bF$buf7  ;
wire _2902_ ;
wire _5794_ ;
wire _5374_ ;
wire _6999_ ;
wire _6579_ ;
wire _6159_ ;
wire _1294_ ;
wire _7940_ ;
wire _7520_ ;
wire _7100_ ;
wire _2499_ ;
wire _2079_ ;
wire _8725_ ;
wire _8305_ ;
wire _3860_ ;
wire _3440_ ;
wire _3020_ ;
wire _4645_ ;
wire _4225_ ;
wire CLK_bF$buf40 ;
wire CLK_bF$buf41 ;
wire CLK_bF$buf42 ;
wire CLK_bF$buf43 ;
wire CLK_bF$buf44 ;
wire CLK_bF$buf45 ;
wire CLK_bF$buf46 ;
wire CLK_bF$buf47 ;
wire CLK_bF$buf48 ;
wire CLK_bF$buf49 ;
wire _9263_ ;
wire _2711_ ;
wire _5183_ ;
wire _3916_ ;
wire _6388_ ;
wire _8954_ ;
wire _8534_ ;
wire _8114_ ;
wire _9319_ ;
wire _4874_ ;
wire _4454_ ;
wire _4034_ ;
wire _5659_ ;
wire _5239_ ;
wire _6600_ ;
wire _9072_ ;
wire _1999_ ;
wire _1579_ ;
wire _1159_ ;
wire _7805_ ;
wire _2940_ ;
wire _2520_ ;
wire _2100_ ;
wire _3725_ ;
wire _3305_ ;
wire _6197_ ;
wire _8763_ ;
wire _8343_ ;
wire _9128_ ;
wire _4683_ ;
wire _4263_ ;
wire _702_ ;
wire _5888_ ;
wire _5468_ ;
wire _5048_ ;
wire _1388_ ;
wire _7614_ ;
wire [31:0] \datapath.registers.1226[0]  ;
wire _299_ ;
wire \datapath.idinstr_20_hier0_bF$buf6  ;
wire _8819_ ;
wire _3954_ ;
wire _3534_ ;
wire _3114_ ;
wire _4739_ ;
wire _4319_ ;
wire _8992_ ;
wire _8572_ ;
wire _8152_ ;
wire _6147__bF$buf0 ;
wire _6147__bF$buf1 ;
wire _6147__bF$buf2 ;
wire _6147__bF$buf3 ;
wire _6147__bF$buf4 ;
wire _18_ ;
wire _1600_ ;
wire _9357_ ;
wire _4492_ ;
wire _4072_ ;
wire \datapath.idinstr_20_bF$buf11  ;
wire _931_ ;
wire _511_ ;
wire _2805_ ;
wire _5697_ ;
wire _5277_ ;
wire _1197_ ;
wire _7843_ ;
wire _7423_ ;
wire _7003_ ;
wire _8628_ ;
wire _8208_ ;
wire _3763_ ;
wire _3343_ ;
wire _4968_ ;
wire _4548_ ;
wire \datapath.idinstr_21_bF$buf20  ;
wire _4128_ ;
wire _8381_ ;
wire _9166_ ;
wire _740_ ;
wire _320_ ;
wire _2614_ ;
wire _5086_ ;
wire \datapath.idinstr_15_bF$buf25  ;
wire _3819_ ;
wire _7652_ ;
wire _7232_ ;
wire _8857_ ;
wire _8437_ ;
wire _8017_ ;
wire _3992_ ;
wire _3572_ ;
wire _3152_ ;
wire _4777_ ;
wire _4357_ ;
wire _8190_ ;
wire \datapath.idinstr_16_bF$buf34  ;
wire _56_ ;
wire _6923_ ;
wire _6503_ ;
wire _9395_ ;
wire _7708_ ;
wire _2843_ ;
wire _2423_ ;
wire _2003_ ;
wire _3628_ ;
wire _3208_ ;
wire _7881_ ;
wire _7461_ ;
wire _7041_ ;
wire _8666_ ;
wire _8246_ ;
wire _3381_ ;
wire _4586_ ;
wire _4166_ ;
wire _605_ ;
wire _6732_ ;
wire _6312_ ;
wire _7937_ ;
wire _7517_ ;
wire _2652_ ;
wire _2232_ ;
wire _3857_ ;
wire _3437_ ;
wire _3017_ ;
wire _7690_ ;
wire _7270_ ;
wire _8895_ ;
wire _8475_ ;
wire _8055_ ;
wire _3190_ ;
wire _1923_ ;
wire _1503_ ;
wire _4395_ ;
wire _834_ ;
wire _414_ ;
wire _2708_ ;
wire _94_ ;
wire _6961_ ;
wire _6541_ ;
wire _6121_ ;
wire _7607__bF$buf0 ;
wire _7607__bF$buf1 ;
wire _7607__bF$buf2 ;
wire _7607__bF$buf3 ;
wire _7607__bF$buf4 ;
wire _7746_ ;
wire _7326_ ;
wire _2881_ ;
wire _2461_ ;
wire _2041_ ;
wire [31:0] \datapath.registers.1226[16]  ;
wire _3666_ ;
wire _3246_ ;
wire _5812_ ;
wire _8284_ ;
wire _1732_ ;
wire _1312_ ;
wire _9069_ ;
wire _643_ ;
wire _223_ ;
wire _2937_ ;
wire _2517_ ;
wire _7611__bF$buf0 ;
wire _7611__bF$buf1 ;
wire _7611__bF$buf2 ;
wire _6770_ ;
wire _7611__bF$buf3 ;
wire _6350_ ;
wire _7611__bF$buf4 ;
wire _7611__bF$buf5 ;
wire _7611__bF$buf6 ;
wire _7611__bF$buf7 ;
wire _7611__bF$buf8 ;
wire _7611__bF$buf9 ;
wire _7975_ ;
wire _7555_ ;
wire _7135_ ;
wire _2690_ ;
wire _2270_ ;
wire _3895_ ;
wire _3475_ ;
wire _3055_ ;
wire [31:0] \datapath.memdataload  ;
wire _5621_ ;
wire _5201_ ;
wire _8093_ ;
wire _6826_ ;
wire _6406_ ;
wire _1961_ ;
wire _1541_ ;
wire _1121_ ;
wire _9298_ ;
wire _872_ ;
wire _452_ ;
wire _2746_ ;
wire _2326_ ;
wire _7784_ ;
wire _7364_ ;
wire _8989_ ;
wire _8569_ ;
wire _8149_ ;
wire _3284_ ;
wire _4489_ ;
wire _4069_ ;
wire _5850_ ;
wire _5430_ ;
wire _5010_ ;
wire _928_ ;
wire _508_ ;
wire _6635_ ;
wire _6215_ ;
wire _1770_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _2975_ ;
wire _2555_ ;
wire _2135_ ;
wire _4701_ ;
wire _7593_ ;
wire _7173_ ;
wire \datapath.idinstr_21_bF$buf17  ;
wire _5906_ ;
wire _8798_ ;
wire _8378_ ;
wire _3093_ ;
wire _1826_ ;
wire _1406_ ;
wire _4298_ ;
wire _737_ ;
wire _317_ ;
wire \datapath.idinstr_17_bF$buf2  ;
wire _6864_ ;
wire _6444_ ;
wire _6024_ ;
wire \datapath._60_  ;
wire _490_ ;
wire \datapath.idinstr_22_bF$buf26  ;
wire _7649_ ;
wire _7229_ ;
wire _2784_ ;
wire _2364_ ;
wire _3989_ ;
wire _3569_ ;
wire _3149_ ;
wire _4930_ ;
wire _4510_ ;
wire _5715_ ;
wire _2680__bF$buf0 ;
wire _2680__bF$buf1 ;
wire _2680__bF$buf2 ;
wire _2680__bF$buf3 ;
wire _8187_ ;
wire _1635_ ;
wire _1215_ ;
wire \datapath.idinstr_21_bF$buf2  ;
wire \datapath.idinstr_20_bF$buf46  ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire \datapath.idinstr_15_bF$buf9  ;
wire _6673_ ;
wire _6253_ ;
wire _7878_ ;
wire _7458_ ;
wire _7038_ ;
wire _2593_ ;
wire _2173_ ;
wire _3798_ ;
wire _3378_ ;
wire _5944_ ;
wire _5524_ ;
wire _5104_ ;
wire _6729_ ;
wire _6309_ ;
wire _1864_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire [31:0] \datapath.registers.regb_data  ;
wire _2649_ ;
wire _2229_ ;
wire _6482_ ;
wire _6062_ ;
wire _7687_ ;
wire _7267_ ;
wire _3187_ ;
wire _9413_ ;
wire _5753_ ;
wire _5333_ ;
wire _6958_ ;
wire _6538_ ;
wire _6118_ ;
wire _1673_ ;
wire _1253_ ;
wire _584_ ;
wire _164_ ;
wire _2878_ ;
wire _2458_ ;
wire _2038_ ;
wire _6291_ ;
wire _4604_ ;
wire _7496_ ;
wire _7076_ ;
wire _5759__bF$buf0 ;
wire _5759__bF$buf1 ;
wire _5759__bF$buf2 ;
wire _5759__bF$buf3 ;
wire _5759__bF$buf4 ;
wire _5809_ ;
wire _9222_ ;
wire _1729_ ;
wire _1309_ ;
wire _5982_ ;
wire _5562_ ;
wire _5142_ ;
wire _6767_ ;
wire _6347_ ;
wire _1482_ ;
wire _1062_ ;
wire _393_ ;
wire \datapath.idinstr_24_bF$buf5  ;
wire _2687_ ;
wire _2267_ ;
wire _8913_ ;
wire _617__bF$buf0 ;
wire _617__bF$buf1 ;
wire _617__bF$buf2 ;
wire _617__bF$buf3 ;
wire _617__bF$buf4 ;
wire _4833_ ;
wire _4413_ ;
wire _5618_ ;
wire _9031_ ;
wire \datapath.alu.b_2_bF$buf4  ;
wire _1958_ ;
wire _1538_ ;
wire _1118_ ;
wire _5791_ ;
wire _5371_ ;
wire _869_ ;
wire _449_ ;
wire _6996_ ;
wire _6576_ ;
wire _6156_ ;
wire _1291_ ;
wire _2496_ ;
wire _2076_ ;
wire _8722_ ;
wire _8302_ ;
wire _4642_ ;
wire _4222_ ;
wire CLK_bF$buf10 ;
wire CLK_bF$buf11 ;
wire CLK_bF$buf12 ;
wire CLK_bF$buf13 ;
wire CLK_bF$buf14 ;
wire CLK_bF$buf15 ;
wire CLK_bF$buf16 ;
wire CLK_bF$buf17 ;
wire CLK_bF$buf18 ;
wire CLK_bF$buf19 ;
wire _5847_ ;
wire _5427_ ;
wire _5007_ ;
wire _9260_ ;
wire _1767_ ;
wire _1347_ ;
wire _5180_ ;
wire _678_ ;
wire _258_ ;
wire _3913_ ;
wire _6385_ ;
wire _5546__bF$buf0 ;
wire _5546__bF$buf1 ;
wire _5546__bF$buf2 ;
wire _5546__bF$buf3 ;
wire _5546__bF$buf4 ;
wire _5546__bF$buf5 ;
wire _8951_ ;
wire _5546__bF$buf6 ;
wire _8531_ ;
wire _5546__bF$buf7 ;
wire _8111_ ;
wire _5546__bF$buf8 ;
wire _5546__bF$buf9 ;
wire _9316_ ;
wire _4871_ ;
wire _4451_ ;
wire _4031_ ;
wire _5656_ ;
wire _5236_ ;
wire _1996_ ;
wire _1576_ ;
wire _1156_ ;
wire _7802_ ;
wire _487_ ;
wire [31:0] DMEM_DATA_L ;
wire _3722_ ;
wire _3302_ ;
wire [31:0] DMEM_DATA_S ;
wire _6194_ ;
wire _4927_ ;
wire _4507_ ;
wire _7399_ ;
wire _8760_ ;
wire _8340_ ;
wire _9125_ ;
wire _4680_ ;
wire _4260_ ;
wire _5885_ ;
wire _5465_ ;
wire _5045_ ;
wire _1385_ ;
wire _7611_ ;
wire _296_ ;
wire \datapath.idinstr_20_hier0_bF$buf3  ;
wire _8816_ ;
wire _3951_ ;
wire _3531_ ;
wire _3111_ ;
wire _4736_ ;
wire _4316_ ;
wire _15_ ;
wire _9354_ ;
wire _2802_ ;
wire _5694_ ;
wire _5274_ ;
wire _6899_ ;
wire _6479_ ;
wire _6059_ ;
wire _1194_ ;
wire _7840_ ;
wire _7420_ ;
wire _7000_ ;
wire _2399_ ;
wire _8625_ ;
wire _8205_ ;
wire _3760_ ;
wire _3340_ ;
wire _4965_ ;
wire _4545_ ;
wire _4125_ ;
wire _9163_ ;
wire _2611_ ;
wire _5083_ ;
wire [31:0] \datapath.registers.1226[31]  ;
wire \datapath.idinstr_15_bF$buf22  ;
wire _3816_ ;
wire _6288_ ;
wire _8854_ ;
wire _8434_ ;
wire _8014_ ;
wire _9219_ ;
wire _4774_ ;
wire _4354_ ;
wire [31:0] \datapath.abypass  ;
wire _5979_ ;
wire _5559_ ;
wire _5139_ ;
wire \datapath.idinstr_16_bF$buf31  ;
wire _53_ ;
wire _6920_ ;
wire _6500_ ;
wire _9392_ ;
wire _1899_ ;
wire _1479_ ;
wire _1059_ ;
wire _7705_ ;
wire _2840_ ;
wire _2420_ ;
wire _2000_ ;
wire _3625_ ;
wire _3205_ ;
wire _6097_ ;
wire _8663_ ;
wire _8243_ ;
wire \datapath.idinstr_17_bF$buf40  ;
wire _9028_ ;
wire _4583_ ;
wire _4163_ ;
wire _602_ ;
wire _5788_ ;
wire _5368_ ;
wire _1288_ ;
wire _7934_ ;
wire _7514_ ;
wire _199_ ;
wire _8719_ ;
wire _3854_ ;
wire _3434_ ;
wire _3014_ ;
wire _4639_ ;
wire _4219_ ;
wire _8892_ ;
wire _8472_ ;
wire _8052_ ;
wire [31:0] \datapath.regcsrmem  ;
wire _1920_ ;
wire _1500_ ;
wire _9257_ ;
wire _4392_ ;
wire _831_ ;
wire _411_ ;
wire _2705_ ;
wire _5597_ ;
wire _5177_ ;
wire _91_ ;
wire _1097_ ;
wire _7743_ ;
wire _7323_ ;
wire _494__bF$buf0 ;
wire _494__bF$buf1 ;
wire _494__bF$buf2 ;
wire _8948_ ;
wire _494__bF$buf3 ;
wire _8528_ ;
wire _494__bF$buf4 ;
wire _8108_ ;
wire _3663_ ;
wire _3243_ ;
wire _4868_ ;
wire _4448_ ;
wire _4028_ ;
wire _8281_ ;
wire _9066_ ;
wire _640_ ;
wire _220_ ;
wire _2934_ ;
wire _2514_ ;
wire _3719_ ;
wire _7972_ ;
wire _7552_ ;
wire _7132_ ;
wire _8757_ ;
wire _8337_ ;
wire _3892_ ;
wire _3472_ ;
wire _3052_ ;
wire _4677_ ;
wire _4257_ ;
wire _8090_ ;
wire _6823_ ;
wire _6403_ ;
wire _9295_ ;
wire _3796__bF$buf0 ;
wire _3796__bF$buf1 ;
wire _3796__bF$buf2 ;
wire _3796__bF$buf3 ;
wire _3796__bF$buf4 ;
wire CLK_hier0_bF$buf10 ;
wire CLK_hier0_bF$buf11 ;
wire _7608_ ;
wire _2743_ ;
wire _2323_ ;
wire _3948_ ;
wire _3528_ ;
wire _3108_ ;
wire _9_ ;
wire _7781_ ;
wire _7361_ ;
wire _8986_ ;
wire _8566_ ;
wire _8146_ ;
wire _3281_ ;
wire _4486_ ;
wire _4066_ ;
wire _925_ ;
wire _505_ ;
wire _6632_ ;
wire _6212_ ;
wire _7837_ ;
wire _7417_ ;
wire _2972_ ;
wire _2552_ ;
wire _2132_ ;
wire _3757_ ;
wire _3337_ ;
wire _7590_ ;
wire _7170_ ;
wire \datapath.idinstr_21_bF$buf14  ;
wire _5903_ ;
wire _8795_ ;
wire _8375_ ;
wire _3090_ ;
wire \datapath.regmret_bF$buf3  ;
wire _1823_ ;
wire _1403_ ;
wire _4295_ ;
wire _734_ ;
wire _314_ ;
wire _2608_ ;
wire _6861_ ;
wire _6441_ ;
wire _6021_ ;
wire \datapath.idinstr_15_bF$buf19  ;
wire \datapath.idinstr_22_bF$buf23  ;
wire _7646_ ;
wire _7226_ ;
wire _2781_ ;
wire _2361_ ;
wire _3986_ ;
wire _3566_ ;
wire _7614__bF$buf0 ;
wire _3146_ ;
wire _7614__bF$buf1 ;
wire _7614__bF$buf2 ;
wire _7614__bF$buf3 ;
wire _7614__bF$buf4 ;
wire _5712_ ;
wire _8184_ ;
wire \datapath.idinstr_16_bF$buf28  ;
wire _6917_ ;
wire _1632_ ;
wire _1212_ ;
wire _9389_ ;
wire \datapath.idinstr_20_bF$buf43  ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _2837_ ;
wire \datapath.idinstr_15_bF$buf6  ;
wire _2417_ ;
wire _6670_ ;
wire _6250_ ;
wire _7875_ ;
wire _7455_ ;
wire _7035_ ;
wire _2590_ ;
wire _2170_ ;
wire _3795_ ;
wire _3375_ ;
wire \datapath.idinstr_17_bF$buf37  ;
wire _5941_ ;
wire _5521_ ;
wire _5101_ ;
wire _6726_ ;
wire _6306_ ;
wire _1861_ ;
wire _1441_ ;
wire _1021_ ;
wire _9198_ ;
wire _772_ ;
wire _352_ ;
wire _2646_ ;
wire _2226_ ;
wire _7684_ ;
wire _7264_ ;
wire [31:0] \datapath.registers.1226[7]  ;
wire _8889_ ;
wire _8469_ ;
wire _8049_ ;
wire _3184_ ;
wire _9410_ ;
wire _1917_ ;
wire _4389_ ;
wire _5750_ ;
wire _5330_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _6955_ ;
wire _6535_ ;
wire _6115_ ;
wire _1670_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _2875_ ;
wire _2455_ ;
wire _2035_ ;
wire _4601_ ;
wire _7493_ ;
wire _7073_ ;
wire _5806_ ;
wire _8698_ ;
wire _8278_ ;
wire _1726_ ;
wire _1306_ ;
wire _4198_ ;
wire _637_ ;
wire _217_ ;
wire _5486__bF$buf0 ;
wire _5486__bF$buf1 ;
wire _5486__bF$buf2 ;
wire _5486__bF$buf3 ;
wire _6764_ ;
wire _5486__bF$buf4 ;
wire _6344_ ;
wire \datapath._50_  ;
wire _390_ ;
wire _7969_ ;
wire _7549_ ;
wire _7129_ ;
wire \datapath.idinstr_24_bF$buf2  ;
wire _2684_ ;
wire _2264_ ;
wire _8910_ ;
wire _3889_ ;
wire _3469_ ;
wire _3049_ ;
wire _4830_ ;
wire _4410_ ;
wire _5615_ ;
wire _8087_ ;
wire \datapath.alu.b_2_bF$buf1  ;
wire _1955_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire _5490__bF$buf0 ;
wire _5490__bF$buf1 ;
wire _5490__bF$buf2 ;
wire _5490__bF$buf3 ;
wire _5490__bF$buf4 ;
wire \datapath.tkbranch  ;
wire _6993_ ;
wire _6573_ ;
wire _6153_ ;
wire _7778_ ;
wire _7358_ ;
wire _2493_ ;
wire _2073_ ;
wire \datapath.idinstr_22_bF$buf9  ;
wire _3698_ ;
wire _3278_ ;
wire _5844_ ;
wire _5424_ ;
wire _5004_ ;
wire _6629_ ;
wire _6209_ ;
wire _1764_ ;
wire _1344_ ;
wire _675_ ;
wire _255_ ;
wire _2969_ ;
wire _2549_ ;
wire _2129_ ;
wire _3910_ ;
wire _6382_ ;
wire _7587_ ;
wire _7167_ ;
wire _3087_ ;
wire _9313_ ;
wire _5653_ ;
wire _5233_ ;
wire _6858_ ;
wire _6438_ ;
wire _6018_ ;
wire _1993_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _2778_ ;
wire _2358_ ;
wire _6191_ ;
wire _4924_ ;
wire _4504_ ;
wire _7396_ ;
wire _5709_ ;
wire _9122_ ;
wire _1629_ ;
wire _1209_ ;
wire _5882_ ;
wire _5462_ ;
wire _5042_ ;
wire \bypassandflushunit.flushid  ;
wire _6667_ ;
wire _6247_ ;
wire _1382_ ;
wire _293_ ;
wire _2587_ ;
wire _2167_ ;
wire \datapath.idinstr_20_hier0_bF$buf0  ;
wire _8813_ ;
wire _4733_ ;
wire _4313_ ;
wire _5938_ ;
wire _5518_ ;
wire _12_ ;
wire _9351_ ;
wire _1858_ ;
wire _1438_ ;
wire _1018_ ;
wire _5691_ ;
wire _5271_ ;
wire _769_ ;
wire _349_ ;
wire _6896_ ;
wire _6476_ ;
wire _6056_ ;
wire _1191_ ;
wire _2396_ ;
wire _8622_ ;
wire _8202_ ;
wire _9407_ ;
wire _4962_ ;
wire _4542_ ;
wire _4122_ ;
wire _5747_ ;
wire _5327_ ;
wire _9160_ ;
wire _1667_ ;
wire _1247_ ;
wire _5080_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _3813_ ;
wire _6285_ ;
wire _8851_ ;
wire _8431_ ;
wire _8011_ ;
wire _9216_ ;
wire _4771_ ;
wire _4351_ ;
wire \datapath.idinstr_21_hier0_bF$buf5  ;
wire _5976_ ;
wire _5556_ ;
wire _5136_ ;
wire _50_ ;
wire _1896_ ;
wire _1476_ ;
wire _1056_ ;
wire _7702_ ;
wire _387_ ;
wire _8907_ ;
wire _3622_ ;
wire _3202_ ;
wire _6094_ ;
wire _4827_ ;
wire _4407_ ;
wire _7299_ ;
wire _8660_ ;
wire _8240_ ;
wire _9025_ ;
wire _4580_ ;
wire _4160_ ;
wire _5785_ ;
wire _5365_ ;
wire _1285_ ;
wire _7931_ ;
wire _7511_ ;
wire _196_ ;
wire _8716_ ;
wire _3851_ ;
wire _3431_ ;
wire _3011_ ;
wire _4636_ ;
wire _4216_ ;
wire _9254_ ;
wire _2702_ ;
wire _5594_ ;
wire _5174_ ;
wire _3907_ ;
wire _6799_ ;
wire _6379_ ;
wire _1094_ ;
wire _7740_ ;
wire _7320_ ;
wire _2299_ ;
wire _8945_ ;
wire _8525_ ;
wire _8105_ ;
wire _3660_ ;
wire _3240_ ;
wire _4865_ ;
wire _4445_ ;
wire _4025_ ;
wire _5434__bF$buf0 ;
wire _5434__bF$buf1 ;
wire _5434__bF$buf2 ;
wire _5434__bF$buf3 ;
wire _9063_ ;
wire _5434__bF$buf4 ;
wire _5434__bF$buf5 ;
wire _5434__bF$buf6 ;
wire _5434__bF$buf7 ;
wire _5434__bF$buf8 ;
wire _5434__bF$buf9 ;
wire _2931_ ;
wire _2511_ ;
wire [31:0] \datapath.registers.1226[21]  ;
wire _3716_ ;
wire _6188_ ;
wire _8754_ ;
wire _8334_ ;
wire _9119_ ;
wire _4674_ ;
wire _4254_ ;
wire _5927__bF$buf0 ;
wire _5927__bF$buf1 ;
wire _5927__bF$buf2 ;
wire _5927__bF$buf3 ;
wire _5927__bF$buf4 ;
wire _5879_ ;
wire _5459_ ;
wire _5039_ ;
wire _6820_ ;
wire _6400_ ;
wire _9292_ ;
wire _1799_ ;
wire _1379_ ;
wire _7605_ ;
wire _2740_ ;
wire _2320_ ;
wire _3945_ ;
wire _3525_ ;
wire _3105_ ;
wire _6_ ;
wire _8983_ ;
wire _8563_ ;
wire _8143_ ;
wire _9348_ ;
wire _4483_ ;
wire _4063_ ;
wire _922_ ;
wire _502_ ;
wire _5688_ ;
wire _5268_ ;
wire _1188_ ;
wire _7834_ ;
wire _7414_ ;
wire _8619_ ;
wire _3754_ ;
wire _3334_ ;
wire _4959_ ;
wire _4539_ ;
wire \datapath.idinstr_21_bF$buf11  ;
wire _4119_ ;
wire _5900_ ;
wire _8792_ ;
wire _8372_ ;
wire \datapath.regmret_bF$buf0  ;
wire _497__bF$buf0 ;
wire _497__bF$buf1 ;
wire _497__bF$buf2 ;
wire _497__bF$buf3 ;
wire _497__bF$buf4 ;
wire _1820_ ;
wire _1400_ ;
wire _9157_ ;
wire _4292_ ;
wire _731_ ;
wire _311_ ;
wire _2605_ ;
wire _5497_ ;
wire _5077_ ;
wire \datapath.idinstr_15_bF$buf16  ;
wire \datapath.idinstr_15_hier0_bF$buf4  ;
wire \datapath.idinstr_22_bF$buf20  ;
wire _7643_ ;
wire _7223_ ;
wire _8848_ ;
wire _8428_ ;
wire _8008_ ;
wire _3983_ ;
wire _3563_ ;
wire _3143_ ;
wire _4768_ ;
wire _4348_ ;
wire _8181_ ;
wire \datapath.idinstr_16_bF$buf25  ;
wire _47_ ;
wire _6914_ ;
wire _9386_ ;
wire _6141__bF$buf10 ;
wire \datapath.idinstr_20_bF$buf40  ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _2834_ ;
wire \datapath.idinstr_15_bF$buf3  ;
wire _2414_ ;
wire _3619_ ;
wire _7872_ ;
wire _7452_ ;
wire _7032_ ;
wire _8657_ ;
wire _8237_ ;
wire _3792_ ;
wire _3372_ ;
wire \datapath.idinstr_17_bF$buf34  ;
wire _4997_ ;
wire _4577_ ;
wire _4157_ ;
wire _6723_ ;
wire _6303_ ;
wire _9195_ ;
wire _7928_ ;
wire _7508_ ;
wire _2643_ ;
wire _2223_ ;
wire _5546__bF$buf10 ;
wire _5546__bF$buf11 ;
wire _5546__bF$buf12 ;
wire _5546__bF$buf13 ;
wire _5546__bF$buf14 ;
wire _5546__bF$buf15 ;
wire _3848_ ;
wire _3428_ ;
wire _3008_ ;
wire _7681_ ;
wire _7261_ ;
wire _8886_ ;
wire _8466_ ;
wire _8046_ ;
wire _3181_ ;
wire _1914_ ;
wire _4386_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _6952_ ;
wire _6532_ ;
wire _6112_ ;
wire _7737_ ;
wire _7317_ ;
wire _2872_ ;
wire _2452_ ;
wire _2032_ ;
wire _3657_ ;
wire _3237_ ;
wire _7490_ ;
wire _7070_ ;
wire _5803_ ;
wire _8695_ ;
wire _8275_ ;
wire _1723_ ;
wire _1303_ ;
wire _4195_ ;
wire _634_ ;
wire _214_ ;
wire _2928_ ;
wire _2508_ ;
wire _6761_ ;
wire _6341_ ;
wire _9244__bF$buf0 ;
wire _9244__bF$buf1 ;
wire _9244__bF$buf2 ;
wire _9244__bF$buf3 ;
wire _9244__bF$buf4 ;
wire _7966_ ;
wire _7546_ ;
wire _7126_ ;
wire _2681_ ;
wire _2261_ ;
wire \datapath.idinstr_18_bF$buf6  ;
wire _3886_ ;
wire _3466_ ;
wire _3046_ ;
wire _5612_ ;
wire _8084_ ;
wire \datapath.pcstall_bF$buf5  ;
wire _6817_ ;
wire _1952_ ;
wire _1532_ ;
wire _1112_ ;
wire _9289_ ;
wire _863_ ;
wire _443_ ;
wire _2737_ ;
wire _2317_ ;
wire _6990_ ;
wire _6570_ ;
wire _6150_ ;
wire _7775_ ;
wire _7355_ ;
wire _2490_ ;
wire _2070_ ;
wire \datapath.idinstr_22_bF$buf6  ;
wire _3695_ ;
wire _3275_ ;
wire _5841_ ;
wire _5421_ ;
wire _5001_ ;
wire _919_ ;
wire _6626_ ;
wire _6206_ ;
wire _1761_ ;
wire _1341_ ;
wire _9098_ ;
wire _672_ ;
wire _252_ ;
wire _2966_ ;
wire _2546_ ;
wire _2126_ ;
wire _7584_ ;
wire _7164_ ;
wire _8789_ ;
wire _8369_ ;
wire _3084_ ;
wire _9310_ ;
wire _1817_ ;
wire _4289_ ;
wire _5650_ ;
wire _5230_ ;
wire _728_ ;
wire _308_ ;
wire [1:0] \controlunit.pc_sel  ;
wire _6855_ ;
wire _6435_ ;
wire _6015_ ;
wire _1990_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire \datapath.idinstr_22_bF$buf17  ;
wire _2775_ ;
wire _2355_ ;
wire _4921_ ;
wire _4501_ ;
wire _7393_ ;
wire _5706_ ;
wire _8598_ ;
wire _8178_ ;
wire _1626_ ;
wire _1206_ ;
wire _4098_ ;
wire \datapath.idinstr_20_bF$buf37  ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire _6664_ ;
wire _6244_ ;
wire _290_ ;
wire _7869_ ;
wire _7449_ ;
wire _7029_ ;
wire _2584_ ;
wire _2164_ ;
wire _8810_ ;
wire _3789_ ;
wire _3369_ ;
wire _4730_ ;
wire _4310_ ;
wire _5935_ ;
wire _5515_ ;
wire \datapath.alu.b_0_bF$buf7  ;
wire _1855_ ;
wire _1435_ ;
wire _1015_ ;
wire _766_ ;
wire _346_ ;
wire _6893_ ;
wire _6473_ ;
wire _6053_ ;
wire _7678_ ;
wire _7258_ ;
wire _2393_ ;
wire _3598_ ;
wire _3178_ ;
wire _9404_ ;
wire _5744_ ;
wire _5324_ ;
wire [29:0] \datapath.csr._26_  ;
wire _6949_ ;
wire _6529_ ;
wire _6109_ ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire _2869_ ;
wire _2449_ ;
wire _2029_ ;
wire _3810_ ;
wire _6282_ ;
wire _7487_ ;
wire _7067_ ;
wire _9213_ ;
wire \datapath.idinstr_21_hier0_bF$buf2  ;
wire _5973_ ;
wire _5553_ ;
wire _5133_ ;
wire _6758_ ;
wire _6338_ ;
wire _1893_ ;
wire _1473_ ;
wire _1053_ ;
wire _384_ ;
wire _2678_ ;
wire _2258_ ;
wire _8904_ ;
wire _6091_ ;
wire _4824_ ;
wire _4404_ ;
wire _7296_ ;
wire _5609_ ;
wire _9442_ ;
wire _9022_ ;
wire _1949_ ;
wire _1529_ ;
wire _1109_ ;
wire _5782_ ;
wire _5362_ ;
wire [1:0] \controlunit.wb_sel  ;
wire _6987_ ;
wire _6567_ ;
wire _6147_ ;
wire _1282_ ;
wire _193_ ;
wire _2487_ ;
wire _2067_ ;
wire _8713_ ;
wire _4633_ ;
wire _4213_ ;
wire _5838_ ;
wire _5418_ ;
wire _9251_ ;
wire _1758_ ;
wire _1338_ ;
wire _5591_ ;
wire _5171_ ;
wire _669_ ;
wire [31:0] _249_ ;
wire _3904_ ;
wire _6796_ ;
wire _6376_ ;
wire _1091_ ;
wire _2296_ ;
wire _8942_ ;
wire _8522_ ;
wire _8102_ ;
wire [31:0] \datapath.alupc  ;
wire _9307_ ;
wire _4862_ ;
wire _4442_ ;
wire _4022_ ;
wire _5647_ ;
wire _5227_ ;
wire _9060_ ;
wire _1987_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _3713_ ;
wire _6185_ ;
wire _4918_ ;
wire _8751_ ;
wire _8331_ ;
wire _9116_ ;
wire _4671_ ;
wire _4251_ ;
wire _5876_ ;
wire _5456_ ;
wire _5036_ ;
wire _1796_ ;
wire _1376_ ;
wire _7602_ ;
wire _287_ ;
wire _8807_ ;
wire _3942_ ;
wire _3522_ ;
wire _3102_ ;
wire _3_ ;
wire _4727_ ;
wire _4307_ ;
wire _7199_ ;
wire _8980_ ;
wire _8560_ ;
wire _8140_ ;
wire _9345_ ;
wire _4480_ ;
wire _4060_ ;
wire _5685_ ;
wire _5265_ ;
wire _1185_ ;
wire _7831_ ;
wire _7411_ ;
wire _8616_ ;
wire _3751_ ;
wire _3331_ ;
wire _4956_ ;
wire _4536_ ;
wire _4116_ ;
wire _9154_ ;
wire _2602_ ;
wire _5494_ ;
wire _5074_ ;
wire CLK_bF$buf130 ;
wire CLK_bF$buf131 ;
wire CLK_bF$buf132 ;
wire CLK_bF$buf133 ;
wire CLK_bF$buf134 ;
wire CLK_bF$buf135 ;
wire \datapath.idinstr_15_bF$buf13  ;
wire CLK_bF$buf136 ;
wire CLK_bF$buf137 ;
wire CLK_bF$buf138 ;
wire _3807_ ;
wire CLK_bF$buf139 ;
wire \datapath.idinstr_15_hier0_bF$buf1  ;
wire _6699_ ;
wire _6279_ ;
wire _7640_ ;
wire _7220_ ;
wire _2199_ ;
wire _8845_ ;
wire _8425_ ;
wire _8005_ ;
wire _3980_ ;
wire _3560_ ;
wire _3140_ ;
wire _4765_ ;
wire _4345_ ;
wire \datapath.idinstr_16_bF$buf22  ;
wire _44_ ;
wire _6911_ ;
wire _9383_ ;
wire _2831_ ;
wire \datapath.idinstr_15_bF$buf0  ;
wire _2411_ ;
wire [31:0] \datapath.registers.1226[11]  ;
wire _3616_ ;
wire _6088_ ;
wire _8654_ ;
wire _8234_ ;
wire \datapath.idinstr_17_bF$buf31  ;
wire _9439_ ;
wire _9019_ ;
wire _4994_ ;
wire _4574_ ;
wire _4154_ ;
wire _5779_ ;
wire _5359_ ;
wire _6720_ ;
wire _6300_ ;
wire _9192_ ;
wire _1699_ ;
wire _1279_ ;
wire _7925_ ;
wire _7505_ ;
wire _2640_ ;
wire _2220_ ;
wire \datapath.idinstr_15_bF$buf51  ;
wire _3845_ ;
wire _3425_ ;
wire _3005_ ;
wire _8883_ ;
wire _8463_ ;
wire _8043_ ;
wire _9109__bF$buf0 ;
wire _9109__bF$buf1 ;
wire _9109__bF$buf2 ;
wire _9109__bF$buf3 ;
wire _9109__bF$buf4 ;
wire _1911_ ;
wire _9248_ ;
wire _4383_ ;
wire _822_ ;
wire _402_ ;
wire _5588_ ;
wire _5168_ ;
wire _82_ ;
wire _1088_ ;
wire _7734_ ;
wire _7314_ ;
wire _8939_ ;
wire _8519_ ;
wire _3654_ ;
wire _3234_ ;
wire _4859_ ;
wire _4439_ ;
wire _4019_ ;
wire _5800_ ;
wire _8692_ ;
wire _8272_ ;
wire _1720_ ;
wire _1300_ ;
wire _9057_ ;
wire _4192_ ;
wire _631_ ;
wire _211_ ;
wire _2925_ ;
wire _2505_ ;
wire _5397_ ;
wire _7963_ ;
wire _7543_ ;
wire _7123_ ;
wire \datapath.idinstr_18_bF$buf3  ;
wire _8748_ ;
wire _8328_ ;
wire _3883_ ;
wire _3463_ ;
wire _3043_ ;
wire _0__1_bF$buf0 ;
wire _0__1_bF$buf1 ;
wire _0__1_bF$buf2 ;
wire _0__1_bF$buf3 ;
wire _0__1_bF$buf4 ;
wire _0__1_bF$buf5 ;
wire _0__1_bF$buf6 ;
wire _0__1_bF$buf7 ;
wire _4668_ ;
wire _0__1_bF$buf8 ;
wire _4248_ ;
wire _0__1_bF$buf9 ;
wire _8081_ ;
wire \datapath.pcstall_bF$buf2  ;
wire _6814_ ;
wire _9286_ ;
wire _860_ ;
wire _440_ ;
wire _2734_ ;
wire _2314_ ;
wire _3939_ ;
wire _3519_ ;
wire _7772_ ;
wire _7352_ ;
wire \datapath.idinstr_22_bF$buf3  ;
wire _8977_ ;
wire _8557_ ;
wire _8137_ ;
wire _3692_ ;
wire _3272_ ;
wire _4897_ ;
wire _4477_ ;
wire _4057_ ;
wire _916_ ;
wire _6623_ ;
wire _6203_ ;
wire _9095_ ;
wire _7828_ ;
wire _7408_ ;
wire _2963_ ;
wire _2543_ ;
wire _2123_ ;
wire _3748_ ;
wire _3328_ ;
wire _7581_ ;
wire _7161_ ;
wire _8786_ ;
wire _8366_ ;
wire _3081_ ;
wire _1814_ ;
wire _4286_ ;
wire _725_ ;
wire _305_ ;
wire _6852_ ;
wire _6432_ ;
wire _6012_ ;
wire \datapath.idinstr_22_bF$buf14  ;
wire _7637_ ;
wire _7217_ ;
wire _2772_ ;
wire _2352_ ;
wire _3977_ ;
wire _3557_ ;
wire _3137_ ;
wire _7390_ ;
wire _5703_ ;
wire _8595_ ;
wire _8175_ ;
wire \datapath.idinstr_16_bF$buf19  ;
wire _6908_ ;
wire _1623_ ;
wire _1203_ ;
wire _4095_ ;
wire \datapath.idinstr_20_bF$buf34  ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _2828_ ;
wire _2408_ ;
wire _6661_ ;
wire _6241_ ;
wire _7866_ ;
wire _7446_ ;
wire _7026_ ;
wire _2581_ ;
wire _2161_ ;
wire [31:0] \datapath.registers.1226[28]  ;
wire _3786_ ;
wire _3366_ ;
wire \datapath.idinstr_17_bF$buf28  ;
wire \datapath.idinstr_21_bF$buf43  ;
wire _5932_ ;
wire _5512_ ;
wire _6717_ ;
wire \datapath.alu.b_0_bF$buf4  ;
wire _1852_ ;
wire _1432_ ;
wire _1012_ ;
wire _9189_ ;
wire _763_ ;
wire _343_ ;
wire _2637_ ;
wire _2217_ ;
wire _6890_ ;
wire _6470_ ;
wire _6050_ ;
wire \datapath.idinstr_15_bF$buf48  ;
wire _7675_ ;
wire _7255_ ;
wire _2390_ ;
wire _3595_ ;
wire _3175_ ;
wire _9401_ ;
wire _1908_ ;
wire _5741_ ;
wire _5321_ ;
wire _819_ ;
wire _79_ ;
wire _6946_ ;
wire _6526_ ;
wire _6106_ ;
wire _1661_ ;
wire _1241_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _2866_ ;
wire _2446_ ;
wire _2026_ ;
wire _7484_ ;
wire _7064_ ;
wire _8689_ ;
wire _8269_ ;
wire _9210_ ;
wire _1717_ ;
wire _4189_ ;
wire _5970_ ;
wire _5550_ ;
wire _5130_ ;
wire _628_ ;
wire _208_ ;
wire _6755_ ;
wire _6335_ ;
wire _1890_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _2675_ ;
wire _2255_ ;
wire _8901_ ;
wire _4821_ ;
wire _4401_ ;
wire _7293_ ;
wire _5606_ ;
wire _8498_ ;
wire _8078_ ;
wire _5496__bF$buf0 ;
wire _5496__bF$buf1 ;
wire _5496__bF$buf2 ;
wire _5496__bF$buf3 ;
wire _5496__bF$buf4 ;
wire _1946_ ;
wire _1526_ ;
wire _1106_ ;
wire _857_ ;
wire _437_ ;
wire _6984_ ;
wire _6564_ ;
wire _6144_ ;
wire [31:0] \datapath._30_  ;
wire _190_ ;
wire _7769_ ;
wire _7349_ ;
wire _2484_ ;
wire _2064_ ;
wire _8710_ ;
wire _3689_ ;
wire _3269_ ;
wire _4630_ ;
wire _4210_ ;
wire _5835_ ;
wire _5415_ ;
wire _1755_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire _3901_ ;
wire _6793_ ;
wire _6373_ ;
wire _7998_ ;
wire _7578_ ;
wire _7158_ ;
wire _2293_ ;
wire _3498_ ;
wire _3078_ ;
wire _9304_ ;
wire _5644_ ;
wire _5224_ ;
wire _6849_ ;
wire _6429_ ;
wire _6009_ ;
wire _1984_ ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _2769_ ;
wire _2349_ ;
wire _3710_ ;
wire _3802__bF$buf0 ;
wire _3802__bF$buf1 ;
wire _6182_ ;
wire _3802__bF$buf2 ;
wire _3802__bF$buf3 ;
wire _3802__bF$buf4 ;
wire _3802__bF$buf5 ;
wire _3802__bF$buf6 ;
wire _4915_ ;
wire _7387_ ;
wire [31:0] \datapath.jumptarget  ;
wire _2480__bF$buf0 ;
wire _2480__bF$buf1 ;
wire _2480__bF$buf2 ;
wire _2480__bF$buf3 ;
wire _2480__bF$buf4 ;
wire _2480__bF$buf5 ;
wire _9113_ ;
wire _5873_ ;
wire _5453_ ;
wire _5033_ ;
wire _6658_ ;
wire [2:0] abpsel ;
wire _6238_ ;
wire _1793_ ;
wire _1373_ ;
wire _284_ ;
wire _2998_ ;
wire _2578_ ;
wire _2158_ ;
wire _8804_ ;
wire [31:0] _0_ ;
wire _4724_ ;
wire _4304_ ;
wire _7196_ ;
wire _5929_ ;
wire _5509_ ;
wire _9342_ ;
wire _1849_ ;
wire _1429_ ;
wire _1009_ ;
wire _5682_ ;
wire _5262_ ;
wire _6887_ ;
wire _6467_ ;
wire _6047_ ;
wire _1182_ ;
wire _2387_ ;
wire _8613_ ;
wire _4953_ ;
wire _4533_ ;
wire _4113_ ;
wire _5738_ ;
wire _5318_ ;
wire _9151_ ;
wire _1658_ ;
wire _1238_ ;
wire _5491_ ;
wire _5071_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire CLK_bF$buf100 ;
wire CLK_bF$buf101 ;
wire CLK_bF$buf102 ;
wire CLK_bF$buf103 ;
wire CLK_bF$buf104 ;
wire CLK_bF$buf105 ;
wire \datapath.idinstr_15_bF$buf10  ;
wire CLK_bF$buf106 ;
wire _5510__bF$buf10 ;
wire CLK_bF$buf107 ;
wire _5510__bF$buf11 ;
wire CLK_bF$buf108 ;
wire _5510__bF$buf12 ;
wire _3804_ ;
wire CLK_bF$buf109 ;
wire _5510__bF$buf13 ;
wire _5510__bF$buf14 ;
wire _5510__bF$buf15 ;
wire _6696_ ;
wire _6276_ ;
wire _2196_ ;
wire _8842_ ;
wire _8422_ ;
wire _8002_ ;
wire _9207_ ;
wire _4762_ ;
wire _4342_ ;
wire _5967_ ;
wire _5547_ ;
wire _5127_ ;
wire _41_ ;
wire _9380_ ;
wire _1887_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _3613_ ;
wire _6085_ ;
wire _4818_ ;
wire _8651_ ;
wire _8231_ ;
wire _9436_ ;
wire _9016_ ;
wire _4991_ ;
wire _4571_ ;
wire _4151_ ;
wire _5776_ ;
wire _5356_ ;
wire _1696_ ;
wire _1276_ ;
wire _7922_ ;
wire _7502_ ;
wire _187_ ;
wire _8707_ ;
wire _3842_ ;
wire _3422_ ;
wire _3002_ ;
wire _4627_ ;
wire _4207_ ;
wire [31:0] \datapath._05_  ;
wire _7099_ ;
wire _8880_ ;
wire _8460_ ;
wire _8040_ ;
wire \datapath.idinstr_16_hier0_bF$buf3  ;
wire [31:0] \datapath.csr.csr_pcaddr  ;
wire _9245_ ;
wire _4380_ ;
wire _5585_ ;
wire _5165_ ;
wire _1085_ ;
wire _7731_ ;
wire _7311_ ;
wire _8936_ ;
wire _8516_ ;
wire _3651_ ;
wire _3231_ ;
wire _4856_ ;
wire _4436_ ;
wire _4016_ ;
wire _9054_ ;
wire _2922_ ;
wire _2502_ ;
wire _5394_ ;
wire _3707_ ;
wire _6599_ ;
wire _6179_ ;
wire _7960_ ;
wire _7540_ ;
wire _7120_ ;
wire \datapath.idinstr_18_bF$buf0  ;
wire _2099_ ;
wire _8745_ ;
wire _8325_ ;
wire _3880_ ;
wire _3460_ ;
wire _3040_ ;
wire _2495__bF$buf0 ;
wire _2495__bF$buf1 ;
wire _2495__bF$buf2 ;
wire _2495__bF$buf3 ;
wire _5444__bF$buf0 ;
wire _2495__bF$buf4 ;
wire _5444__bF$buf1 ;
wire _2495__bF$buf5 ;
wire _5444__bF$buf2 ;
wire _2495__bF$buf6 ;
wire _5444__bF$buf3 ;
wire _5444__bF$buf4 ;
wire _4665_ ;
wire _4245_ ;
wire _6811_ ;
wire _9283_ ;
wire _2731_ ;
wire _2311_ ;
wire _3675__bF$buf0 ;
wire _3675__bF$buf1 ;
wire _3675__bF$buf2 ;
wire _3675__bF$buf3 ;
wire _3675__bF$buf4 ;
wire _3936_ ;
wire _3516_ ;
wire \datapath.idinstr_22_bF$buf0  ;
wire \datapath.idinstr_16_bF$buf7  ;
wire _8974_ ;
wire _8554_ ;
wire _8134_ ;
wire _9339_ ;
wire _4894_ ;
wire _4474_ ;
wire _4054_ ;
wire _913_ ;
wire _5679_ ;
wire _5259_ ;
wire _6620_ ;
wire _6200_ ;
wire _9092_ ;
wire _1599_ ;
wire _1179_ ;
wire _7825_ ;
wire _7405_ ;
wire _2960_ ;
wire _2540_ ;
wire _2120_ ;
wire _3745_ ;
wire _3325_ ;
wire \datapath.idinstr_20_bF$buf7  ;
wire _8783_ ;
wire _8363_ ;
wire _1811_ ;
wire _9148_ ;
wire _4283_ ;
wire _722_ ;
wire _302_ ;
wire _5488_ ;
wire _5068_ ;
wire \datapath.idinstr_22_bF$buf11  ;
wire _7634_ ;
wire _7214_ ;
wire [31:0] \datapath.registers.1226[2]  ;
wire _8839_ ;
wire _8419_ ;
wire _3974_ ;
wire _3554_ ;
wire _3134_ ;
wire [31:0] \datapath.regrs2alu  ;
wire _4759_ ;
wire _4339_ ;
wire _5700_ ;
wire _8592_ ;
wire _8172_ ;
wire \datapath.idinstr_16_bF$buf16  ;
wire _38_ ;
wire _6905_ ;
wire _1620_ ;
wire _1200_ ;
wire _9377_ ;
wire _4092_ ;
wire \datapath.idinstr_20_bF$buf31  ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _2825_ ;
wire _2405_ ;
wire _5297_ ;
wire _7863_ ;
wire _7443_ ;
wire _7023_ ;
wire _8648_ ;
wire _8228_ ;
wire _3783_ ;
wire _3363_ ;
wire \datapath.idinstr_17_bF$buf25  ;
wire _4988_ ;
wire _4568_ ;
wire \datapath.idinstr_21_bF$buf40  ;
wire _4148_ ;
wire [31:0] \datapath.idpc_4  ;
wire [31:0] \datapath.meminstr  ;
wire _6714_ ;
wire \datapath.alu.b_0_bF$buf1  ;
wire _9186_ ;
wire _760_ ;
wire _340_ ;
wire _7919_ ;
wire _2634_ ;
wire _2214_ ;
wire \datapath.idinstr_15_bF$buf45  ;
wire _3839_ ;
wire _3419_ ;
wire _7672_ ;
wire _7252_ ;
wire _8877_ ;
wire _8457_ ;
wire _8037_ ;
wire _3592_ ;
wire _3172_ ;
wire _1905_ ;
wire _4797_ ;
wire _4377_ ;
wire _816_ ;
wire _76_ ;
wire _6943_ ;
wire _6523_ ;
wire _6103_ ;
wire _7728_ ;
wire _7308_ ;
wire _2863_ ;
wire _2443_ ;
wire _2023_ ;
wire _3648_ ;
wire _3228_ ;
wire _7481_ ;
wire _7061_ ;
wire _8686_ ;
wire _8266_ ;
wire _1714_ ;
wire _4186_ ;
wire _625_ ;
wire _205_ ;
wire _2919_ ;
wire _6752_ ;
wire _6332_ ;
wire _7957_ ;
wire _7537_ ;
wire _7117_ ;
wire _2672_ ;
wire _2252_ ;
wire _3877_ ;
wire _3457_ ;
wire _3037_ ;
wire _7290_ ;
wire _5603_ ;
wire _8495_ ;
wire _8075_ ;
wire \datapath.regcsrtrap_bF$buf5  ;
wire _6808_ ;
wire _1943_ ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire _2728_ ;
wire _2308_ ;
wire _6981_ ;
wire _6561_ ;
wire _6141_ ;
wire \datapath.alu.b_3_bF$buf4  ;
wire _7766_ ;
wire _7346_ ;
wire _2481_ ;
wire _2061_ ;
wire [31:0] \datapath.registers.1226[18]  ;
wire _3686_ ;
wire _3266_ ;
wire _5832_ ;
wire _5412_ ;
wire _6617_ ;
wire _1752_ ;
wire _1332_ ;
wire _9089_ ;
wire _663_ ;
wire _243_ ;
wire _2957_ ;
wire _2537_ ;
wire _2117_ ;
wire _6790_ ;
wire _6370_ ;
wire _7995_ ;
wire _7575_ ;
wire _7155_ ;
wire _2290_ ;
wire _3495_ ;
wire _3075_ ;
wire _9301_ ;
wire _1808_ ;
wire _5641_ ;
wire _5221_ ;
wire _719_ ;
wire _6846_ ;
wire _6426_ ;
wire _6006_ ;
wire _1981_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _2766_ ;
wire _2346_ ;
wire _5960__bF$buf0 ;
wire _5960__bF$buf1 ;
wire _5960__bF$buf2 ;
wire _5960__bF$buf3 ;
wire _5960__bF$buf4 ;
wire _4912_ ;
wire _7384_ ;
wire _8589_ ;
wire _8169_ ;
wire _9110_ ;
wire _9041__bF$buf0 ;
wire _9041__bF$buf1 ;
wire _9041__bF$buf2 ;
wire _9041__bF$buf3 ;
wire _9041__bF$buf4 ;
wire _9041__bF$buf5 ;
wire _9041__bF$buf6 ;
wire _9041__bF$buf7 ;
wire _1617_ ;
wire _4089_ ;
wire _5870_ ;
wire _5450_ ;
wire _5030_ ;
wire \datapath.idinstr_20_bF$buf28  ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _6655_ ;
wire _6235_ ;
wire _1790_ ;
wire _1370_ ;
wire _281_ ;
wire _2995_ ;
wire _2575_ ;
wire _2155_ ;
wire _8801_ ;
wire _4721_ ;
wire _4301_ ;
wire _7193_ ;
wire \datapath.idinstr_21_bF$buf37  ;
wire _5926_ ;
wire _5506_ ;
wire _8398_ ;
wire _1846_ ;
wire _1426_ ;
wire _1006_ ;
wire _757_ ;
wire _337_ ;
wire _6884_ ;
wire _6464_ ;
wire _6044_ ;
wire \datapath.idinstr_22_hier0_bF$buf3  ;
wire \datapath._62_  ;
wire _7669_ ;
wire _7249_ ;
wire _2384_ ;
wire _8610_ ;
wire _3589_ ;
wire _3169_ ;
wire _4950_ ;
wire _4530_ ;
wire _4110_ ;
wire _5735_ ;
wire _5315_ ;
wire _1655_ ;
wire _1235_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire _3801_ ;
wire _6693_ ;
wire _6273_ ;
wire _7898_ ;
wire _7478_ ;
wire _7058_ ;
wire _2193_ ;
wire _3398_ ;
wire _9204_ ;
wire _5964_ ;
wire _5544_ ;
wire _5124_ ;
wire _5432__bF$buf0 ;
wire _5432__bF$buf1 ;
wire _5432__bF$buf2 ;
wire _5432__bF$buf3 ;
wire _5432__bF$buf4 ;
wire _6749_ ;
wire _5432__bF$buf5 ;
wire _6329_ ;
wire _5432__bF$buf6 ;
wire _5432__bF$buf7 ;
wire _5432__bF$buf8 ;
wire _1884_ ;
wire _5432__bF$buf9 ;
wire _1464_ ;
wire _1044_ ;
wire _795_ ;
wire _375_ ;
wire _2669_ ;
wire _2249_ ;
wire _3610_ ;
wire _6082_ ;
wire _4815_ ;
wire _7287_ ;
wire _9433_ ;
wire _9013_ ;
wire _5773_ ;
wire _5353_ ;
wire [31:0] \datapath.wbpc_4  ;
wire _6978_ ;
wire _6558_ ;
wire _6138_ ;
wire _1693_ ;
wire _1273_ ;
wire _184_ ;
wire _2898_ ;
wire _2478_ ;
wire _2058_ ;
wire _8704_ ;
wire _4624_ ;
wire _4204_ ;
wire _7096_ ;
wire _5829_ ;
wire _5409_ ;
wire \datapath.idinstr_16_hier0_bF$buf0  ;
wire _9242_ ;
wire _1749_ ;
wire _1329_ ;
wire _5582_ ;
wire _5162_ ;
wire _6787_ ;
wire _6367_ ;
wire _1082_ ;
wire _2287_ ;
wire _8933_ ;
wire _8513_ ;
wire _4853_ ;
wire _4433_ ;
wire _4013_ ;
wire _5638_ ;
wire _5218_ ;
wire _9051_ ;
wire _1978_ ;
wire _1558_ ;
wire _1138_ ;
wire _5391_ ;
wire _889_ ;
wire _469_ ;
wire _3704_ ;
wire _6596_ ;
wire _6176_ ;
wire _4909_ ;
wire _2096_ ;
wire _8742_ ;
wire _8322_ ;
wire _9107_ ;
wire _4662_ ;
wire _4242_ ;
wire _5867_ ;
wire _5447_ ;
wire _5027_ ;
wire _9280_ ;
wire _1787_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _3933_ ;
wire _3513_ ;
wire _4718_ ;
wire \datapath.idinstr_16_bF$buf4  ;
wire _8971_ ;
wire _8551_ ;
wire _8131_ ;
wire _9336_ ;
wire _4891_ ;
wire _4471_ ;
wire _4051_ ;
wire _910_ ;
wire _5676_ ;
wire _5256_ ;
wire _1596_ ;
wire _1176_ ;
wire _7822_ ;
wire _7402_ ;
wire _8607_ ;
wire _3742_ ;
wire _3322_ ;
wire _4947_ ;
wire \datapath.idinstr_20_bF$buf4  ;
wire _4527_ ;
wire _4107_ ;
wire _8780_ ;
wire _8360_ ;
wire _9145_ ;
wire _4280_ ;
wire _5485_ ;
wire _5065_ ;
wire [31:0] \datapath.programcounter._1_  ;
wire _7631_ ;
wire _7211_ ;
wire _8836_ ;
wire _8416_ ;
wire _3971_ ;
wire _3551_ ;
wire _3131_ ;
wire _6040__bF$buf0 ;
wire _6040__bF$buf1 ;
wire _6040__bF$buf2 ;
wire _6040__bF$buf3 ;
wire _6040__bF$buf4 ;
wire _4756_ ;
wire _4336_ ;
wire \datapath.idinstr_16_bF$buf13  ;
wire _35_ ;
wire _6902_ ;
wire _9374_ ;
wire _2822_ ;
wire _2402_ ;
wire _5294_ ;
wire _3607_ ;
wire _6499_ ;
wire _6079_ ;
wire _7860_ ;
wire _7440_ ;
wire _7020_ ;
wire _8645_ ;
wire _8225_ ;
wire _3780_ ;
wire _3360_ ;
wire \datapath.idinstr_17_bF$buf22  ;
wire _4985_ ;
wire _4565_ ;
wire _4145_ ;
wire _6711_ ;
wire _9183_ ;
wire _7916_ ;
wire _2631_ ;
wire _2211_ ;
wire \datapath.idinstr_15_bF$buf42  ;
wire _3836_ ;
wire _3416_ ;
wire _8874_ ;
wire _8454_ ;
wire _8034_ ;
wire _1902_ ;
wire _9239_ ;
wire _4794_ ;
wire _4374_ ;
wire \datapath.idinstr_23_bF$buf7  ;
wire _813_ ;
wire _5999_ ;
wire _5579_ ;
wire _5159_ ;
wire _73_ ;
wire _6940_ ;
wire _6520_ ;
wire _6100_ ;
wire _1499_ ;
wire _1079_ ;
wire _7725_ ;
wire _7305_ ;
wire _2860_ ;
wire _2440_ ;
wire _2020_ ;
wire _3645_ ;
wire _3225_ ;
wire _8683_ ;
wire _8263_ ;
wire _1711_ ;
wire _9048_ ;
wire _4183_ ;
wire _622_ ;
wire _202_ ;
wire _2916_ ;
wire _5388_ ;
wire _7954_ ;
wire _7534_ ;
wire _7114_ ;
wire _8739_ ;
wire _8319_ ;
wire _3874_ ;
wire _3454_ ;
wire _3034_ ;
wire _4659_ ;
wire _4239_ ;
wire _5600_ ;
wire _8492_ ;
wire _8072_ ;
wire \datapath.regcsrtrap_bF$buf2  ;
wire _6805_ ;
wire _1940_ ;
wire _1520_ ;
wire _1100_ ;
wire _9277_ ;
wire _851_ ;
wire _431_ ;
wire _2725_ ;
wire _2305_ ;
wire _5197_ ;
wire \datapath.alu.b_3_bF$buf1  ;
wire _7763_ ;
wire _7343_ ;
wire _8968_ ;
wire _8548_ ;
wire _8128_ ;
wire \datapath.regwbtrap  ;
wire _3683_ ;
wire _3263_ ;
wire _4888_ ;
wire _4468_ ;
wire _4048_ ;
wire _907_ ;
wire _6614_ ;
wire _9086_ ;
wire _660_ ;
wire _240_ ;
wire _7819_ ;
wire _2954_ ;
wire _2534_ ;
wire _2114_ ;
wire _3739_ ;
wire _3319_ ;
wire _7992_ ;
wire _7572_ ;
wire _7152_ ;
wire _8777_ ;
wire _8357_ ;
wire _3492_ ;
wire _3072_ ;
wire _297__bF$buf0 ;
wire _297__bF$buf1 ;
wire _297__bF$buf2 ;
wire _297__bF$buf3 ;
wire _297__bF$buf4 ;
wire _297__bF$buf5 ;
wire _297__bF$buf6 ;
wire _297__bF$buf7 ;
wire _297__bF$buf8 ;
wire _1805_ ;
wire _4697_ ;
wire _4277_ ;
wire _716_ ;
wire _6843_ ;
wire _6423_ ;
wire _6003_ ;
wire _7628_ ;
wire _7208_ ;
wire _2763_ ;
wire _2343_ ;
wire _3968_ ;
wire _3548_ ;
wire _3128_ ;
wire _7381_ ;
wire _8586_ ;
wire _8166_ ;
wire _1614_ ;
wire _4086_ ;
wire \datapath.idinstr_20_bF$buf25  ;
wire _4192__bF$buf0 ;
wire _945_ ;
wire _4192__bF$buf1 ;
wire _525_ ;
wire _4192__bF$buf2 ;
wire _105_ ;
wire _4192__bF$buf3 ;
wire _4192__bF$buf4 ;
wire _2819_ ;
wire _6652_ ;
wire _6232_ ;
wire _7857_ ;
wire _7437_ ;
wire _7017_ ;
wire _2992_ ;
wire _2572_ ;
wire _2152_ ;
wire _3777_ ;
wire _3357_ ;
wire \datapath.idinstr_17_bF$buf19  ;
wire _7190_ ;
wire \datapath.idinstr_21_bF$buf34  ;
wire _5432__bF$buf10 ;
wire _5923_ ;
wire _5503_ ;
wire _8395_ ;
wire _6708_ ;
wire _1843_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire _2628_ ;
wire _2208_ ;
wire _6881_ ;
wire _6461_ ;
wire _6041_ ;
wire \datapath.idinstr_15_bF$buf39  ;
wire \datapath.idinstr_22_hier0_bF$buf0  ;
wire \datapath.idinstr_22_bF$buf43  ;
wire _7666_ ;
wire _7246_ ;
wire _2381_ ;
wire _3586_ ;
wire _3166_ ;
wire _5732_ ;
wire _5312_ ;
wire _6937_ ;
wire _6517_ ;
wire _1652_ ;
wire _1232_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _2857_ ;
wire _2437_ ;
wire _2017_ ;
wire _6690_ ;
wire _6270_ ;
wire [31:0] \datapath.mempc_4  ;
wire _7895_ ;
wire _7475_ ;
wire _7055_ ;
wire _2190_ ;
wire _3395_ ;
wire _9201_ ;
wire _1708_ ;
wire _5961_ ;
wire _5541_ ;
wire _5121_ ;
wire _619_ ;
wire _6746_ ;
wire _6326_ ;
wire _1881_ ;
wire _1461_ ;
wire _1041_ ;
wire _792_ ;
wire _372_ ;
wire _2666_ ;
wire _2246_ ;
wire _5648__bF$buf0 ;
wire _5648__bF$buf1 ;
wire _5648__bF$buf2 ;
wire _5648__bF$buf3 ;
wire _5648__bF$buf4 ;
wire _4812_ ;
wire _7284_ ;
wire [31:0] \datapath.registers.1226[9]  ;
wire _8489_ ;
wire _8069_ ;
wire _9430_ ;
wire _9010_ ;
wire _1937_ ;
wire _1517_ ;
wire _5770_ ;
wire _5350_ ;
wire _848_ ;
wire _428_ ;
wire _6975_ ;
wire _6555_ ;
wire _6135_ ;
wire _1690_ ;
wire _1270_ ;
wire _181_ ;
wire _2895_ ;
wire _2475_ ;
wire _2055_ ;
wire _8701_ ;
wire _4621_ ;
wire _4201_ ;
wire \datapath.alu.b_0_bF$buf10  ;
wire _7093_ ;
wire _5826_ ;
wire _5406_ ;
wire _8298_ ;
wire _1746_ ;
wire _1326_ ;
wire _657_ ;
wire _237_ ;
wire _7611__bF$buf10 ;
wire _6784_ ;
wire _6364_ ;
wire \datapath._52_  ;
wire _7989_ ;
wire _7569_ ;
wire _7149_ ;
wire _2284_ ;
wire _8930_ ;
wire _8510_ ;
wire _3489_ ;
wire _3069_ ;
wire _4850_ ;
wire _4430_ ;
wire _4010_ ;
wire _5635_ ;
wire _5215_ ;
wire _1975_ ;
wire _1555_ ;
wire _1135_ ;
wire _886_ ;
wire _466_ ;
wire _3701_ ;
wire _6593_ ;
wire _6173_ ;
wire _4906_ ;
wire _7798_ ;
wire _7378_ ;
wire _2093_ ;
wire _3298_ ;
wire _9104_ ;
wire _5864_ ;
wire _5444_ ;
wire _5024_ ;
wire _6649_ ;
wire _6229_ ;
wire _1784_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _2989_ ;
wire _2569_ ;
wire _2149_ ;
wire _3930_ ;
wire _3510_ ;
wire _4715_ ;
wire _7187_ ;
wire \datapath.idinstr_16_bF$buf1  ;
wire _9333_ ;
wire _5673_ ;
wire _5253_ ;
wire _6878_ ;
wire _6458_ ;
wire _6038_ ;
wire _1593_ ;
wire _1173_ ;
wire _2798_ ;
wire _2378_ ;
wire _8604_ ;
wire _4944_ ;
wire \datapath.idinstr_20_bF$buf1  ;
wire _4524_ ;
wire _4104_ ;
wire _5729_ ;
wire _5309_ ;
wire _9142_ ;
wire _1649_ ;
wire _1229_ ;
wire _5482_ ;
wire _5062_ ;
wire _498__bF$buf0 ;
wire _498__bF$buf1 ;
wire _498__bF$buf2 ;
wire _498__bF$buf3 ;
wire _498__bF$buf4 ;
wire _6687_ ;
wire _6267_ ;
wire _2187_ ;
wire _8833_ ;
wire _8413_ ;
wire _4753_ ;
wire _4333_ ;
wire _5958_ ;
wire _5538_ ;
wire _5118_ ;
wire \datapath.idinstr_16_bF$buf10  ;
wire _32_ ;
wire _9371_ ;
wire _1878_ ;
wire _1458_ ;
wire _1038_ ;
wire _5291_ ;
wire _789_ ;
wire _369_ ;
wire \datapath.idinstr_17_hier0_bF$buf4  ;
wire _3604_ ;
wire _6496_ ;
wire _6076_ ;
wire _596__bF$buf0 ;
wire _596__bF$buf1 ;
wire _596__bF$buf2 ;
wire _596__bF$buf3 ;
wire _596__bF$buf4 ;
wire _4809_ ;
wire _8642_ ;
wire _8222_ ;
wire _9427_ ;
wire _9007_ ;
wire _4982_ ;
wire _4562_ ;
wire _4142_ ;
wire \datapath.idinstr_19_bF$buf4  ;
wire _5767_ ;
wire _5347_ ;
wire _9180_ ;
wire _1687_ ;
wire _1267_ ;
wire _7913_ ;
wire _598_ ;
wire _178_ ;
wire _3833_ ;
wire _3413_ ;
wire _4618_ ;
wire _8871_ ;
wire _8451_ ;
wire _8031_ ;
wire _9236_ ;
wire _4791_ ;
wire _4371_ ;
wire \datapath.idinstr_23_bF$buf4  ;
wire _810_ ;
wire _5996_ ;
wire _5576_ ;
wire _5156_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _7722_ ;
wire _7302_ ;
wire _8927_ ;
wire _8507_ ;
wire _3642_ ;
wire _3222_ ;
wire _4847_ ;
wire _4427_ ;
wire _4007_ ;
wire _8680_ ;
wire _8260_ ;
wire _9045_ ;
wire _4180_ ;
wire _2913_ ;
wire _5385_ ;
wire _7951_ ;
wire _7531_ ;
wire _7111_ ;
wire _8736_ ;
wire _8316_ ;
wire _3871_ ;
wire _3451_ ;
wire _3031_ ;
wire _4656_ ;
wire _4236_ ;
wire _6802_ ;
wire _9274_ ;
wire _2722_ ;
wire _2302_ ;
wire _5194_ ;
wire _5454__bF$buf0 ;
wire _5454__bF$buf1 ;
wire _3927_ ;
wire _5454__bF$buf2 ;
wire _3507_ ;
wire _5454__bF$buf3 ;
wire _5454__bF$buf4 ;
wire _6399_ ;
wire _7760_ ;
wire _7340_ ;
wire _8965_ ;
wire _8545_ ;
wire _8125_ ;
wire _3680_ ;
wire _3260_ ;
wire _4885_ ;
wire _4465_ ;
wire _4045_ ;
wire _9343__bF$buf0 ;
wire _9343__bF$buf1 ;
wire _9343__bF$buf2 ;
wire _9343__bF$buf3 ;
wire _9343__bF$buf4 ;
wire _9343__bF$buf5 ;
wire _9343__bF$buf6 ;
wire _9343__bF$buf7 ;
wire _904_ ;
wire _3685__bF$buf0 ;
wire _3685__bF$buf1 ;
wire _3685__bF$buf2 ;
wire _3685__bF$buf3 ;
wire _3685__bF$buf4 ;
wire _6611_ ;
wire _9083_ ;
wire \datapath.regcondt  ;
wire _7816_ ;
wire _2951_ ;
wire _2531_ ;
wire _2111_ ;
wire [31:0] \datapath.registers.1226[23]  ;
wire _3736_ ;
wire _3316_ ;
wire \datapath.alu.b_1_bF$buf5  ;
wire _8774_ ;
wire _8354_ ;
wire _1802_ ;
wire _9139_ ;
wire _4694_ ;
wire _4274_ ;
wire _713_ ;
wire _5899_ ;
wire _5479_ ;
wire _5059_ ;
wire _6840_ ;
wire _6420_ ;
wire _6000_ ;
wire [31:0] \datapath.alu.b  ;
wire _1399_ ;
wire _7625_ ;
wire _7205_ ;
wire _2760_ ;
wire _2340_ ;
wire _3965_ ;
wire _3545_ ;
wire _3125_ ;
wire _8583_ ;
wire _8163_ ;
wire _29_ ;
wire _1611_ ;
wire _9368_ ;
wire _4083_ ;
wire \datapath.idinstr_20_bF$buf22  ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _2816_ ;
wire _5288_ ;
wire _7854_ ;
wire _7434_ ;
wire _7014_ ;
wire _8639_ ;
wire _8219_ ;
wire _3774_ ;
wire _3354_ ;
wire \datapath.idinstr_17_bF$buf16  ;
wire _4979_ ;
wire _4559_ ;
wire \datapath.idinstr_21_bF$buf31  ;
wire _4139_ ;
wire _5920_ ;
wire _5500_ ;
wire _8392_ ;
wire _6705_ ;
wire _1840_ ;
wire _1420_ ;
wire _1000_ ;
wire _9177_ ;
wire _751_ ;
wire _331_ ;
wire _2625_ ;
wire _2205_ ;
wire _5097_ ;
wire \datapath.idinstr_15_bF$buf36  ;
wire \datapath.idinstr_22_bF$buf40  ;
wire _7663_ ;
wire _7243_ ;
wire _8868_ ;
wire _8448_ ;
wire _8028_ ;
wire _3583_ ;
wire _3163_ ;
wire _4788_ ;
wire _4368_ ;
wire _807_ ;
wire \datapath.idinstr_16_bF$buf45  ;
wire _67_ ;
wire _6934_ ;
wire _6514_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _7719_ ;
wire _2854_ ;
wire _2434_ ;
wire _2014_ ;
wire _3639_ ;
wire _3219_ ;
wire _7892_ ;
wire _7472_ ;
wire _7052_ ;
wire _8677_ ;
wire _8257_ ;
wire _3392_ ;
wire _1705_ ;
wire _4597_ ;
wire _4177_ ;
wire _616_ ;
wire _6743_ ;
wire _6323_ ;
wire _7948_ ;
wire _7528_ ;
wire _7108_ ;
wire _2663_ ;
wire _2243_ ;
wire _3868_ ;
wire _3448_ ;
wire _3028_ ;
wire \datapath.csr.csr_irq  ;
wire _7281_ ;
wire _8486_ ;
wire _8066_ ;
wire _1934_ ;
wire _1514_ ;
wire _845_ ;
wire _425_ ;
wire _2719_ ;
wire _6972_ ;
wire _6552_ ;
wire _6132_ ;
wire _7757_ ;
wire _7337_ ;
wire _2892_ ;
wire _2472_ ;
wire _2052_ ;
wire _3677_ ;
wire _3257_ ;
wire _7090_ ;
wire _5823_ ;
wire _5403_ ;
wire _8295_ ;
wire _6608_ ;
wire _1743_ ;
wire _1323_ ;
wire _654_ ;
wire _234_ ;
wire _2948_ ;
wire _2528_ ;
wire _2108_ ;
wire _6781_ ;
wire _6361_ ;
wire _7986_ ;
wire _7566_ ;
wire _7146_ ;
wire _2281_ ;
wire _3486_ ;
wire _3066_ ;
wire _5632_ ;
wire _5212_ ;
wire _6837_ ;
wire _6417_ ;
wire _1972_ ;
wire _1552_ ;
wire _1132_ ;
wire _883_ ;
wire _463_ ;
wire _2757_ ;
wire _2337_ ;
wire _6590_ ;
wire _6170_ ;
wire _4903_ ;
wire _7795_ ;
wire _7375_ ;
wire _2090_ ;
wire _3295_ ;
wire _9101_ ;
wire _1608_ ;
wire _5861_ ;
wire _5441_ ;
wire _5021_ ;
wire \datapath.idinstr_20_bF$buf19  ;
wire _939_ ;
wire _519_ ;
wire _6646_ ;
wire _6226_ ;
wire _1781_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _2986_ ;
wire _2566_ ;
wire _2146_ ;
wire _4712_ ;
wire _7184_ ;
wire \datapath.idinstr_21_bF$buf28  ;
wire _5917_ ;
wire _8389_ ;
wire _9330_ ;
wire _1837_ ;
wire _1417_ ;
wire _5670_ ;
wire _5250_ ;
wire _748_ ;
wire _328_ ;
wire _6875_ ;
wire _6455_ ;
wire _6035_ ;
wire _1590_ ;
wire _1170_ ;
wire \datapath.idinstr_22_bF$buf37  ;
wire _2795_ ;
wire _2375_ ;
wire _8601_ ;
wire _4941_ ;
wire _4521_ ;
wire _4101_ ;
wire \bypassandflushunit.stall_bF$buf7  ;
wire _5726_ ;
wire _5306_ ;
wire _8198_ ;
wire _1646_ ;
wire _1226_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire _6684_ ;
wire _6264_ ;
wire [31:0] \datapath.aluinstr  ;
wire _7889_ ;
wire _7469_ ;
wire _7049_ ;
wire _2184_ ;
wire _8830_ ;
wire _8410_ ;
wire _3389_ ;
wire _4750_ ;
wire _2489__bF$buf0 ;
wire _4330_ ;
wire _2489__bF$buf1 ;
wire _2489__bF$buf2 ;
wire _2489__bF$buf3 ;
wire _5438__bF$buf0 ;
wire _2489__bF$buf4 ;
wire _5438__bF$buf1 ;
wire _2489__bF$buf5 ;
wire _5438__bF$buf2 ;
wire _2489__bF$buf6 ;
wire _5438__bF$buf3 ;
wire _2489__bF$buf7 ;
wire _5438__bF$buf4 ;
wire _5955_ ;
wire _5535_ ;
wire _5115_ ;
wire _611__bF$buf0 ;
wire _611__bF$buf1 ;
wire _611__bF$buf2 ;
wire _611__bF$buf3 ;
wire _611__bF$buf4 ;
wire _1875_ ;
wire _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire \datapath.idinstr_17_hier0_bF$buf1  ;
wire _3601_ ;
wire _6493_ ;
wire _6073_ ;
wire _4806_ ;
wire _7698_ ;
wire _7278_ ;
wire _3198_ ;
wire _5442__bF$buf0 ;
wire _5442__bF$buf1 ;
wire _5442__bF$buf2 ;
wire _5442__bF$buf3 ;
wire _5442__bF$buf4 ;
wire _9424_ ;
wire _9004_ ;
wire \datapath.idinstr_19_bF$buf1  ;
wire _1238__bF$buf0 ;
wire _1238__bF$buf1 ;
wire _1238__bF$buf2 ;
wire _5764_ ;
wire _1238__bF$buf3 ;
wire _5344_ ;
wire _1238__bF$buf4 ;
wire _6969_ ;
wire _6549_ ;
wire _6129_ ;
wire _1684_ ;
wire _1264_ ;
wire _7910_ ;
wire _595_ ;
wire _175_ ;
wire _2889_ ;
wire _2469_ ;
wire _2049_ ;
wire _3830_ ;
wire _3410_ ;
wire _4615_ ;
wire _7087_ ;
wire _9233_ ;
wire \datapath.idinstr_23_bF$buf1  ;
wire _1242__bF$buf0 ;
wire _1242__bF$buf1 ;
wire _1242__bF$buf2 ;
wire _1242__bF$buf3 ;
wire _1242__bF$buf4 ;
wire _5993_ ;
wire _5573_ ;
wire _5153_ ;
wire _6778_ ;
wire _6358_ ;
wire _1493_ ;
wire _1073_ ;
wire _2698_ ;
wire _2278_ ;
wire _8924_ ;
wire _8504_ ;
wire _4844_ ;
wire _4424_ ;
wire _4004_ ;
wire _5629_ ;
wire _5209_ ;
wire _9042_ ;
wire _1969_ ;
wire _1549_ ;
wire _1129_ ;
wire _2910_ ;
wire _5382_ ;
wire _6587_ ;
wire _6167_ ;
wire _2087_ ;
wire _8733_ ;
wire _8313_ ;
wire _4653_ ;
wire _4233_ ;
wire _5858_ ;
wire _5438_ ;
wire _5018_ ;
wire _9271_ ;
wire _1778_ ;
wire _1358_ ;
wire _5191_ ;
wire _689_ ;
wire _269_ ;
wire _3924_ ;
wire _3504_ ;
wire _6396_ ;
wire _4709_ ;
wire _8962_ ;
wire _8542_ ;
wire _8122_ ;
wire _9327_ ;
wire _4882_ ;
wire _4462_ ;
wire _4042_ ;
wire _901_ ;
wire _5667_ ;
wire _5247_ ;
wire _9080_ ;
wire _1587_ ;
wire _1167_ ;
wire _7813_ ;
wire _498_ ;
wire _3733_ ;
wire _3313_ ;
wire \datapath.alu.b_1_bF$buf2  ;
wire _4938_ ;
wire _4518_ ;
wire _8771_ ;
wire _8351_ ;
wire _9136_ ;
wire _4691_ ;
wire _4271_ ;
wire _710_ ;
wire _5896_ ;
wire _5476_ ;
wire _5056_ ;
wire _1396_ ;
wire _7622_ ;
wire _7202_ ;
wire _8827_ ;
wire _8407_ ;
wire _3962_ ;
wire _3542_ ;
wire _3122_ ;
wire _4747_ ;
wire _4327_ ;
wire _8580_ ;
wire _8160_ ;
wire _26_ ;
wire _9365_ ;
wire _4080_ ;
wire _2813_ ;
wire _5285_ ;
wire _7851_ ;
wire _7431_ ;
wire _7011_ ;
wire _8636_ ;
wire _8216_ ;
wire _3771_ ;
wire _3351_ ;
wire \datapath.idinstr_17_bF$buf13  ;
wire _4976_ ;
wire _4556_ ;
wire _4136_ ;
wire _6702_ ;
wire _9174_ ;
wire _7907_ ;
wire _2622_ ;
wire _2202_ ;
wire _5094_ ;
wire \datapath.idinstr_15_bF$buf33  ;
wire _3827_ ;
wire _3407_ ;
wire _6299_ ;
wire _7660_ ;
wire _7240_ ;
wire _8865_ ;
wire _8445_ ;
wire _8025_ ;
wire _3580_ ;
wire _3160_ ;
wire _4785_ ;
wire _4365_ ;
wire _804_ ;
wire \datapath.idinstr_16_bF$buf42  ;
wire _64_ ;
wire _6931_ ;
wire _6511_ ;
wire _7716_ ;
wire _2851_ ;
wire _2431_ ;
wire _2011_ ;
wire [31:0] \datapath.registers.1226[13]  ;
wire _3636_ ;
wire _3216_ ;
wire _8674_ ;
wire _8254_ ;
wire \controlunit.csrfile_trap_wen  ;
wire _1702_ ;
wire _9039_ ;
wire _4594_ ;
wire _4174_ ;
wire _613_ ;
wire _2907_ ;
wire _5799_ ;
wire _5379_ ;
wire _6740_ ;
wire _6320_ ;
wire _1299_ ;
wire _7945_ ;
wire _7525_ ;
wire _7105_ ;
wire _2660_ ;
wire _2240_ ;
wire _3865_ ;
wire _3445_ ;
wire _3025_ ;
wire _8483_ ;
wire CLK_bF$buf90 ;
wire _8063_ ;
wire CLK_bF$buf91 ;
wire CLK_bF$buf92 ;
wire CLK_bF$buf93 ;
wire CLK_bF$buf94 ;
wire CLK_bF$buf95 ;
wire CLK_bF$buf96 ;
wire CLK_bF$buf97 ;
wire CLK_bF$buf98 ;
wire CLK_bF$buf99 ;
wire _1931_ ;
wire _1511_ ;
wire _9268_ ;
wire _842_ ;
wire _422_ ;
wire _2716_ ;
wire _5188_ ;
wire _7754_ ;
wire _7334_ ;
wire _8959_ ;
wire _8539_ ;
wire _8119_ ;
wire _3674_ ;
wire _3254_ ;
wire _4879_ ;
wire _4459_ ;
wire _4039_ ;
wire _5820_ ;
wire _5400_ ;
wire _8292_ ;
wire _6605_ ;
wire _1740_ ;
wire _1320_ ;
wire _9077_ ;
wire _651_ ;
wire _231_ ;
wire _2945_ ;
wire _2525_ ;
wire _2105_ ;
wire _7983_ ;
wire _7563_ ;
wire _7143_ ;
wire _8768_ ;
wire _8348_ ;
wire _3483_ ;
wire _3063_ ;
wire _4688_ ;
wire _4268_ ;
wire _707_ ;
wire _6834_ ;
wire _6414_ ;
wire \controlunit.ecall  ;
wire _880_ ;
wire _460_ ;
wire _7619_ ;
wire _2754_ ;
wire _2334_ ;
wire _3959_ ;
wire _3539_ ;
wire _3119_ ;
wire _4900_ ;
wire _7792_ ;
wire _7372_ ;
wire _4198__bF$buf0 ;
wire _4198__bF$buf1 ;
wire _4198__bF$buf2 ;
wire _8997_ ;
wire _4198__bF$buf3 ;
wire _8577_ ;
wire _4198__bF$buf4 ;
wire _8157_ ;
wire _3292_ ;
wire _1605_ ;
wire _4497_ ;
wire _4077_ ;
wire \datapath.idinstr_20_bF$buf16  ;
wire _936_ ;
wire _516_ ;
wire _6643_ ;
wire _6223_ ;
wire _7848_ ;
wire _7428_ ;
wire _7008_ ;
wire _2983_ ;
wire _2563_ ;
wire _2143_ ;
wire _3768_ ;
wire _3348_ ;
wire _7181_ ;
wire \datapath.idinstr_21_bF$buf25  ;
wire _5914_ ;
wire _8386_ ;
wire _1834_ ;
wire _1414_ ;
wire _745_ ;
wire _325_ ;
wire _2619_ ;
wire _6872_ ;
wire _6452_ ;
wire _6032_ ;
wire \datapath.idinstr_22_bF$buf34  ;
wire _7657_ ;
wire _7237_ ;
wire _2792_ ;
wire _2372_ ;
wire _3997_ ;
wire _3577_ ;
wire _3157_ ;
wire \bypassandflushunit.stall_bF$buf4  ;
wire _5723_ ;
wire _5303_ ;
wire _8195_ ;
wire \datapath.idinstr_16_bF$buf39  ;
wire _6928_ ;
wire _6508_ ;
wire _1643_ ;
wire _1223_ ;
wire \datapath.idinstr_20_bF$buf54  ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire _2848_ ;
wire _2428_ ;
wire _2008_ ;
wire _6681_ ;
wire _6261_ ;
wire _7886_ ;
wire _7466_ ;
wire _7046_ ;
wire _2181_ ;
wire _3386_ ;
wire _5952_ ;
wire _5532_ ;
wire _5112_ ;
wire _6737_ ;
wire _6317_ ;
wire _1872_ ;
wire _1452_ ;
wire _1032_ ;
wire _783_ ;
wire _363_ ;
wire _2657_ ;
wire _2237_ ;
wire _6490_ ;
wire _6070_ ;
wire _4803_ ;
wire _7695_ ;
wire _7275_ ;
wire _3195_ ;
wire _9421_ ;
wire _9001_ ;
wire _1928_ ;
wire _1508_ ;
wire _5761_ ;
wire _5341_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _6966_ ;
wire _6546_ ;
wire _6126_ ;
wire _1681_ ;
wire _1261_ ;
wire _592_ ;
wire _172_ ;
wire _2886_ ;
wire _2466_ ;
wire _2046_ ;
wire _4612_ ;
wire _7084_ ;
wire _5817_ ;
wire _8289_ ;
wire _9230_ ;
wire _1737_ ;
wire _1317_ ;
wire _5990_ ;
wire _5570_ ;
wire _5150_ ;
wire _648_ ;
wire _228_ ;
wire _6775_ ;
wire _6355_ ;
wire _1490_ ;
wire _1070_ ;
wire _2695_ ;
wire _2275_ ;
wire _8921_ ;
wire _8501_ ;
wire _4841_ ;
wire _4421_ ;
wire _4001_ ;
wire _5626_ ;
wire _5206_ ;
wire _8098_ ;
wire _1966_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire _614__bF$buf0 ;
wire _614__bF$buf1 ;
wire _614__bF$buf2 ;
wire _614__bF$buf3 ;
wire _614__bF$buf4 ;
wire _6584_ ;
wire _6164_ ;
wire _5760__bF$buf0 ;
wire _5760__bF$buf1 ;
wire _5760__bF$buf2 ;
wire _5760__bF$buf3 ;
wire _5760__bF$buf4 ;
wire _5760__bF$buf5 ;
wire _5760__bF$buf6 ;
wire _5760__bF$buf7 ;
wire _5760__bF$buf8 ;
wire [1:0] \datapath._32_  ;
wire _7789_ ;
wire _7369_ ;
wire _2084_ ;
wire _8730_ ;
wire _8310_ ;
wire \datapath.immediatedecoder._12_  ;
wire _3289_ ;
wire _4650_ ;
wire _4230_ ;
wire _5855_ ;
wire _5435_ ;
wire _5015_ ;
wire _1775_ ;
wire _1355_ ;
wire _686_ ;
wire [31:0] \datapath.imm  ;
wire _266_ ;
wire _3921_ ;
wire _3501_ ;
wire _6393_ ;
wire _4706_ ;
wire _7598_ ;
wire _7178_ ;
wire _3098_ ;
wire _9324_ ;
wire [31:0] \datapath.regimmalu  ;
wire _5664_ ;
wire _5244_ ;
wire \datapath.idinstr_17_bF$buf7  ;
wire _965__bF$buf0 ;
wire _965__bF$buf1 ;
wire _965__bF$buf2 ;
wire _965__bF$buf3 ;
wire _965__bF$buf4 ;
wire _6869_ ;
wire _6449_ ;
wire _6029_ ;
wire _1584_ ;
wire _1164_ ;
wire _7810_ ;
wire CLK ;
wire _495_ ;
wire _2789_ ;
wire _2369_ ;
wire _3730_ ;
wire _3310_ ;
wire _4935_ ;
wire _4515_ ;
wire _9133_ ;
wire \datapath.idinstr_21_bF$buf7  ;
wire _5893_ ;
wire _5473_ ;
wire _5053_ ;
wire _6678_ ;
wire _6258_ ;
wire _1393_ ;
wire _2598_ ;
wire _2178_ ;
wire _8824_ ;
wire _8404_ ;
wire _4744_ ;
wire _4324_ ;
wire _5949_ ;
wire _5529_ ;
wire _5109_ ;
wire _23_ ;
wire _9362_ ;
wire _1869_ ;
wire _1449_ ;
wire _1029_ ;
wire _2810_ ;
wire _5894__bF$buf0 ;
wire _5894__bF$buf1 ;
wire _5894__bF$buf2 ;
wire _5894__bF$buf3 ;
wire _5894__bF$buf4 ;
wire _5894__bF$buf5 ;
wire _5894__bF$buf6 ;
wire _5894__bF$buf7 ;
wire _5282_ ;
wire _5894__bF$buf8 ;
wire _6487_ ;
wire _6067_ ;
wire _8633_ ;
wire _8213_ ;
wire \datapath.idinstr_17_bF$buf10  ;
wire _3463__bF$buf0 ;
wire _3463__bF$buf1 ;
wire _3463__bF$buf2 ;
wire _3463__bF$buf3 ;
wire _3463__bF$buf4 ;
wire _3463__bF$buf5 ;
wire _3463__bF$buf6 ;
wire _9418_ ;
wire _4973_ ;
wire _4553_ ;
wire _4133_ ;
wire _5758_ ;
wire _5338_ ;
wire _9171_ ;
wire _1678_ ;
wire _1258_ ;
wire _7904_ ;
wire _5091_ ;
wire _589_ ;
wire _169_ ;
wire \datapath.idinstr_15_bF$buf30  ;
wire _3824_ ;
wire _3404_ ;
wire _6296_ ;
wire _4609_ ;
wire _8862_ ;
wire _8442_ ;
wire _8022_ ;
wire \datapath.alu.b_4_bF$buf2  ;
wire _9227_ ;
wire _4782_ ;
wire _4362_ ;
wire _801_ ;
wire _5987_ ;
wire _5567_ ;
wire _5147_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _7713_ ;
wire _398_ ;
wire _8918_ ;
wire _3633_ ;
wire _3213_ ;
wire _4838_ ;
wire _4418_ ;
wire _8671_ ;
wire _8251_ ;
wire _9036_ ;
wire _4591_ ;
wire _4171_ ;
wire _610_ ;
wire _2904_ ;
wire _5681__bF$buf0 ;
wire _5681__bF$buf1 ;
wire _5681__bF$buf2 ;
wire _5681__bF$buf3 ;
wire _5681__bF$buf4 ;
wire _5796_ ;
wire _5376_ ;
wire _1296_ ;
wire _7942_ ;
wire _7522_ ;
wire _7102_ ;
wire _8727_ ;
wire _8307_ ;
wire _3862_ ;
wire _3442_ ;
wire _3022_ ;
wire _3250__bF$buf0 ;
wire _3250__bF$buf1 ;
wire _3250__bF$buf2 ;
wire _3250__bF$buf3 ;
wire _3250__bF$buf4 ;
wire _3250__bF$buf5 ;
wire _4647_ ;
wire _4227_ ;
wire [14:0] \datapath._49_  ;
wire _8480_ ;
wire CLK_bF$buf60 ;
wire _8060_ ;
wire CLK_bF$buf61 ;
wire CLK_bF$buf62 ;
wire CLK_bF$buf63 ;
wire CLK_bF$buf64 ;
wire CLK_bF$buf65 ;
wire CLK_bF$buf66 ;
wire CLK_bF$buf67 ;
wire CLK_bF$buf68 ;
wire CLK_bF$buf69 ;
wire _9265_ ;
wire _2713_ ;
wire _5185_ ;
wire [31:0] \datapath.rd  ;
wire _3918_ ;
wire _7751_ ;
wire _7331_ ;
wire _8956_ ;
wire _8536_ ;
wire _8116_ ;
wire _3671_ ;
wire _3251_ ;
wire _4876_ ;
wire _4456_ ;
wire _4036_ ;
wire _5464__bF$buf0 ;
wire _5464__bF$buf1 ;
wire _5464__bF$buf2 ;
wire _5464__bF$buf3 ;
wire _6602_ ;
wire _5464__bF$buf4 ;
wire _9074_ ;
wire _7807_ ;
wire _2942_ ;
wire _2522_ ;
wire _2102_ ;
wire _3727_ ;
wire _3307_ ;
wire _6199_ ;
wire _7980_ ;
wire _7560_ ;
wire _7140_ ;
wire _8765_ ;
wire _8345_ ;
wire _3480_ ;
wire _3060_ ;
wire _4685_ ;
wire _4265_ ;
wire _704_ ;
wire _6831_ ;
wire _6411_ ;
wire _7616_ ;
wire _2751_ ;
wire _2331_ ;
wire _3956_ ;
wire _3536_ ;
wire _3116_ ;
wire _8994_ ;
wire _8574_ ;
wire _8154_ ;
wire _1602_ ;
wire _9359_ ;
wire _4494_ ;
wire _4074_ ;
wire \datapath.idinstr_20_bF$buf13  ;
wire _933_ ;
wire _513_ ;
wire _2807_ ;
wire _5699_ ;
wire _5279_ ;
wire _6640_ ;
wire _6220_ ;
wire _1199_ ;
wire _7845_ ;
wire _7425_ ;
wire _7005_ ;
wire _2980_ ;
wire _2560_ ;
wire _2140_ ;
wire _3765_ ;
wire _3345_ ;
wire \datapath.idinstr_21_bF$buf22  ;
wire _5911_ ;
wire _8383_ ;
wire _1831_ ;
wire _1411_ ;
wire _9168_ ;
wire _742_ ;
wire _322_ ;
wire _2616_ ;
wire _5088_ ;
wire \datapath.idinstr_15_bF$buf27  ;
wire \datapath.idinstr_22_bF$buf31  ;
wire _7654_ ;
wire _7234_ ;
wire [31:0] \datapath.registers.1226[4]  ;
wire _8859_ ;
wire _8439_ ;
wire _8019_ ;
wire _3994_ ;
wire _3574_ ;
wire _3154_ ;
wire [31:0] IMEM_ADDR ;
wire \bypassandflushunit.stall_bF$buf1  ;
wire _4779_ ;
wire _4359_ ;
wire _5720_ ;
wire _5300_ ;
wire _8192_ ;
wire \datapath.idinstr_16_bF$buf36  ;
wire _58_ ;
wire _6925_ ;
wire _6505_ ;
wire _1640_ ;
wire _1220_ ;
wire _6144__bF$buf10 ;
wire _9397_ ;
wire \datapath.idinstr_20_bF$buf51  ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _2845_ ;
wire _2425_ ;
wire _2005_ ;
wire _7883_ ;
wire _7463_ ;
wire _7043_ ;
wire _8668_ ;
wire _8248_ ;
wire _3383_ ;
wire _4588_ ;
wire _4168_ ;
wire _607_ ;
wire _6734_ ;
wire _6314_ ;
wire _780_ ;
wire _360_ ;
wire _7939_ ;
wire _7519_ ;
wire _2654_ ;
wire _2234_ ;
wire _3859_ ;
wire _3439_ ;
wire _3019_ ;
wire _4800_ ;
wire _7692_ ;
wire _7272_ ;
wire _8897_ ;
wire _8477_ ;
wire _8057_ ;
wire _3192_ ;
wire _1925_ ;
wire _1505_ ;
wire [3:0] \datapath.excpt_cause  ;
wire _4397_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _6963_ ;
wire _6543_ ;
wire _6123_ ;
wire _7748_ ;
wire _7328_ ;
wire _2883_ ;
wire _2463_ ;
wire _2043_ ;
wire _3668_ ;
wire _3248_ ;
wire _7081_ ;
wire _5814_ ;
wire _8286_ ;
wire _1734_ ;
wire _1314_ ;
wire _645_ ;
wire _225_ ;
wire _2939_ ;
wire _2519_ ;
wire _6772_ ;
wire _6352_ ;
wire _7977_ ;
wire _7557_ ;
wire _7137_ ;
wire _2692_ ;
wire _2272_ ;
wire _3897_ ;
wire _3477_ ;
wire _3057_ ;
wire _5623_ ;
wire _5203_ ;
wire _8095_ ;
wire _6828_ ;
wire _6408_ ;
wire _1963_ ;
wire _1543_ ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _2748_ ;
wire _2328_ ;
wire _6581_ ;
wire _6161_ ;
wire _7786_ ;
wire _7366_ ;
wire _2081_ ;
wire _3286_ ;
wire _5852_ ;
wire _5432_ ;
wire _5012_ ;
wire _6637_ ;
wire _6217_ ;
wire _1772_ ;
wire _1352_ ;
wire _683_ ;
wire _263_ ;
wire _2977_ ;
wire _2557_ ;
wire _2137_ ;
wire _6390_ ;
wire _4703_ ;
wire _7595_ ;
wire _7175_ ;
wire \datapath.idinstr_21_bF$buf19  ;
wire _5908_ ;
wire _3095_ ;
wire _9321_ ;
wire _1828_ ;
wire _1408_ ;
wire \bypassandflushunit.flushalu  ;
wire _5661_ ;
wire _5241_ ;
wire _739_ ;
wire _319_ ;
wire \datapath.idinstr_17_bF$buf4  ;
wire _6866_ ;
wire _6446_ ;
wire _6026_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire \datapath.idinstr_22_bF$buf28  ;
wire _2786_ ;
wire _2366_ ;
wire _4932_ ;
wire _4512_ ;
wire _5717_ ;
wire _8189_ ;
wire _9130_ ;
wire _1637_ ;
wire _1217_ ;
wire \datapath.idinstr_21_bF$buf4  ;
wire _5890_ ;
wire _5470_ ;
wire _5050_ ;
wire \datapath.idinstr_20_bF$buf48  ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _6675_ ;
wire _6255_ ;
wire _1390_ ;
wire _2595_ ;
wire _2175_ ;
wire _8821_ ;
wire _8401_ ;
wire _4741_ ;
wire _4321_ ;
wire _5946_ ;
wire _5526_ ;
wire _5106_ ;
wire _20_ ;
wire _1866_ ;
wire _1446_ ;
wire _1026_ ;
wire _6041__bF$buf0 ;
wire _6041__bF$buf1 ;
wire _6041__bF$buf2 ;
wire _6041__bF$buf3 ;
wire _6041__bF$buf4 ;
wire _6041__bF$buf5 ;
wire _6041__bF$buf6 ;
wire _6041__bF$buf7 ;
wire _6041__bF$buf8 ;
wire _777_ ;
wire _357_ ;
wire _6484_ ;
wire _6064_ ;
wire _5448__bF$buf0 ;
wire _5448__bF$buf1 ;
wire _5448__bF$buf2 ;
wire _5448__bF$buf3 ;
wire _5448__bF$buf4 ;
wire _7689_ ;
wire _7269_ ;
wire _8630_ ;
wire _8210_ ;
wire _3189_ ;
wire _9415_ ;
wire _4970_ ;
wire _4550_ ;
wire _4130_ ;
wire _5755_ ;
wire _5335_ ;
wire _1675_ ;
wire _1255_ ;
wire _7901_ ;
wire _586_ ;
wire _166_ ;
wire _3821_ ;
wire _3401_ ;
wire _5452__bF$buf0 ;
wire _6293_ ;
wire _5452__bF$buf1 ;
wire _5452__bF$buf2 ;
wire _5452__bF$buf3 ;
wire _5452__bF$buf4 ;
wire _4606_ ;
wire _7498_ ;
wire _7078_ ;
wire _9224_ ;
wire _5984_ ;
wire _5564_ ;
wire _5144_ ;
wire _6769_ ;
wire _6349_ ;
wire _1484_ ;
wire _1064_ ;
wire _7710_ ;
wire _395_ ;
wire _2689_ ;
wire _2269_ ;
wire _8915_ ;
wire [31:0] \datapath.programcounter.jumps  ;
wire _3630_ ;
wire _3210_ ;
wire _4835_ ;
wire _4415_ ;
wire _9033_ ;
wire \datapath.alu.b_2_bF$buf6  ;
wire _2901_ ;
wire _5793_ ;
wire _5373_ ;
wire _6998_ ;
wire _6578_ ;
wire _6158_ ;
wire _1293_ ;
wire _2498_ ;
wire _2078_ ;
wire _8724_ ;
wire _8304_ ;
wire _4644_ ;
wire _4224_ ;
wire CLK_bF$buf30 ;
wire CLK_bF$buf31 ;
wire CLK_bF$buf32 ;
wire CLK_bF$buf33 ;
wire CLK_bF$buf34 ;
wire CLK_bF$buf35 ;
wire CLK_bF$buf36 ;
wire CLK_bF$buf37 ;
wire CLK_bF$buf38 ;
wire CLK_bF$buf39 ;
wire _5849_ ;
wire _5429_ ;
wire _5009_ ;
wire _9262_ ;
wire _1769_ ;
wire _1349_ ;
wire _2710_ ;
wire _5182_ ;
wire _3915_ ;
wire _6387_ ;
wire _8953_ ;
wire _8533_ ;
wire _8113_ ;
wire _9318_ ;
wire _4873_ ;
wire _4453_ ;
wire _4033_ ;
wire _5658_ ;
wire _5238_ ;
wire _9071_ ;
wire _9076__bF$buf0 ;
wire _9076__bF$buf1 ;
wire _9076__bF$buf2 ;
wire _9076__bF$buf3 ;
wire _9076__bF$buf4 ;
wire _9076__bF$buf5 ;
wire _9076__bF$buf6 ;
wire _9076__bF$buf7 ;
wire _9076__bF$buf8 ;
wire _1998_ ;
wire _1578_ ;
wire _1158_ ;
wire _7804_ ;
wire _489_ ;
wire _5826__bF$buf0 ;
wire _5826__bF$buf1 ;
wire _5826__bF$buf2 ;
wire _5826__bF$buf3 ;
wire _5826__bF$buf4 ;
wire _3724_ ;
wire _3304_ ;
wire _6196_ ;
wire _4929_ ;
wire _4509_ ;
wire _8762_ ;
wire _8342_ ;
wire _9127_ ;
wire _4682_ ;
wire _4262_ ;
wire _701_ ;
wire _5887_ ;
wire _5467_ ;
wire _5047_ ;
wire _298__bF$buf0 ;
wire _298__bF$buf1 ;
wire _298__bF$buf2 ;
wire _298__bF$buf3 ;
wire _298__bF$buf4 ;
wire _1387_ ;
wire _7613_ ;
wire _298_ ;
wire \datapath.idinstr_20_hier0_bF$buf5  ;
wire _8818_ ;
wire _3953_ ;
wire _3533_ ;
wire _3113_ ;
wire _4738_ ;
wire _4318_ ;
wire _8991_ ;
wire _8571_ ;
wire _8151_ ;
wire _17_ ;
wire _9356_ ;
wire _4491_ ;
wire _4071_ ;
wire \datapath.idinstr_20_bF$buf10  ;
wire _930_ ;
wire _510_ ;
wire _2804_ ;
wire _5696_ ;
wire _5276_ ;
wire _1196_ ;
wire _7842_ ;
wire _7422_ ;
wire _7002_ ;
wire _8627_ ;
wire _8207_ ;
wire _3762_ ;
wire _3342_ ;
wire _4967_ ;
wire _4547_ ;
wire _4127_ ;
wire _8380_ ;
wire _9165_ ;
wire _2613_ ;
wire _5085_ ;
wire \datapath.idinstr_15_bF$buf24  ;
wire _3818_ ;
wire _7651_ ;
wire _7231_ ;
wire _8856_ ;
wire _8436_ ;
wire _8016_ ;
wire _3991_ ;
wire _3571_ ;
wire _3151_ ;
wire _4776_ ;
wire _4356_ ;
wire \datapath.idinstr_16_bF$buf33  ;
wire _55_ ;
wire _6922_ ;
wire _6502_ ;
wire _9394_ ;
wire _7707_ ;
wire _2842_ ;
wire _2422_ ;
wire _2002_ ;
wire _3627_ ;
wire _3207_ ;
wire _6099_ ;
wire _7880_ ;
wire _7460_ ;
wire _7040_ ;
wire _8665_ ;
wire _8245_ ;
wire _3380_ ;
wire _4585_ ;
wire _4165_ ;
wire _604_ ;
wire _6731_ ;
wire _6311_ ;
wire _7936_ ;
wire _7516_ ;
wire _2651_ ;
wire _2231_ ;
wire _3856_ ;
wire _3436_ ;
wire _3016_ ;
wire _8894_ ;
wire _8474_ ;
wire _8054_ ;
wire _1922_ ;
wire _1502_ ;
wire _9259_ ;
wire _4394_ ;
wire _833_ ;
wire _413_ ;
wire _2707_ ;
wire _5599_ ;
wire _5179_ ;
wire _93_ ;
wire _6960_ ;
wire _6540_ ;
wire _6120_ ;
wire _1099_ ;
wire _7745_ ;
wire _7325_ ;
wire _2880_ ;
wire _2460_ ;
wire _2040_ ;
wire _3665_ ;
wire _3245_ ;
wire _5811_ ;
wire _8283_ ;
wire _1731_ ;
wire _1311_ ;
wire _9068_ ;
wire _642_ ;
wire _222_ ;
wire _2936_ ;
wire _2516_ ;
wire _7974_ ;
wire _7554_ ;
wire _7134_ ;
wire _8759_ ;
wire _8339_ ;
wire _3894_ ;
wire _3474_ ;
wire _3054_ ;
wire _4679_ ;
wire _4259_ ;
wire _5620_ ;
wire _5200_ ;
wire _8092_ ;
wire _6825_ ;
wire _6405_ ;
wire _1960_ ;
wire _1540_ ;
wire _1120_ ;
wire _9297_ ;
wire _871_ ;
wire _451_ ;
wire _2745_ ;
wire _2325_ ;
wire _7783_ ;
wire _7363_ ;
wire _8988_ ;
wire _8568_ ;
wire _8148_ ;
wire _3283_ ;
wire _4488_ ;
wire _4068_ ;
wire _927_ ;
wire _507_ ;
wire _6634_ ;
wire _6214_ ;
wire _680_ ;
wire _260_ ;
wire _7839_ ;
wire _7419_ ;
wire _2974_ ;
wire _2554_ ;
wire _2134_ ;
wire _3759_ ;
wire _3339_ ;
wire _4700_ ;
wire _7592_ ;
wire _7172_ ;
wire \datapath.idinstr_21_bF$buf16  ;
wire _5905_ ;
wire _8797_ ;
wire _8377_ ;
wire _3092_ ;
wire _1825_ ;
wire _1405_ ;
wire _4297_ ;
wire _736_ ;
wire _316_ ;
wire \datapath.idinstr_17_bF$buf1  ;
wire _6863_ ;
wire _6443_ ;
wire _6023_ ;
wire [31:0] \datapath.rs2bypass  ;
wire \datapath.idinstr_22_bF$buf25  ;
wire _7648_ ;
wire _7228_ ;
wire _2783_ ;
wire _2363_ ;
wire _3988_ ;
wire _3568_ ;
wire _3148_ ;
wire _9277__bF$buf0 ;
wire _9277__bF$buf1 ;
wire _9277__bF$buf2 ;
wire _9277__bF$buf3 ;
wire _9277__bF$buf4 ;
wire _5714_ ;
wire _8186_ ;
wire _6919_ ;
wire _1634_ ;
wire _1214_ ;
wire \datapath.idinstr_21_bF$buf1  ;
wire _5434__bF$buf10 ;
wire _5434__bF$buf11 ;
wire \datapath.idinstr_20_bF$buf45  ;
wire _5434__bF$buf12 ;
wire _5434__bF$buf13 ;
wire _965_ ;
wire _5434__bF$buf14 ;
wire _545_ ;
wire _125_ ;
wire _2839_ ;
wire \datapath.idinstr_15_bF$buf8  ;
wire _2419_ ;
wire _6672_ ;
wire _6252_ ;
wire _7877_ ;
wire _7457_ ;
wire _7037_ ;
wire _2592_ ;
wire _2172_ ;
wire _3797_ ;
wire _3377_ ;
wire \datapath.idinstr_17_bF$buf39  ;
wire _5943_ ;
wire _5523_ ;
wire _5103_ ;
wire _6728_ ;
wire _6308_ ;
wire _1863_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _2648_ ;
wire _2228_ ;
wire _6481_ ;
wire _6061_ ;
wire _7686_ ;
wire _7266_ ;
wire _3186_ ;
wire _9412_ ;
wire _1919_ ;
wire _597__bF$buf0 ;
wire _597__bF$buf1 ;
wire _597__bF$buf2 ;
wire _597__bF$buf3 ;
wire _597__bF$buf4 ;
wire _5752_ ;
wire _5332_ ;
wire _6957_ ;
wire _6537_ ;
wire _6117_ ;
wire _1672_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _2877_ ;
wire _2457_ ;
wire _2037_ ;
wire _6290_ ;
wire _4603_ ;
wire _7495_ ;
wire _7075_ ;
wire _5808_ ;
wire _9221_ ;
wire _1728_ ;
wire _1308_ ;
wire _5981_ ;
wire _5561_ ;
wire _5141_ ;
wire _639_ ;
wire _219_ ;
wire [31:0] DMEM_ADDR ;
wire _6766_ ;
wire _6346_ ;
wire _1481_ ;
wire _1061_ ;
wire _392_ ;
wire \datapath.idinstr_24_bF$buf4  ;
wire _2686_ ;
wire _2266_ ;
wire _8912_ ;
wire _4832_ ;
wire _4412_ ;
wire _5617_ ;
wire _8089_ ;
wire _9030_ ;
wire \datapath.alu.b_2_bF$buf3  ;
wire _1957_ ;
wire _1537_ ;
wire _1117_ ;
wire _5790_ ;
wire _5370_ ;
wire _868_ ;
wire _448_ ;
wire _6995_ ;
wire _6575_ ;
wire _6155_ ;
wire _1290_ ;
wire _2495_ ;
wire _2075_ ;
wire _8721_ ;
wire _8301_ ;
wire _4641_ ;
wire _4221_ ;
wire _5846_ ;
wire _5426_ ;
wire _5006_ ;
wire _1766_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire _3912_ ;
wire _6384_ ;
wire _7589_ ;
wire _7169_ ;
wire _8950_ ;
wire _8530_ ;
wire _8110_ ;
wire _3089_ ;
wire _9315_ ;
wire _4870_ ;
wire _4450_ ;
wire _4030_ ;
wire _5655_ ;
wire _5235_ ;
wire _1995_ ;
wire _1575_ ;
wire _1155_ ;
wire _7801_ ;
wire _486_ ;
wire _3721_ ;
wire _3301_ ;
wire _6193_ ;
wire _4926_ ;
wire _4506_ ;
wire _7398_ ;
wire _9124_ ;
wire _5884_ ;
wire _5464_ ;
wire _5044_ ;
wire _6669_ ;
wire _6249_ ;
wire _1384_ ;
wire _7610_ ;
wire _295_ ;
wire _2589_ ;
wire _3690__bF$buf0 ;
wire _2169_ ;
wire _3690__bF$buf1 ;
wire _3690__bF$buf2 ;
wire _3690__bF$buf3 ;
wire \datapath.idinstr_20_hier0_bF$buf2  ;
wire _3690__bF$buf4 ;
wire _8815_ ;
wire _3950_ ;
wire _3530_ ;
wire _3110_ ;
wire _4735_ ;
wire _4315_ ;
wire _14_ ;
wire _9353_ ;
wire _2801_ ;
wire _5693_ ;
wire _5273_ ;
wire _6898_ ;
wire _6478_ ;
wire _6058_ ;
wire _1193_ ;
wire _2398_ ;
wire _8624_ ;
wire _8204_ ;
wire _9409_ ;
wire _4964_ ;
wire _4544_ ;
wire _4124_ ;
wire _5749_ ;
wire _5329_ ;
wire _9162_ ;
wire _1669_ ;
wire _1249_ ;
wire _2610_ ;
wire _5082_ ;
wire \datapath.idinstr_15_bF$buf21  ;
wire _3815_ ;
wire _6287_ ;
wire _8853_ ;
wire _8433_ ;
wire _8013_ ;
wire _9218_ ;
wire _4773_ ;
wire _4353_ ;
wire _5978_ ;
wire _5558_ ;
wire _5138_ ;
wire \datapath.idinstr_16_bF$buf30  ;
wire _52_ ;
wire _9391_ ;
wire _1898_ ;
wire _1478_ ;
wire _1058_ ;
wire _7704_ ;
wire _389_ ;
wire _8909_ ;
wire _3624_ ;
wire _3204_ ;
wire _6096_ ;
wire _4829_ ;
wire _4409_ ;
wire _8662_ ;
wire _8242_ ;
wire _9027_ ;
wire _4582_ ;
wire _4162_ ;
wire _601_ ;
wire _5787_ ;
wire _5367_ ;
wire _1287_ ;
wire _7933_ ;
wire _7513_ ;
wire _198_ ;
wire _8718_ ;
wire _3853_ ;
wire _3433_ ;
wire _3013_ ;
wire _4638_ ;
wire _4218_ ;
wire _8891_ ;
wire _8471_ ;
wire _8051_ ;
wire _9256_ ;
wire _4391_ ;
wire _830_ ;
wire _410_ ;
wire _2704_ ;
wire _5596_ ;
wire _5176_ ;
wire _90_ ;
wire _3909_ ;
wire _1096_ ;
wire _7742_ ;
wire _7322_ ;
wire _8947_ ;
wire _8527_ ;
wire _8107_ ;
wire _3662_ ;
wire _3242_ ;
wire _4867_ ;
wire _4447_ ;
wire _4027_ ;
wire [2:0] \datapath._29_  ;
wire _8280_ ;
wire \datapath.immediatedecoder._09_  ;
wire _9065_ ;
wire _2933_ ;
wire _2513_ ;
wire _3718_ ;
wire _7971_ ;
wire _7551_ ;
wire _7131_ ;
wire _8756_ ;
wire _8336_ ;
wire _3891_ ;
wire _3471_ ;
wire _3051_ ;
wire _5474__bF$buf0 ;
wire _5474__bF$buf1 ;
wire _5474__bF$buf2 ;
wire _5474__bF$buf3 ;
wire _5474__bF$buf4 ;
wire _4676_ ;
wire _4256_ ;
wire _6822_ ;
wire _6402_ ;
wire _9294_ ;
wire _7607_ ;
wire _2742_ ;
wire _2322_ ;
wire _3947_ ;
wire _3527_ ;
wire _3107_ ;
wire _8_ ;
wire _7780_ ;
wire _7360_ ;
wire _8985_ ;
wire _8565_ ;
wire _8145_ ;
wire _3280_ ;
wire _4485_ ;
wire _4065_ ;
wire _924_ ;
wire _504_ ;
wire _6631_ ;
wire _6211_ ;
wire _7836_ ;
wire _7416_ ;
wire _2971_ ;
wire _2551_ ;
wire _2131_ ;
wire [31:0] \datapath.registers.1226[25]  ;
wire _3756_ ;
wire _3336_ ;
wire \datapath.idinstr_21_bF$buf13  ;
wire _5902_ ;
wire _8794_ ;
wire _8374_ ;
wire \datapath.regmret_bF$buf2  ;
wire _1822_ ;
wire _1402_ ;
wire _9159_ ;
wire _4294_ ;
wire _733_ ;
wire _313_ ;
wire _2607_ ;
wire _5499_ ;
wire _5079_ ;
wire _6860_ ;
wire _6440_ ;
wire _6020_ ;
wire \datapath.idinstr_15_bF$buf18  ;
wire \datapath.idinstr_15_hier0_bF$buf6  ;
wire \datapath.idinstr_22_bF$buf22  ;
wire _7645_ ;
wire _7225_ ;
wire _2780_ ;
wire _2360_ ;
wire _3985_ ;
wire _3565_ ;
wire _3145_ ;
wire _5711_ ;
wire _8183_ ;
wire \datapath.idinstr_16_bF$buf27  ;
wire _49_ ;
wire _6916_ ;
wire _1631_ ;
wire _1211_ ;
wire _9388_ ;
wire \datapath.idinstr_20_bF$buf42  ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _2836_ ;
wire \datapath.idinstr_15_bF$buf5  ;
wire _2416_ ;
wire _7874_ ;
wire _7454_ ;
wire _7034_ ;
wire _8659_ ;
wire _8239_ ;
wire _3794_ ;
wire _3374_ ;
wire \datapath.idinstr_17_bF$buf36  ;
wire _4999_ ;
wire _4579_ ;
wire _4159_ ;
wire _5940_ ;
wire _5520_ ;
wire _5100_ ;
wire _6725_ ;
wire _6305_ ;
wire _1860_ ;
wire _1440_ ;
wire _1020_ ;
wire _9197_ ;
wire _771_ ;
wire _351_ ;
wire _2645_ ;
wire _2225_ ;
wire _7683_ ;
wire _7263_ ;
wire _8888_ ;
wire _8468_ ;
wire _8048_ ;
wire _3183_ ;
wire _1916_ ;
wire _4388_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _6954_ ;
wire _6534_ ;
wire _6114_ ;
wire _580_ ;
wire _160_ ;
wire _7739_ ;
wire _7319_ ;
wire _2874_ ;
wire _2454_ ;
wire _2034_ ;
wire _3659_ ;
wire _3239_ ;
wire _4600_ ;
wire _7492_ ;
wire _7072_ ;
wire _5805_ ;
wire _8697_ ;
wire _8277_ ;
wire _1725_ ;
wire _1305_ ;
wire _4197_ ;
wire _636_ ;
wire _216_ ;
wire _6763_ ;
wire _6343_ ;
wire _7968_ ;
wire _7548_ ;
wire _7128_ ;
wire \datapath.idinstr_24_bF$buf1  ;
wire _2683_ ;
wire _2263_ ;
wire _3888_ ;
wire _3468_ ;
wire _3048_ ;
wire _5614_ ;
wire _8086_ ;
wire [31:0] \datapath.csr._13_  ;
wire \datapath.pcstall_bF$buf7  ;
wire \datapath.alu.b_2_bF$buf0  ;
wire _6819_ ;
wire _1954_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire _2739_ ;
wire _2319_ ;
wire _6992_ ;
wire _6572_ ;
wire _6152_ ;
wire _7777_ ;
wire _7357_ ;
wire _2492_ ;
wire _2072_ ;
wire \datapath.idinstr_22_bF$buf8  ;
wire _3697_ ;
wire _3277_ ;
wire _5843_ ;
wire _5423_ ;
wire _5003_ ;
wire _6628_ ;
wire _6208_ ;
wire _1763_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _2968_ ;
wire _2548_ ;
wire _2128_ ;
wire _6381_ ;
wire _7586_ ;
wire _7166_ ;
wire _3086_ ;
wire _9312_ ;
wire _1819_ ;
wire _5652_ ;
wire _5232_ ;
wire _6857_ ;
wire _6437_ ;
wire _6017_ ;
wire _1992_ ;
wire _1572_ ;
wire _1152_ ;
wire _483_ ;
wire \datapath.idinstr_22_bF$buf19  ;
wire _2777_ ;
wire _2357_ ;
wire _6190_ ;
wire _4923_ ;
wire _4503_ ;
wire _7395_ ;
wire _5708_ ;
wire _9121_ ;
wire _1628_ ;
wire _1208_ ;
wire _5881_ ;
wire _5461_ ;
wire _5041_ ;
wire \datapath.idinstr_20_bF$buf39  ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _6666_ ;
wire _6246_ ;
wire _1381_ ;
wire _292_ ;
wire _2586_ ;
wire _2166_ ;
wire _8812_ ;
wire _4732_ ;
wire _4312_ ;
wire _5937_ ;
wire _5517_ ;
wire _11_ ;
wire _9350_ ;
wire \datapath.alu.b_0_bF$buf9  ;
wire _1857_ ;
wire _1437_ ;
wire _1017_ ;
wire _5690_ ;
wire _5270_ ;
wire _768_ ;
wire _348_ ;
wire _6895_ ;
wire _6475_ ;
wire _6055_ ;
wire _1190_ ;
wire _2395_ ;
wire _8621_ ;
wire _8201_ ;
wire _9406_ ;
wire _4961_ ;
wire _4541_ ;
wire _4121_ ;
wire [1:0] \datapath.csr.mstatus  ;
wire _5746_ ;
wire _5326_ ;
wire _6145__bF$buf0 ;
wire _6145__bF$buf1 ;
wire _6145__bF$buf2 ;
wire _6145__bF$buf3 ;
wire _6145__bF$buf4 ;
wire _6145__bF$buf5 ;
wire \controlunit.ill_op  ;
wire _6145__bF$buf6 ;
wire _6145__bF$buf7 ;
wire _5458__bF$buf0 ;
wire _5458__bF$buf1 ;
wire _5458__bF$buf2 ;
wire _5458__bF$buf3 ;
wire _5458__bF$buf4 ;
wire _1666_ ;
wire _1246_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _3812_ ;
wire _6284_ ;
wire _7489_ ;
wire _7069_ ;
wire _8850_ ;
wire _8430_ ;
wire _8010_ ;
wire _9215_ ;
wire _4770_ ;
wire _4350_ ;
wire \datapath.idinstr_21_hier0_bF$buf4  ;
wire _5975_ ;
wire _5555_ ;
wire _5135_ ;
wire _5462__bF$buf0 ;
wire _5462__bF$buf1 ;
wire _5462__bF$buf2 ;
wire _5462__bF$buf3 ;
wire _5462__bF$buf4 ;
wire _1895_ ;
wire _1475_ ;
wire _1055_ ;
wire _7701_ ;
wire _386_ ;
wire _8906_ ;
wire _3621_ ;
wire _3201_ ;
wire _6093_ ;
wire _4826_ ;
wire _4406_ ;
wire _7298_ ;
wire _9024_ ;
wire _5784_ ;
wire _5364_ ;
wire _982__bF$buf0 ;
wire _982__bF$buf1 ;
wire _982__bF$buf2 ;
wire _982__bF$buf3 ;
wire _982__bF$buf4 ;
wire _6989_ ;
wire _6569_ ;
wire _6149_ ;
wire _1284_ ;
wire _7930_ ;
wire _7510_ ;
wire _195_ ;
wire _2489_ ;
wire _2069_ ;
wire _8715_ ;
wire _3850_ ;
wire _3430_ ;
wire _3010_ ;
wire _4635_ ;
wire _4215_ ;
wire _9253_ ;
wire _2701_ ;
wire _5593_ ;
wire _5173_ ;
wire _3906_ ;
wire _6798_ ;
wire _6378_ ;
wire _1093_ ;
wire _2298_ ;
wire _8944_ ;
wire _8524_ ;
wire _8104_ ;
wire _9309_ ;
wire _4864_ ;
wire _4444_ ;
wire _4024_ ;
wire _5649_ ;
wire _5229_ ;
wire _9062_ ;
wire _1989_ ;
wire _1569_ ;
wire _1149_ ;
wire _2930_ ;
wire _2510_ ;
wire _3715_ ;
wire _6187_ ;
wire _8753_ ;
wire _8333_ ;
wire _9118_ ;
wire _4673_ ;
wire _4253_ ;
wire _5878_ ;
wire _5458_ ;
wire _5038_ ;
wire _9291_ ;
wire _1798_ ;
wire _1378_ ;
wire _7604_ ;
wire _289_ ;
wire _8809_ ;
wire _3944_ ;
wire _3524_ ;
wire _3104_ ;
wire _5_ ;
wire _4729_ ;
wire _4309_ ;
wire _8982_ ;
wire _8562_ ;
wire _8142_ ;
wire _9347_ ;
wire _4482_ ;
wire _4062_ ;
wire _921_ ;
wire _501_ ;
wire _5687_ ;
wire _5267_ ;
wire _1187_ ;
wire _7833_ ;
wire _7413_ ;
wire _8618_ ;
wire _3753_ ;
wire _3333_ ;
wire _4958_ ;
wire _4538_ ;
wire \datapath.idinstr_21_bF$buf10  ;
wire _4118_ ;
wire _8791_ ;
wire _8371_ ;
wire _9156_ ;
wire _4291_ ;
wire _730_ ;
wire _310_ ;
wire _2604_ ;
wire _5496_ ;
wire _5076_ ;
wire CLK_bF$buf150 ;
wire CLK_bF$buf151 ;
wire CLK_bF$buf152 ;
wire CLK_bF$buf153 ;
wire \datapath.idinstr_15_bF$buf15  ;
wire _3809_ ;
wire \datapath.idinstr_15_hier0_bF$buf3  ;
wire _7642_ ;
wire _7222_ ;
wire _8847_ ;
wire _8427_ ;
wire _8007_ ;
wire _3982_ ;
wire _3562_ ;
wire _3142_ ;
wire _4767_ ;
wire _4347_ ;
wire _8180_ ;
wire \datapath.idinstr_16_bF$buf24  ;
wire _46_ ;
wire _6913_ ;
wire _9385_ ;
wire _2833_ ;
wire \datapath.idinstr_15_bF$buf2  ;
wire _2413_ ;
wire _3618_ ;
wire _7871_ ;
wire _7451_ ;
wire _7031_ ;
wire _8656_ ;
wire _8236_ ;
wire _3791_ ;
wire _3371_ ;
wire \datapath.idinstr_17_bF$buf33  ;
wire \datapath.regmret  ;
wire _4996_ ;
wire _4576_ ;
wire _4156_ ;
wire _6722_ ;
wire _6302_ ;
wire _9194_ ;
wire _7927_ ;
wire _7507_ ;
wire _2642_ ;
wire _2222_ ;
wire \datapath.idinstr_15_bF$buf53  ;
wire _3847_ ;
wire _3427_ ;
wire _3007_ ;
wire _7680_ ;
wire _7260_ ;
wire _8885_ ;
wire _8465_ ;
wire _8045_ ;
wire _3180_ ;
wire _1913_ ;
wire _4385_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _6951_ ;
wire _6531_ ;
wire _6111_ ;
wire _7736_ ;
wire _7316_ ;
wire _2871_ ;
wire _2451_ ;
wire _2031_ ;
wire [31:0] \datapath.registers.1226[15]  ;
wire _3656_ ;
wire _3236_ ;
wire _5802_ ;
wire _8694_ ;
wire _8274_ ;
wire _1722_ ;
wire _1302_ ;
wire _9059_ ;
wire _4194_ ;
wire _633_ ;
wire _213_ ;
wire _2927_ ;
wire _2507_ ;
wire _5399_ ;
wire _6760_ ;
wire _6340_ ;
wire _7965_ ;
wire _7545_ ;
wire _7125_ ;
wire _2680_ ;
wire _2260_ ;
wire \datapath.idinstr_18_bF$buf5  ;
wire _3885_ ;
wire _3465_ ;
wire _3045_ ;
wire _5611_ ;
wire _8083_ ;
wire \datapath.pcstall_bF$buf4  ;
wire _6816_ ;
wire _1951_ ;
wire _1531_ ;
wire _1111_ ;
wire _9288_ ;
wire _862_ ;
wire _442_ ;
wire _2736_ ;
wire _2316_ ;
wire _7774_ ;
wire _7354_ ;
wire \datapath.idinstr_22_bF$buf5  ;
wire _8979_ ;
wire _8559_ ;
wire _8139_ ;
wire _3694_ ;
wire _3274_ ;
wire _4899_ ;
wire _4479_ ;
wire _4059_ ;
wire _5840_ ;
wire _5420_ ;
wire _5000_ ;
wire _918_ ;
wire _6625_ ;
wire _6205_ ;
wire _1760_ ;
wire _1340_ ;
wire _9097_ ;
wire _671_ ;
wire _251_ ;
wire _2965_ ;
wire _2545_ ;
wire _2125_ ;
wire _7583_ ;
wire _7163_ ;
wire _8788_ ;
wire _8368_ ;
wire _3083_ ;
wire _1816_ ;
wire _4288_ ;
wire _727_ ;
wire _307_ ;
wire _6854_ ;
wire _6434_ ;
wire _6014_ ;
wire _480_ ;
wire \datapath.idinstr_22_bF$buf16  ;
wire _7639_ ;
wire _7219_ ;
wire _2774_ ;
wire _2354_ ;
wire _3979_ ;
wire _3559_ ;
wire _3139_ ;
wire _4920_ ;
wire _4500_ ;
wire _7392_ ;
wire _5705_ ;
wire _8597_ ;
wire _8177_ ;
wire _1625_ ;
wire _1205_ ;
wire _4097_ ;
wire \datapath.idinstr_20_bF$buf36  ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _6663_ ;
wire _6243_ ;
wire _7868_ ;
wire _7448_ ;
wire _7028_ ;
wire _2583_ ;
wire _2163_ ;
wire _3788_ ;
wire _3368_ ;
wire _5934_ ;
wire _5514_ ;
wire _6719_ ;
wire \datapath.alu.b_0_bF$buf6  ;
wire _1854_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _2639_ ;
wire _2219_ ;
wire _6892_ ;
wire _6472_ ;
wire _6052_ ;
wire _7677_ ;
wire _7257_ ;
wire _2392_ ;
wire _3597_ ;
wire _3177_ ;
wire _9403_ ;
wire _5743_ ;
wire _5323_ ;
wire _6948_ ;
wire _6528_ ;
wire _6108_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _2868_ ;
wire _2448_ ;
wire _2028_ ;
wire _6281_ ;
wire _7486_ ;
wire _7066_ ;
wire _5993__bF$buf0 ;
wire _5993__bF$buf1 ;
wire _5993__bF$buf2 ;
wire _5993__bF$buf3 ;
wire _5993__bF$buf4 ;
wire _5993__bF$buf5 ;
wire _5993__bF$buf6 ;
wire _5993__bF$buf7 ;
wire _9212_ ;
wire _1719_ ;
wire \datapath.idinstr_21_hier0_bF$buf1  ;
wire _5972_ ;
wire _5552_ ;
wire _5132_ ;
wire _6757_ ;
wire _6337_ ;
wire _1892_ ;
wire _1472_ ;
wire _1052_ ;
wire _383_ ;
wire _2677_ ;
wire _2257_ ;
wire _8903_ ;
wire _6090_ ;
wire \controlunit.regfile_wen  ;
wire _4823_ ;
wire _4403_ ;
wire _7295_ ;
wire _5608_ ;
wire \datapath.pcstall  ;
wire _9441_ ;
wire _9021_ ;
wire _1948_ ;
wire _1528_ ;
wire _1108_ ;
wire _5781_ ;
wire _5361_ ;
wire _859_ ;
wire _439_ ;
wire _6986_ ;
wire _6566_ ;
wire _6146_ ;
wire _1281_ ;
wire _192_ ;
wire _2486_ ;
wire _2066_ ;
wire _8712_ ;
wire _4632_ ;
wire _4212_ ;
wire _5837_ ;
wire _5417_ ;
wire _9250_ ;
wire _1757_ ;
wire _1337_ ;
wire _5590_ ;
wire _5170_ ;
wire _668_ ;
wire [31:0] _248_ ;
wire _3903_ ;
wire _6795_ ;
wire _6375_ ;
wire _1090_ ;
wire _2295_ ;
wire _8941_ ;
wire _8521_ ;
wire _8101_ ;
wire _9306_ ;
wire _4861_ ;
wire _4441_ ;
wire _4021_ ;
wire _5646_ ;
wire _5226_ ;
wire _1986_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _3712_ ;
wire _6184_ ;
wire _4917_ ;
wire _7389_ ;
wire _8750_ ;
wire _8330_ ;
wire _9115_ ;
wire _4670_ ;
wire _4250_ ;
wire _5875_ ;
wire _5455_ ;
wire _5035_ ;
wire _1795_ ;
wire _1375_ ;
wire _7601_ ;
wire _286_ ;
wire [31:0] \datapath.csr.mcause  ;
wire _8806_ ;
wire _3941_ ;
wire _3521_ ;
wire _3101_ ;
wire _2_ ;
wire _4726_ ;
wire _4306_ ;
wire _7198_ ;
wire _9344_ ;
wire _5684_ ;
wire _5264_ ;
wire _6889_ ;
wire _6469_ ;
wire _6049_ ;
wire _1184_ ;
wire _7830_ ;
wire _7410_ ;
wire _2389_ ;
wire _8615_ ;
wire _3750_ ;
wire _3330_ ;
wire _4955_ ;
wire _4535_ ;
wire _4115_ ;
wire _9153_ ;
wire _2601_ ;
wire _5493_ ;
wire _5073_ ;
wire CLK_bF$buf120 ;
wire CLK_bF$buf121 ;
wire [31:0] \datapath.registers.1226[30]  ;
wire CLK_bF$buf122 ;
wire CLK_bF$buf123 ;
wire CLK_bF$buf124 ;
wire CLK_bF$buf125 ;
wire \datapath.idinstr_15_bF$buf12  ;
wire CLK_bF$buf126 ;
wire CLK_bF$buf127 ;
wire CLK_bF$buf128 ;
wire _3806_ ;
wire CLK_bF$buf129 ;
wire \datapath.idinstr_15_hier0_bF$buf0  ;
wire _6698_ ;
wire _6278_ ;
wire _2198_ ;
wire _8844_ ;
wire _8424_ ;
wire _8004_ ;
wire _7608__bF$buf0 ;
wire _7608__bF$buf1 ;
wire _7608__bF$buf2 ;
wire _7608__bF$buf3 ;
wire _7608__bF$buf4 ;
wire _7608__bF$buf5 ;
wire _7608__bF$buf6 ;
wire _7608__bF$buf7 ;
wire _7608__bF$buf8 ;
wire _7608__bF$buf9 ;
wire _9209_ ;
wire _4764_ ;
wire _4344_ ;
wire _5969_ ;
wire _5549_ ;
wire _5129_ ;
wire \datapath.idinstr_16_bF$buf21  ;
wire _43_ ;
wire _6910_ ;
wire _9382_ ;
wire _1889_ ;
wire _1469_ ;
wire _1049_ ;
wire _2830_ ;
wire _2410_ ;
wire _3615_ ;
wire _6087_ ;
wire _8653_ ;
wire _8233_ ;
wire \datapath.idinstr_17_bF$buf30  ;
wire _7612__bF$buf0 ;
wire _7612__bF$buf1 ;
wire _7612__bF$buf2 ;
wire _7612__bF$buf3 ;
wire _7612__bF$buf4 ;
wire _7612__bF$buf5 ;
wire _7612__bF$buf6 ;
wire _7612__bF$buf7 ;
wire _9438_ ;
wire _9018_ ;
wire _4993_ ;
wire _4573_ ;
wire _4153_ ;
wire _5778_ ;
wire _5358_ ;
wire _9191_ ;
wire _1698_ ;
wire _1278_ ;
wire _7924_ ;
wire _7504_ ;
wire _189_ ;
wire _8709_ ;
wire \datapath.idinstr_15_bF$buf50  ;
wire _3844_ ;
wire _3424_ ;
wire _3004_ ;
wire _4629_ ;
wire _4209_ ;
wire _8882_ ;
wire _8462_ ;
wire _8042_ ;
wire \datapath.idinstr_16_hier0_bF$buf5  ;
wire _1910_ ;
wire _9247_ ;
wire _4382_ ;
wire _821_ ;
wire _401_ ;
wire _5587_ ;
wire _5167_ ;
wire _81_ ;
wire _1087_ ;
wire _7733_ ;
wire _7313_ ;
wire _8938_ ;
wire _8518_ ;
wire _3653_ ;
wire _3233_ ;
wire _4858_ ;
wire _4438_ ;
wire _4018_ ;
wire _8691_ ;
wire _8271_ ;
wire _9056_ ;
wire _4191_ ;
wire _630_ ;
wire _210_ ;
wire _2924_ ;
wire _2504_ ;
wire _5396_ ;
wire _3709_ ;
wire _7962_ ;
wire _7542_ ;
wire _7122_ ;
wire \datapath.idinstr_18_bF$buf2  ;
wire _8747_ ;
wire _8327_ ;
wire _3882_ ;
wire _3462_ ;
wire _3042_ ;
wire [31:0] \datapath.regcsrwb  ;
wire _4667_ ;
wire _4247_ ;
wire _8080_ ;
wire \datapath.pcstall_bF$buf1  ;
wire _6813_ ;
wire _9285_ ;
wire _2733_ ;
wire _2313_ ;
wire _5484__bF$buf0 ;
wire _5484__bF$buf1 ;
wire _5484__bF$buf2 ;
wire _5484__bF$buf3 ;
wire _5484__bF$buf4 ;
wire _3938_ ;
wire _3518_ ;
wire _7771_ ;
wire _7351_ ;
wire \datapath.idinstr_22_bF$buf2  ;
wire \datapath.idinstr_16_bF$buf9  ;
wire _8976_ ;
wire _8556_ ;
wire _8136_ ;
wire _3691_ ;
wire _3271_ ;
wire _4896_ ;
wire _4476_ ;
wire _4056_ ;
wire _915_ ;
wire _6622_ ;
wire _6202_ ;
wire _9094_ ;
wire _7827_ ;
wire _7407_ ;
wire _2962_ ;
wire _2542_ ;
wire _2122_ ;
wire _3747_ ;
wire _3327_ ;
wire _7580_ ;
wire _7160_ ;
wire \datapath.idinstr_20_bF$buf9  ;
wire _8785_ ;
wire _8365_ ;
wire _3080_ ;
wire _1813_ ;
wire _4285_ ;
wire _724_ ;
wire _304_ ;
wire _6851_ ;
wire _6431_ ;
wire _6011_ ;
wire [31:0] \datapath.bbypass  ;
wire \datapath.idinstr_22_bF$buf13  ;
wire _7636_ ;
wire _7216_ ;
wire _2771_ ;
wire _2351_ ;
wire _3976_ ;
wire _3556_ ;
wire _3136_ ;
wire _5702_ ;
wire _8594_ ;
wire _8174_ ;
wire \datapath.idinstr_16_bF$buf18  ;
wire _6907_ ;
wire _1622_ ;
wire _1202_ ;
wire _9379_ ;
wire _4094_ ;
wire \datapath.idinstr_20_bF$buf33  ;
wire _953_ ;
wire _533_ ;
wire _113_ ;
wire _2827_ ;
wire _2407_ ;
wire _5299_ ;
wire _6660_ ;
wire _6240_ ;
wire _7865_ ;
wire _7445_ ;
wire _7025_ ;
wire _2580_ ;
wire _2160_ ;
wire _3785_ ;
wire _3365_ ;
wire \datapath.idinstr_17_bF$buf27  ;
wire \datapath.idinstr_21_bF$buf42  ;
wire _5931_ ;
wire _5511_ ;
wire _6716_ ;
wire \datapath.alu.b_0_bF$buf3  ;
wire _1851_ ;
wire _1431_ ;
wire _1011_ ;
wire _9188_ ;
wire _762_ ;
wire _342_ ;
wire _2636_ ;
wire _2216_ ;
wire \datapath.idinstr_15_bF$buf47  ;
wire _7674_ ;
wire _7254_ ;
wire [31:0] \datapath.registers.1226[6]  ;
wire _8879_ ;
wire _8459_ ;
wire _8039_ ;
wire _3594_ ;
wire _3174_ ;
wire _9400_ ;
wire _1907_ ;
wire _4799_ ;
wire _4379_ ;
wire _5740_ ;
wire _5320_ ;
wire _818_ ;
wire _78_ ;
wire _6945_ ;
wire _6525_ ;
wire _6105_ ;
wire _1660_ ;
wire _1240_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _2865_ ;
wire _2445_ ;
wire _2025_ ;
wire _7483_ ;
wire _7063_ ;
wire _6140__bF$buf0 ;
wire _6140__bF$buf1 ;
wire _6140__bF$buf2 ;
wire _6140__bF$buf3 ;
wire _6140__bF$buf4 ;
wire _8688_ ;
wire _8268_ ;
wire _7608__bF$buf10 ;
wire _1716_ ;
wire _4188_ ;
wire _627_ ;
wire _207_ ;
wire _6754_ ;
wire _6334_ ;
wire _380_ ;
wire _7959_ ;
wire _7539_ ;
wire _7119_ ;
wire _2674_ ;
wire _2254_ ;
wire _8900_ ;
wire _3879_ ;
wire _3459_ ;
wire _3039_ ;
wire _4820_ ;
wire _4400_ ;
wire _7292_ ;
wire _5605_ ;
wire _8497_ ;
wire _8077_ ;
wire \datapath.regcsrtrap_bF$buf7  ;
wire _1945_ ;
wire _1525_ ;
wire _1105_ ;
wire _856_ ;
wire _436_ ;
wire _6983_ ;
wire _6563_ ;
wire _6143_ ;
wire \datapath.alu.b_3_bF$buf6  ;
wire _7768_ ;
wire _7348_ ;
wire _2483_ ;
wire _2063_ ;
wire _3688_ ;
wire _3268_ ;
wire _5834_ ;
wire _5414_ ;
wire _6619_ ;
wire _1754_ ;
wire _1334_ ;
wire _665_ ;
wire _245_ ;
wire _2959_ ;
wire _2539_ ;
wire _2119_ ;
wire [29:0] \datapath.csr.mepc  ;
wire _3900_ ;
wire _6792_ ;
wire _6372_ ;
wire _7997_ ;
wire _7577_ ;
wire _7157_ ;
wire _2292_ ;
wire _3497_ ;
wire _3077_ ;
wire _9303_ ;
wire _5643_ ;
wire _5223_ ;
wire _6848_ ;
wire _6428_ ;
wire _6008_ ;
wire _1983_ ;
wire _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _2768_ ;
wire _2348_ ;
wire _6181_ ;
wire _4914_ ;
wire _7386_ ;
wire _9112_ ;
wire _1619_ ;
wire _5872_ ;
wire _5452_ ;
wire _5032_ ;
wire _6657_ ;
wire _6237_ ;
wire _1792_ ;
wire _1372_ ;
wire CLK_hier0_bF$buf0 ;
wire CLK_hier0_bF$buf1 ;
wire CLK_hier0_bF$buf2 ;
wire CLK_hier0_bF$buf3 ;
wire CLK_hier0_bF$buf4 ;
wire CLK_hier0_bF$buf5 ;
wire CLK_hier0_bF$buf6 ;
wire CLK_hier0_bF$buf7 ;
wire CLK_hier0_bF$buf8 ;
wire CLK_hier0_bF$buf9 ;
wire _283_ ;
wire _2997_ ;
wire _2577_ ;
wire _2157_ ;
wire _8803_ ;
wire _4723_ ;
wire _4303_ ;
wire _7195_ ;
wire _9175__bF$buf0 ;
wire _9175__bF$buf1 ;
wire _9175__bF$buf2 ;
wire _9175__bF$buf3 ;
wire _9175__bF$buf4 ;
wire _9175__bF$buf5 ;
wire _9175__bF$buf6 ;
wire _9175__bF$buf7 ;
wire \datapath.idinstr_21_bF$buf39  ;
wire _5928_ ;
wire _5508_ ;
wire _9341_ ;
wire _1848_ ;
wire _1428_ ;
wire _1008_ ;
wire _5681_ ;
wire _5261_ ;
wire _759_ ;
wire _339_ ;
wire _6886_ ;
wire _6466_ ;
wire _6046_ ;
wire _1181_ ;
wire \datapath.idinstr_22_hier0_bF$buf5  ;
wire _2386_ ;
wire _8612_ ;
wire _4952_ ;
wire _4532_ ;
wire _4112_ ;
wire _5737_ ;
wire _5317_ ;
wire _9150_ ;
wire _1657_ ;
wire _1237_ ;
wire _5490_ ;
wire _5070_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _3803_ ;
wire _6695_ ;
wire _6275_ ;
wire _2195_ ;
wire _8841_ ;
wire _8421_ ;
wire _8001_ ;
wire _5614__bF$buf0 ;
wire _5614__bF$buf1 ;
wire _5614__bF$buf2 ;
wire _5614__bF$buf3 ;
wire _5614__bF$buf4 ;
wire _5468__bF$buf0 ;
wire _5468__bF$buf1 ;
wire _5468__bF$buf2 ;
wire _9206_ ;
wire _5468__bF$buf3 ;
wire _5468__bF$buf4 ;
wire _4761_ ;
wire _4341_ ;
wire _5966_ ;
wire _5546_ ;
wire _5126_ ;
wire _495__bF$buf0 ;
wire _495__bF$buf1 ;
wire _495__bF$buf2 ;
wire _495__bF$buf3 ;
wire _40_ ;
wire _495__bF$buf4 ;
wire _1886_ ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire _3612_ ;
wire _6084_ ;
wire _4817_ ;
wire _7289_ ;
wire _8650_ ;
wire _8230_ ;
wire _5472__bF$buf0 ;
wire _5472__bF$buf1 ;
wire _5472__bF$buf2 ;
wire _5472__bF$buf3 ;
wire _5472__bF$buf4 ;
wire _9435_ ;
wire _9015_ ;
wire _4990_ ;
wire _4570_ ;
wire _4150_ ;
wire _5775_ ;
wire _5355_ ;
wire _1695_ ;
wire _1275_ ;
wire _7921_ ;
wire _7501_ ;
wire _186_ ;
wire _8706_ ;
wire _3841_ ;
wire _3421_ ;
wire _3001_ ;
wire _4626_ ;
wire _4206_ ;
wire _7098_ ;
wire \datapath.idinstr_16_hier0_bF$buf2  ;
wire _9244_ ;
wire _5584_ ;
wire _5164_ ;
wire _6789_ ;
wire _6369_ ;
wire _1084_ ;
wire _7730_ ;
wire _7310_ ;
wire _2289_ ;
wire _8935_ ;
wire _8515_ ;
wire _3650_ ;
wire _3230_ ;
wire _4855_ ;
wire _4435_ ;
wire _4015_ ;
wire _9053_ ;
wire _2921_ ;
wire _2501_ ;
wire _5393_ ;
wire [31:0] \datapath.registers.1226[20]  ;
wire _3706_ ;
wire _6598_ ;
wire _6178_ ;
wire _2098_ ;
wire _8744_ ;
wire _8324_ ;
wire _9109_ ;
wire _4664_ ;
wire _4244_ ;
wire _5869_ ;
wire _5449_ ;
wire _5029_ ;
wire _6810_ ;
wire _9282_ ;
wire _1789_ ;
wire _1369_ ;
wire _2730_ ;
wire _2310_ ;
wire _3935_ ;
wire _3515_ ;
wire \datapath.idinstr_16_bF$buf6  ;
wire _8973_ ;
wire _8553_ ;
wire _8133_ ;
wire _9338_ ;
wire _4893_ ;
wire _4473_ ;
wire _4053_ ;
wire _912_ ;
wire _5678_ ;
wire _5258_ ;
wire _9091_ ;
wire _1598_ ;
wire _1178_ ;
wire _7824_ ;
wire _7404_ ;
wire _8609_ ;
wire _3744_ ;
wire _3324_ ;
wire _4949_ ;
wire \datapath.idinstr_20_bF$buf6  ;
wire _4529_ ;
wire _4109_ ;
wire _8782_ ;
wire _8362_ ;
wire _1810_ ;
wire _9147_ ;
wire _4282_ ;
wire _721_ ;
wire _301_ ;
wire _5487_ ;
wire _5067_ ;
wire \datapath.idinstr_22_bF$buf10  ;
wire _7633_ ;
wire _7213_ ;
wire _8838_ ;
wire _8418_ ;
wire _3973_ ;
wire _3553_ ;
wire _3133_ ;
wire _4758_ ;
wire _4338_ ;
wire _8591_ ;
wire _8171_ ;
wire \datapath.idinstr_16_bF$buf15  ;
wire _37_ ;
wire _6904_ ;
wire _9376_ ;
wire _4091_ ;
wire \datapath.idinstr_20_bF$buf30  ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _2824_ ;
wire _2404_ ;
wire _5296_ ;
wire _3609_ ;
wire _7862_ ;
wire _7442_ ;
wire _7022_ ;
wire _8647_ ;
wire _8227_ ;
wire _3782_ ;
wire _3362_ ;
wire \datapath.idinstr_17_bF$buf24  ;
wire _4987_ ;
wire _4567_ ;
wire _4147_ ;
wire _6713_ ;
wire \datapath.alu.b_0_bF$buf0  ;
wire _9185_ ;
wire _7918_ ;
wire _2633_ ;
wire _2213_ ;
wire \datapath.idinstr_15_bF$buf44  ;
wire _3838_ ;
wire _3418_ ;
wire _7671_ ;
wire _7251_ ;
wire _8876_ ;
wire _8456_ ;
wire _8036_ ;
wire _3591_ ;
wire _3171_ ;
wire _1904_ ;
wire _4796_ ;
wire _4376_ ;
wire _815_ ;
wire _75_ ;
wire _6942_ ;
wire _6522_ ;
wire _6102_ ;
wire _7727_ ;
wire _7307_ ;
wire _2862_ ;
wire _2442_ ;
wire _2022_ ;
wire _3647_ ;
wire _3227_ ;
wire _7480_ ;
wire _7060_ ;
wire _8685_ ;
wire _8265_ ;
wire _1713_ ;
wire _4185_ ;
wire _624_ ;
wire _204_ ;
wire _2918_ ;
wire _6751_ ;
wire _6331_ ;
wire _7956_ ;
wire _7536_ ;
wire _7116_ ;
wire _2671_ ;
wire _2251_ ;
wire _3876_ ;
wire _3456_ ;
wire _3036_ ;
wire _5602_ ;
wire _8494_ ;
wire _8074_ ;
wire \datapath.regcsrtrap_bF$buf4  ;
wire _6807_ ;
wire _1942_ ;
wire _1522_ ;
wire _1102_ ;
wire _9279_ ;
wire _853_ ;
wire _433_ ;
wire _2727_ ;
wire _2307_ ;
wire _5199_ ;
wire _6980_ ;
wire _6560_ ;
wire _6140_ ;
wire \datapath.alu.b_3_bF$buf3  ;
wire _7765_ ;
wire _7345_ ;
wire _2480_ ;
wire _2060_ ;
wire [31:0] \datapath.programcounter.pc  ;
wire _3685_ ;
wire _3265_ ;
wire _5831_ ;
wire _5411_ ;
wire _909_ ;
wire _6616_ ;
wire _1751_ ;
wire _1331_ ;
wire _9088_ ;
wire _662_ ;
wire _242_ ;
wire _2956_ ;
wire _2536_ ;
wire _2116_ ;
wire _7994_ ;
wire _7574_ ;
wire _7154_ ;
wire _8779_ ;
wire _8359_ ;
wire _3494_ ;
wire _3074_ ;
wire _9300_ ;
wire _1807_ ;
wire _4699_ ;
wire _4279_ ;
wire _5640_ ;
wire _5220_ ;
wire _718_ ;
wire _6143__bF$buf0 ;
wire _6143__bF$buf1 ;
wire _6143__bF$buf2 ;
wire _6143__bF$buf3 ;
wire _6143__bF$buf4 ;
wire _6845_ ;
wire _6425_ ;
wire _6005_ ;
wire _1980_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _2765_ ;
wire _2345_ ;
wire _4911_ ;
wire _7383_ ;
wire _8588_ ;
wire _8168_ ;
wire _1616_ ;
wire _4088_ ;
wire \datapath.idinstr_20_bF$buf27  ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _6654_ ;
wire _6234_ ;
wire _280_ ;
wire _7859_ ;
wire _7439_ ;
wire _7019_ ;
wire _2994_ ;
wire _2574_ ;
wire _2154_ ;
wire _8800_ ;
wire _3779_ ;
wire _3359_ ;
wire _4720_ ;
wire _4300_ ;
wire _7192_ ;
wire \datapath.idinstr_21_bF$buf36  ;
wire _5925_ ;
wire _5505_ ;
wire _8397_ ;
wire _1845_ ;
wire _1425_ ;
wire _1005_ ;
wire _756_ ;
wire _336_ ;
wire _6883_ ;
wire _6463_ ;
wire _6043_ ;
wire \datapath.idinstr_22_hier0_bF$buf2  ;
wire _7668_ ;
wire _7248_ ;
wire _2383_ ;
wire _3588_ ;
wire _3168_ ;
wire _5734_ ;
wire _5314_ ;
wire _6939_ ;
wire _6519_ ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _2859_ ;
wire _2439_ ;
wire _2019_ ;
wire _3800_ ;
wire _6692_ ;
wire _6272_ ;
wire _7897_ ;
wire _7477_ ;
wire _7057_ ;
wire _2192_ ;
wire _3397_ ;
wire _9203_ ;
wire _5963_ ;
wire _5543_ ;
wire _5123_ ;
wire _6748_ ;
wire _6328_ ;
wire _1883_ ;
wire _1463_ ;
wire _1043_ ;
wire _794_ ;
wire _374_ ;
wire _2668_ ;
wire _2248_ ;
wire _6081_ ;
wire _4814_ ;
wire _7286_ ;
wire _9432_ ;
wire _9012_ ;
wire _1939_ ;
wire _1519_ ;
wire _5772_ ;
wire _5352_ ;
wire _6977_ ;
wire _6557_ ;
wire _6137_ ;
wire _1692_ ;
wire _1272_ ;
wire _183_ ;
wire _2897_ ;
wire _2477_ ;
wire _2057_ ;
wire _8703_ ;
wire _4623_ ;
wire _4203_ ;
wire _7095_ ;
wire _5828_ ;
wire _5408_ ;
wire _9241_ ;
wire _1748_ ;
wire _1328_ ;
wire _5581_ ;
wire _5161_ ;
wire _659_ ;
wire _239_ ;
wire [31:0] \datapath.memoryinterface.data_store  ;
wire _6786_ ;
wire _6366_ ;
wire _1081_ ;
wire _2286_ ;
wire _8932_ ;
wire _8512_ ;
wire _4852_ ;
wire _4432_ ;
wire _4012_ ;
wire _5637_ ;
wire _5217_ ;
wire \datapath.regcsrtrap  ;
wire _9050_ ;
wire _1977_ ;
wire _1557_ ;
wire _1137_ ;
wire _5390_ ;
wire _888_ ;
wire _468_ ;
wire _3703_ ;
wire _6595_ ;
wire _6175_ ;
wire _4908_ ;
wire _2095_ ;
wire _8741_ ;
wire _8321_ ;
wire _9106_ ;
wire _4661_ ;
wire _4241_ ;
wire _5866_ ;
wire _5446_ ;
wire _5026_ ;
wire _1786_ ;
wire _1366_ ;
wire _5715__bF$buf0 ;
wire _5715__bF$buf1 ;
wire _5715__bF$buf2 ;
wire _5715__bF$buf3 ;
wire _5715__bF$buf4 ;
wire _5715__bF$buf5 ;
wire _5715__bF$buf6 ;
wire _5715__bF$buf7 ;
wire _697_ ;
wire _277_ ;
wire _3932_ ;
wire _3512_ ;
wire _4717_ ;
wire _7189_ ;
wire \datapath.idinstr_16_bF$buf3  ;
wire _8970_ ;
wire _8550_ ;
wire _8130_ ;
wire _9335_ ;
wire _4890_ ;
wire _4470_ ;
wire _4050_ ;
wire _0__0_bF$buf0 ;
wire _5675_ ;
wire _0__0_bF$buf1 ;
wire _5255_ ;
wire _0__0_bF$buf2 ;
wire _0__0_bF$buf3 ;
wire _0__0_bF$buf4 ;
wire _1595_ ;
wire _1175_ ;
wire _7821_ ;
wire _7401_ ;
wire _8606_ ;
wire _3741_ ;
wire _3321_ ;
wire _4946_ ;
wire \datapath.idinstr_20_bF$buf3  ;
wire _4526_ ;
wire _4106_ ;
wire _9144_ ;
wire \datapath.allowcsrwrite  ;
wire _5484_ ;
wire _5064_ ;
wire _6689_ ;
wire _6269_ ;
wire _7630_ ;
wire _7210_ ;
wire _2189_ ;
wire _8835_ ;
wire _8415_ ;
wire _3970_ ;
wire _3550_ ;
wire _3130_ ;
wire _4755_ ;
wire _4335_ ;
wire \datapath.idinstr_16_bF$buf12  ;
wire _34_ ;
wire _6901_ ;
wire _9373_ ;
wire _2821_ ;
wire _2401_ ;
wire _5293_ ;
wire [3:0] \datapath.csr.csr_mcause  ;
wire [31:0] \datapath.registers.1226[10]  ;
wire _3606_ ;
wire _6498_ ;
wire _6078_ ;
wire _8644_ ;
wire _8224_ ;
wire \datapath.idinstr_17_bF$buf21  ;
wire _9429_ ;
wire _9009_ ;
wire _4984_ ;
wire _4564_ ;
wire _4144_ ;
wire _5769_ ;
wire _5349_ ;
wire _6710_ ;
wire _9182_ ;
wire _1689_ ;
wire _1269_ ;
wire _7915_ ;
wire _2630_ ;
wire _2210_ ;
wire \datapath.idinstr_15_bF$buf41  ;
wire _3835_ ;
wire _3415_ ;
wire _8873_ ;
wire _8453_ ;
wire _8033_ ;
wire _1901_ ;
wire _9238_ ;
wire _4793_ ;
wire _4373_ ;
wire \datapath.idinstr_23_bF$buf6  ;
wire _812_ ;
wire _5998_ ;
wire _5578_ ;
wire _5158_ ;
wire _72_ ;
wire _1498_ ;
wire _1078_ ;
wire _7724_ ;
wire _7304_ ;
wire _8929_ ;
wire _8509_ ;
wire _3644_ ;
wire _3224_ ;
wire _4849_ ;
wire _4429_ ;
wire _4009_ ;
wire _8682_ ;
wire _8262_ ;
wire _1710_ ;
wire _9047_ ;
wire _4182_ ;
wire _621_ ;
wire _201_ ;
wire _2915_ ;
wire _5387_ ;
wire _7953_ ;
wire _7533_ ;
wire _7113_ ;
wire _8738_ ;
wire _8318_ ;
wire _3873_ ;
wire _3453_ ;
wire _3033_ ;
wire _4658_ ;
wire _4238_ ;
wire _8491_ ;
wire _8071_ ;
wire \datapath.regcsrtrap_bF$buf1  ;
wire _6804_ ;
wire _9276_ ;
wire _850_ ;
wire _430_ ;
wire _2724_ ;
wire _2304_ ;
wire _5196_ ;
wire _3929_ ;
wire _3509_ ;
wire \datapath.alu.b_3_bF$buf0  ;
wire _7762_ ;
wire _7342_ ;
wire _8967_ ;
wire _8547_ ;
wire _8127_ ;
wire _3682_ ;
wire _3262_ ;
wire _4887_ ;
wire _4467_ ;
wire _4047_ ;
wire _906_ ;
wire _5494__bF$buf0 ;
wire _5494__bF$buf1 ;
wire _5494__bF$buf2 ;
wire _5494__bF$buf3 ;
wire _5494__bF$buf4 ;
wire _6613_ ;
wire _9085_ ;
wire _7818_ ;
wire _2953_ ;
wire _2533_ ;
wire _2113_ ;
wire _3738_ ;
wire _3318_ ;
wire _7991_ ;
wire _7571_ ;
wire _7151_ ;
wire _8776_ ;
wire _8356_ ;
wire _3491_ ;
wire _3071_ ;
wire _1804_ ;
wire _4696_ ;
wire _4276_ ;
wire _715_ ;
wire _6842_ ;
wire _6422_ ;
wire _6002_ ;
wire _7627_ ;
wire _7207_ ;
wire _2762_ ;
wire _2342_ ;
wire _3967_ ;
wire _3547_ ;
wire _3127_ ;
wire _7380_ ;
wire _8585_ ;
wire _8165_ ;
wire _1613_ ;
wire _4085_ ;
wire \datapath.idinstr_20_bF$buf24  ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire _2818_ ;
wire _6651_ ;
wire _6231_ ;
wire _7856_ ;
wire _7436_ ;
wire _7016_ ;
wire _2991_ ;
wire _2571_ ;
wire _2151_ ;
wire _3800__bF$buf0 ;
wire [31:0] \datapath.registers.1226[27]  ;
wire _3800__bF$buf1 ;
wire _3800__bF$buf2 ;
wire _3800__bF$buf3 ;
wire _3800__bF$buf4 ;
wire _3800__bF$buf5 ;
wire _3800__bF$buf6 ;
wire _3800__bF$buf7 ;
wire _3776_ ;
wire _3356_ ;
wire \datapath.idinstr_17_bF$buf18  ;
wire \datapath.idinstr_21_bF$buf33  ;
wire _5922_ ;
wire _5502_ ;
wire _8394_ ;
wire _6707_ ;
wire _1842_ ;
wire _1422_ ;
wire _1002_ ;
wire _9179_ ;
wire _753_ ;
wire _333_ ;
wire _2627_ ;
wire _2207_ ;
wire _5099_ ;
wire _6880_ ;
wire _6460_ ;
wire _6040_ ;
wire _3339__bF$buf0 ;
wire _3339__bF$buf1 ;
wire _3339__bF$buf2 ;
wire _3339__bF$buf3 ;
wire _3339__bF$buf4 ;
wire _3339__bF$buf5 ;
wire \datapath.idinstr_15_bF$buf38  ;
wire _3339__bF$buf6 ;
wire \datapath.idinstr_22_bF$buf42  ;
wire _7665_ ;
wire _7245_ ;
wire _2380_ ;
wire _9410__bF$buf0 ;
wire _9410__bF$buf1 ;
wire _9410__bF$buf2 ;
wire _9410__bF$buf3 ;
wire _9410__bF$buf4 ;
wire _3585_ ;
wire _3165_ ;
wire _5731_ ;
wire _5311_ ;
wire [31:0] \datapath.registers.rega_data  ;
wire _809_ ;
wire _69_ ;
wire _6936_ ;
wire _6516_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _2856_ ;
wire _2436_ ;
wire _2016_ ;
wire _7894_ ;
wire _7474_ ;
wire _7054_ ;
wire _8679_ ;
wire _8259_ ;
wire _3394_ ;
wire _486__bF$buf0 ;
wire _486__bF$buf1 ;
wire _486__bF$buf2 ;
wire _486__bF$buf3 ;
wire _486__bF$buf4 ;
wire _9200_ ;
wire _1707_ ;
wire _4599_ ;
wire _4179_ ;
wire _5960_ ;
wire _5540_ ;
wire _5120_ ;
wire _618_ ;
wire _6745_ ;
wire _6325_ ;
wire _1880_ ;
wire _1460_ ;
wire _1040_ ;
wire _791_ ;
wire _371_ ;
wire _2665_ ;
wire _2245_ ;
wire _4811_ ;
wire _7283_ ;
wire _490__bF$buf0 ;
wire _490__bF$buf1 ;
wire _490__bF$buf2 ;
wire _490__bF$buf3 ;
wire _490__bF$buf4 ;
wire _8488_ ;
wire _8068_ ;
wire _1936_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire _6974_ ;
wire _6554_ ;
wire _6134_ ;
wire _180_ ;
wire _7759_ ;
wire _7339_ ;
wire _2894_ ;
wire _2474_ ;
wire _2054_ ;
wire _8700_ ;
wire _3679_ ;
wire _3259_ ;
wire _4620_ ;
wire _4200_ ;
wire _7092_ ;
wire _5825_ ;
wire _5405_ ;
wire _8297_ ;
wire _1745_ ;
wire _1325_ ;
wire _656_ ;
wire _236_ ;
wire _6783_ ;
wire _6363_ ;
wire _7988_ ;
wire _7568_ ;
wire _7148_ ;
wire _2283_ ;
wire _3488_ ;
wire _3068_ ;
wire _5634_ ;
wire _5214_ ;
wire _6839_ ;
wire _6419_ ;
wire _1974_ ;
wire _1554_ ;
wire _1134_ ;
wire _885_ ;
wire _465_ ;
wire _2759_ ;
wire _2339_ ;
wire _3700_ ;
wire _6592_ ;
wire _6172_ ;
wire _4905_ ;
wire _7797_ ;
wire _7377_ ;
wire _2092_ ;
wire _3297_ ;
wire _9103_ ;
wire _5863_ ;
wire _5443_ ;
wire _5023_ ;
wire _6648_ ;
wire _6228_ ;
wire _1783_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _2988_ ;
wire _2568_ ;
wire _2148_ ;
wire _4714_ ;
wire _7186_ ;
wire \datapath.idinstr_16_bF$buf0  ;
wire _5919_ ;
wire _9332_ ;
wire _1839_ ;
wire _1419_ ;
wire _5672_ ;
wire _5252_ ;
wire _6877_ ;
wire _6457_ ;
wire _6037_ ;
wire _1592_ ;
wire _1172_ ;
wire \datapath.idinstr_22_bF$buf39  ;
wire _2797_ ;
wire _2377_ ;
wire _8603_ ;
wire _4943_ ;
wire \datapath.idinstr_20_bF$buf0  ;
wire _4523_ ;
wire _4103_ ;
wire \bypassandflushunit.stall_bF$buf9  ;
wire _5728_ ;
wire _5308_ ;
wire _9141_ ;
wire _1648_ ;
wire _1228_ ;
wire _5481_ ;
wire _5061_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _6686_ ;
wire _6266_ ;
wire _2186_ ;
wire _8832_ ;
wire _8412_ ;
wire _5793__bF$buf0 ;
wire _5793__bF$buf1 ;
wire _5793__bF$buf2 ;
wire _5793__bF$buf3 ;
wire _5793__bF$buf4 ;
wire _4752_ ;
wire _4332_ ;
wire _5957_ ;
wire _5537_ ;
wire _5117_ ;
wire _31_ ;
wire _9370_ ;
wire _1877_ ;
wire _1457_ ;
wire _1037_ ;
wire _5290_ ;
wire _788_ ;
wire _368_ ;
wire \datapath.idinstr_17_hier0_bF$buf3  ;
wire _3603_ ;
wire _6495_ ;
wire _6075_ ;
wire _5478__bF$buf0 ;
wire _5478__bF$buf1 ;
wire _5478__bF$buf2 ;
wire _5478__bF$buf3 ;
wire _5478__bF$buf4 ;
wire _4808_ ;
wire _8641_ ;
wire _8221_ ;
wire _9426_ ;
wire _9006_ ;
wire _4981_ ;
wire _4561_ ;
wire _4141_ ;
wire \datapath.idinstr_19_bF$buf3  ;
wire _5766_ ;
wire _5346_ ;
wire _1686_ ;
wire _1266_ ;
wire _7912_ ;
wire _597_ ;
wire _177_ ;
wire _5482__bF$buf0 ;
wire _3832_ ;
wire _5482__bF$buf1 ;
wire _3412_ ;
wire _5482__bF$buf2 ;
wire _5482__bF$buf3 ;
wire _5482__bF$buf4 ;
wire _4617_ ;
wire _7089_ ;
wire _8870_ ;
wire _8450_ ;
wire _8030_ ;
wire _9235_ ;
wire _4790_ ;
wire _4370_ ;
wire \datapath.idinstr_23_bF$buf3  ;
wire _5995_ ;
wire _5575_ ;
wire _5155_ ;
wire _1495_ ;
wire _1075_ ;
wire _7721_ ;
wire _7301_ ;
wire _8926_ ;
wire _8506_ ;
wire _3641_ ;
wire _3221_ ;
wire _5580__bF$buf0 ;
wire _5580__bF$buf1 ;
wire _5580__bF$buf2 ;
wire _5580__bF$buf3 ;
wire _5580__bF$buf4 ;
wire _4846_ ;
wire _4426_ ;
wire _4006_ ;
wire _9044_ ;
wire _2912_ ;
wire _5384_ ;
wire _6589_ ;
wire _6169_ ;
wire _7950_ ;
wire _7530_ ;
wire _7110_ ;
wire _5505__bF$buf0 ;
wire _5505__bF$buf1 ;
wire _5505__bF$buf2 ;
wire _5505__bF$buf3 ;
wire _2089_ ;
wire _5505__bF$buf4 ;
wire _5505__bF$buf5 ;
wire _5505__bF$buf6 ;
wire _5505__bF$buf7 ;
wire _8735_ ;
wire _8315_ ;
wire _3870_ ;
wire _3450_ ;
wire _3030_ ;
wire _4655_ ;
wire _4235_ ;
wire _6801_ ;
wire _9273_ ;
wire _2721_ ;
wire _2301_ ;
wire _5193_ ;
wire _3926_ ;
wire _3506_ ;
wire _6398_ ;
wire _8964_ ;
wire _8544_ ;
wire _8124_ ;
wire _9329_ ;
wire _4884_ ;
wire _4464_ ;
wire _4044_ ;
wire _903_ ;
wire _5669_ ;
wire _5249_ ;
wire _6610_ ;
wire _9082_ ;
wire _1589_ ;
wire _1169_ ;
wire _7815_ ;
wire _2950_ ;
wire _2530_ ;
wire _2110_ ;
wire _3735_ ;
wire _3315_ ;
wire \datapath.alu.b_1_bF$buf4  ;
wire [31:0] \datapath.mempc  ;
wire _8773_ ;
wire _8353_ ;
wire _1801_ ;
wire _9138_ ;
wire _4693_ ;
wire _4273_ ;
wire _712_ ;
wire _5898_ ;
wire _5478_ ;
wire _5058_ ;
wire [31:0] \datapath.alu.a  ;
wire _1398_ ;
wire _7624_ ;
wire _7204_ ;
wire [31:0] \datapath.registers.1226[1]  ;
wire _8829_ ;
wire _8409_ ;
wire _3964_ ;
wire _3544_ ;
wire _3124_ ;
wire _4749_ ;
wire _4329_ ;
wire _8582_ ;
wire _8162_ ;
wire _28_ ;
wire _1610_ ;
wire _9367_ ;
wire _4082_ ;
wire \datapath.idinstr_20_bF$buf21  ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _2815_ ;
wire \controlunit.ebreak  ;
wire _5287_ ;
wire _7853_ ;
wire _7433_ ;
wire _7013_ ;
wire _8638_ ;
wire _8218_ ;
wire _3773_ ;
wire _3353_ ;
wire \datapath.idinstr_17_bF$buf15  ;
wire _4978_ ;
wire _4558_ ;
wire \datapath.idinstr_21_bF$buf30  ;
wire _4138_ ;
wire _8391_ ;
wire _6704_ ;
wire _9176_ ;
wire _750_ ;
wire _330_ ;
wire _7909_ ;
wire _2624_ ;
wire _2204_ ;
wire _5096_ ;
wire \datapath.idinstr_15_bF$buf35  ;
wire _3829_ ;
wire _3409_ ;
wire _7662_ ;
wire _7242_ ;
wire _8867_ ;
wire _8447_ ;
wire _8027_ ;
wire _3582_ ;
wire _3162_ ;
wire _4787_ ;
wire _4367_ ;
wire _806_ ;
wire \datapath.idinstr_16_bF$buf44  ;
wire _66_ ;
wire _6933_ ;
wire _6513_ ;
wire _7718_ ;
wire _2853_ ;
wire _2433_ ;
wire _2013_ ;
wire _3638_ ;
wire _3218_ ;
wire _7891_ ;
wire _7471_ ;
wire _7051_ ;
wire \bypassandflushunit.flushsystem  ;
wire _8676_ ;
wire _8256_ ;
wire _3391_ ;
wire _1704_ ;
wire _4596_ ;
wire _4176_ ;
wire _615_ ;
wire _2909_ ;
wire _6742_ ;
wire _6322_ ;
wire _7947_ ;
wire _7527_ ;
wire _7107_ ;
wire _2662_ ;
wire _2242_ ;
wire _3867_ ;
wire _3447_ ;
wire _3027_ ;
wire _7280_ ;
wire _8485_ ;
wire _8065_ ;
wire _1933_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire _2718_ ;
wire _6971_ ;
wire _6551_ ;
wire _6131_ ;
wire _7756_ ;
wire _7336_ ;
wire _2891_ ;
wire _2471_ ;
wire _2051_ ;
wire [31:0] \datapath.registers.1226[17]  ;
wire _3676_ ;
wire _3256_ ;
wire _5822_ ;
wire _5402_ ;
wire _8294_ ;
wire [31:0] \datapath.idinstr  ;
wire _6607_ ;
wire _1742_ ;
wire _1322_ ;
wire _9079_ ;
wire _653_ ;
wire _233_ ;
wire _2947_ ;
wire _2527_ ;
wire _2107_ ;
wire _6780_ ;
wire _6360_ ;
wire _7985_ ;
wire _7565_ ;
wire _7145_ ;
wire _2280_ ;
wire _3485_ ;
wire _3065_ ;
wire _5631_ ;
wire _5211_ ;
wire _709_ ;
wire _6836_ ;
wire _6416_ ;
wire _1971_ ;
wire _1551_ ;
wire _1131_ ;
wire _882_ ;
wire _462_ ;
wire _2756_ ;
wire _2336_ ;
wire _4902_ ;
wire _7794_ ;
wire _7374_ ;
wire _8999_ ;
wire _8579_ ;
wire _8159_ ;
wire _3294_ ;
wire _9100_ ;
wire _1607_ ;
wire _4499_ ;
wire _4079_ ;
wire _5860_ ;
wire _5440_ ;
wire _5020_ ;
wire \datapath.idinstr_20_bF$buf18  ;
wire _938_ ;
wire _518_ ;
wire _6645_ ;
wire _6225_ ;
wire _1780_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _2985_ ;
wire _2565_ ;
wire _2145_ ;
wire _4711_ ;
wire _7183_ ;
wire \datapath.idinstr_21_bF$buf27  ;
wire _5916_ ;
wire _8388_ ;
wire _1836_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _6874_ ;
wire _6454_ ;
wire _6034_ ;
wire \datapath.idinstr_22_bF$buf36  ;
wire _7659_ ;
wire _7239_ ;
wire _2794_ ;
wire _2374_ ;
wire _8600_ ;
wire _3999_ ;
wire _3579_ ;
wire _3159_ ;
wire _4940_ ;
wire _4520_ ;
wire _4100_ ;
wire \bypassandflushunit.stall_bF$buf6  ;
wire _5725_ ;
wire _5305_ ;
wire _8197_ ;
wire _1645_ ;
wire _1225_ ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire _6683_ ;
wire _6263_ ;
wire _7888_ ;
wire _7468_ ;
wire _7048_ ;
wire _2183_ ;
wire _3388_ ;
wire _5954_ ;
wire _5534_ ;
wire _5114_ ;
wire _6739_ ;
wire _6319_ ;
wire _1874_ ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _2659_ ;
wire _2239_ ;
wire \datapath.idinstr_17_hier0_bF$buf0  ;
wire _3600_ ;
wire _6492_ ;
wire _6072_ ;
wire _4805_ ;
wire _7697_ ;
wire _7277_ ;
wire [31:0] \datapath.regloadwb  ;
wire _3197_ ;
wire _9423_ ;
wire _9003_ ;
wire \datapath.idinstr_19_bF$buf0  ;
wire _5763_ ;
wire _5343_ ;
wire _6968_ ;
wire _6548_ ;
wire _6128_ ;
wire _1683_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _2888_ ;
wire _2468_ ;
wire _2048_ ;
wire _4614_ ;
wire _7086_ ;
wire _5819_ ;
wire _9232_ ;
wire _1739_ ;
wire _1319_ ;
wire \datapath.idinstr_23_bF$buf0  ;
wire _5992_ ;
wire _5572_ ;
wire _5152_ ;
wire _6777_ ;
wire _6357_ ;
wire _1492_ ;
wire _1072_ ;
wire _2697_ ;
wire _2277_ ;
wire _8923_ ;
wire _8503_ ;
wire _4843_ ;
wire _4423_ ;
wire _4003_ ;
wire _5628_ ;
wire _5208_ ;
wire _9041_ ;
wire _1968_ ;
wire _1548_ ;
wire _1128_ ;
wire _5381_ ;
wire _879_ ;
wire _459_ ;
wire _6586_ ;
wire _6166_ ;
wire _2086_ ;
wire _8732_ ;
wire _8312_ ;
wire _4652_ ;
wire _4232_ ;
wire _5857_ ;
wire _5437_ ;
wire _5017_ ;
wire _9270_ ;
wire _1777_ ;
wire _1357_ ;
wire _5190_ ;
wire _688_ ;
wire _268_ ;
wire _3923_ ;
wire _3503_ ;
wire _6395_ ;
wire _4708_ ;
wire _8961_ ;
wire _8541_ ;
wire _8121_ ;
wire _9326_ ;
wire _4881_ ;
wire _4461_ ;
wire _4041_ ;
wire [3:0] \datapath.alu.funsel  ;
wire _5579__bF$buf0 ;
wire _5579__bF$buf1 ;
wire _900_ ;
wire _5579__bF$buf2 ;
wire _5579__bF$buf3 ;
wire _5579__bF$buf4 ;
wire _5579__bF$buf5 ;
wire _5666_ ;
wire _5246_ ;
wire \datapath.idinstr_17_bF$buf9  ;
wire _1586_ ;
wire _1166_ ;
wire _7812_ ;
wire _497_ ;
wire _3732_ ;
wire _3312_ ;
wire \datapath.alu.b_1_bF$buf1  ;
wire _4937_ ;
wire _4517_ ;
wire _8770_ ;
wire _8350_ ;
wire _9135_ ;
wire _4690_ ;
wire _4270_ ;
wire \datapath.idinstr_21_bF$buf9  ;
wire _5895_ ;
wire _5475_ ;
wire _5055_ ;
wire _1395_ ;
wire _7621_ ;
wire _7201_ ;
wire _8826_ ;
wire _8406_ ;
wire _3961_ ;
wire _3541_ ;
wire _3121_ ;
wire _4746_ ;
wire _4326_ ;
wire [2:0] \datapath.aluexecptions  ;
wire _25_ ;
wire _9364_ ;
wire _2812_ ;
wire _5284_ ;
wire _6489_ ;
wire _6069_ ;
wire _7850_ ;
wire _7430_ ;
wire _7010_ ;
wire _8635_ ;
wire _8215_ ;
wire _3770_ ;
wire _3350_ ;
wire \datapath.idinstr_17_bF$buf12  ;
wire _4975_ ;
wire _4555_ ;
wire _4135_ ;
wire _6701_ ;
wire _9173_ ;
wire _7906_ ;
wire _2621_ ;
wire _2201_ ;
wire _5093_ ;
wire \datapath.idinstr_15_bF$buf32  ;
wire _3826_ ;
wire _3406_ ;
wire _6298_ ;
wire _8864_ ;
wire _8444_ ;
wire _8024_ ;
wire _5859__bF$buf0 ;
wire _5859__bF$buf1 ;
wire _5859__bF$buf2 ;
wire _5859__bF$buf3 ;
wire _5859__bF$buf4 ;
wire _5859__bF$buf5 ;
wire _5859__bF$buf6 ;
wire _5859__bF$buf7 ;
wire \datapath.alu.b_4_bF$buf4  ;
wire _9229_ ;
wire _4784_ ;
wire _4364_ ;
wire _803_ ;
wire _5989_ ;
wire _5569_ ;
wire _5149_ ;
wire \datapath.idinstr_16_bF$buf41  ;
wire _63_ ;
wire _6930_ ;
wire _6510_ ;
wire _1489_ ;
wire _1069_ ;
wire _7715_ ;
wire _2850_ ;
wire _2430_ ;
wire _2010_ ;
wire _3635_ ;
wire _3215_ ;
wire _8673_ ;
wire _8253_ ;
wire _1701_ ;
wire _9038_ ;
wire _4593_ ;
wire _4173_ ;
wire _612_ ;
wire _2906_ ;
wire _5798_ ;
wire _5378_ ;
wire [1:0] bsel ;
wire _1298_ ;
wire _7944_ ;
wire _7524_ ;
wire _7104_ ;
wire _8729_ ;
wire _8309_ ;
wire _3864_ ;
wire _3444_ ;
wire _3024_ ;
wire _4649_ ;
wire _4229_ ;
wire _8482_ ;
wire CLK_bF$buf80 ;
wire _8062_ ;
wire CLK_bF$buf81 ;
wire CLK_bF$buf82 ;
wire CLK_bF$buf83 ;
wire CLK_bF$buf84 ;
wire CLK_bF$buf85 ;
wire CLK_bF$buf86 ;
wire CLK_bF$buf87 ;
wire CLK_bF$buf88 ;
wire CLK_bF$buf89 ;
wire _1930_ ;
wire _1510_ ;
wire _9267_ ;
wire _841_ ;
wire _421_ ;
wire _2715_ ;
wire _5187_ ;
wire _7753_ ;
wire _7333_ ;
wire _8958_ ;
wire _8538_ ;
wire _8118_ ;
wire _3673_ ;
wire _3253_ ;
wire _4878_ ;
wire _4458_ ;
wire _4038_ ;
wire _8291_ ;
wire _6604_ ;
wire _9076_ ;
wire _650_ ;
wire _230_ ;
wire _7809_ ;
wire _2944_ ;
wire _2524_ ;
wire _2104_ ;
wire _3729_ ;
wire _3309_ ;
wire _7982_ ;
wire _7562_ ;
wire _7142_ ;
wire _8767_ ;
wire _8347_ ;
wire _3482_ ;
wire _3062_ ;
wire _4687_ ;
wire _4267_ ;
wire _706_ ;
wire _6833_ ;
wire _6413_ ;
wire _7618_ ;
wire _2753_ ;
wire _2333_ ;
wire _3958_ ;
wire _3538_ ;
wire _3118_ ;
wire _5429__bF$buf0 ;
wire _5429__bF$buf1 ;
wire _7791_ ;
wire _5429__bF$buf2 ;
wire _7371_ ;
wire _5429__bF$buf3 ;
wire _5429__bF$buf4 ;
wire _8996_ ;
wire _8576_ ;
wire _8156_ ;
wire \datapath.csr._20_  ;
wire _3291_ ;
wire _1604_ ;
wire _4496_ ;
wire _4076_ ;
wire \datapath.idinstr_20_bF$buf15  ;
wire _935_ ;
wire _515_ ;
wire _2809_ ;
wire _6642_ ;
wire _6222_ ;
wire _7847_ ;
wire _7427_ ;
wire _7007_ ;
wire _2982_ ;
wire _2562_ ;
wire _2142_ ;
wire _3767_ ;
wire _3347_ ;
wire _7180_ ;
wire \datapath.idinstr_21_bF$buf24  ;
wire _5913_ ;
wire _8385_ ;
wire [2:0] \controlunit.imm_sel  ;
wire _1833_ ;
wire _1413_ ;
wire _744_ ;
wire _324_ ;
wire _2618_ ;
wire _6871_ ;
wire _6451_ ;
wire _6031_ ;
wire \datapath.idinstr_15_bF$buf29  ;
wire \datapath.idinstr_22_bF$buf33  ;
wire _7656_ ;
wire _7236_ ;
wire _2791_ ;
wire _2371_ ;
wire _3996_ ;
wire _3576_ ;
wire _3156_ ;
wire \bypassandflushunit.stall_bF$buf3  ;
wire _5722_ ;
wire _5302_ ;
wire _8194_ ;
wire \datapath.idinstr_16_bF$buf38  ;
wire _6927_ ;
wire _6507_ ;
wire _1642_ ;
wire _1222_ ;
wire _9399_ ;
wire \datapath.idinstr_20_bF$buf53  ;
wire _973_ ;
wire _553_ ;
wire _133_ ;
wire _2847_ ;
wire _2427_ ;
wire _2007_ ;
wire _6680_ ;
wire _6260_ ;
wire _7885_ ;
wire _7465_ ;
wire _7045_ ;
wire _2180_ ;
wire _3385_ ;
wire _5951_ ;
wire _5531_ ;
wire _5111_ ;
wire _609_ ;
wire _6736_ ;
wire _6316_ ;
wire _1871_ ;
wire _1451_ ;
wire _1031_ ;
wire _782_ ;
wire _362_ ;
wire _2656_ ;
wire _2236_ ;
wire _4802_ ;
wire _7694_ ;
wire _7274_ ;
wire [31:0] \datapath.registers.1226[8]  ;
wire _8899_ ;
wire _8479_ ;
wire _8059_ ;
wire _3194_ ;
wire _9420_ ;
wire _9000_ ;
wire _1927_ ;
wire _1507_ ;
wire _4399_ ;
wire _5760_ ;
wire _5340_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _6965_ ;
wire _6545_ ;
wire _6125_ ;
wire _1680_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _2885_ ;
wire _2465_ ;
wire _2045_ ;
wire _4611_ ;
wire _7083_ ;
wire _5816_ ;
wire _8288_ ;
wire _1736_ ;
wire _1316_ ;
wire _3798__bF$buf0 ;
wire _3798__bF$buf1 ;
wire _3798__bF$buf2 ;
wire _3798__bF$buf3 ;
wire _3798__bF$buf4 ;
wire _647_ ;
wire _227_ ;
wire _6774_ ;
wire _6354_ ;
wire \datapath._51_  ;
wire _7979_ ;
wire _7559_ ;
wire _7139_ ;
wire _2694_ ;
wire _2274_ ;
wire _8920_ ;
wire _8500_ ;
wire _3899_ ;
wire _3479_ ;
wire _3059_ ;
wire _4840_ ;
wire _4420_ ;
wire _4000_ ;
wire _5625_ ;
wire _5205_ ;
wire _8097_ ;
wire _1965_ ;
wire _1545_ ;
wire _1125_ ;
wire [31:0] \datapath.wbinstr  ;
wire _876_ ;
wire _456_ ;
wire _6583_ ;
wire _6163_ ;
wire _7788_ ;
wire _7368_ ;
wire _2083_ ;
wire _3288_ ;
wire _5854_ ;
wire _5434_ ;
wire _5014_ ;
wire [1:0] \datapath.csr._37_  ;
wire _6639_ ;
wire _6219_ ;
wire _1774_ ;
wire _1354_ ;
wire _685_ ;
wire _265_ ;
wire _2979_ ;
wire _2559_ ;
wire _2139_ ;
wire _3920_ ;
wire _3500_ ;
wire _6392_ ;
wire _4705_ ;
wire _7597_ ;
wire _7177_ ;
wire _3097_ ;
wire _9323_ ;
wire _5663_ ;
wire _5243_ ;
wire \datapath.idinstr_17_bF$buf6  ;
wire _6868_ ;
wire _6448_ ;
wire _6028_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _2788_ ;
wire _2368_ ;
wire [31:0] \datapath.nextpc  ;
wire _4934_ ;
wire _4514_ ;
wire _5719_ ;
wire _9132_ ;
wire _1639_ ;
wire _1219_ ;
wire \datapath.idinstr_21_bF$buf6  ;
wire _5892_ ;
wire _5472_ ;
wire _5052_ ;
wire _6677_ ;
wire _6257_ ;
wire _1392_ ;
wire _2597_ ;
wire _2177_ ;
wire _8823_ ;
wire _8403_ ;
wire _4743_ ;
wire _4323_ ;
wire _5948_ ;
wire _5528_ ;
wire _5108_ ;
wire _22_ ;
wire _9361_ ;
wire _1868_ ;
wire _1448_ ;
wire _1028_ ;
wire _5281_ ;
wire _779_ ;
wire _359_ ;
wire _6486_ ;
wire _6066_ ;
wire _8632_ ;
wire _8212_ ;

BUFX2 BUFX2_insert1463 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [16]),
    .Y(\datapath.idinstr_16_hier0_bF$buf0 )
);

BUFX2 BUFX2_insert1462 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [16]),
    .Y(\datapath.idinstr_16_hier0_bF$buf1 )
);

BUFX2 BUFX2_insert1461 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [16]),
    .Y(\datapath.idinstr_16_hier0_bF$buf2 )
);

BUFX2 BUFX2_insert1460 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [16]),
    .Y(\datapath.idinstr_16_hier0_bF$buf3 )
);

BUFX2 BUFX2_insert1459 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [16]),
    .Y(\datapath.idinstr_16_hier0_bF$buf4 )
);

BUFX2 BUFX2_insert1458 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [16]),
    .Y(\datapath.idinstr_16_hier0_bF$buf5 )
);

BUFX2 BUFX2_insert1457 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [22]),
    .Y(\datapath.idinstr_22_hier0_bF$buf0 )
);

BUFX2 BUFX2_insert1456 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [22]),
    .Y(\datapath.idinstr_22_hier0_bF$buf1 )
);

BUFX2 BUFX2_insert1455 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [22]),
    .Y(\datapath.idinstr_22_hier0_bF$buf2 )
);

BUFX2 BUFX2_insert1454 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [22]),
    .Y(\datapath.idinstr_22_hier0_bF$buf3 )
);

BUFX2 BUFX2_insert1453 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [22]),
    .Y(\datapath.idinstr_22_hier0_bF$buf4 )
);

BUFX2 BUFX2_insert1452 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [22]),
    .Y(\datapath.idinstr_22_hier0_bF$buf5 )
);

CLKBUF1 CLKBUF1_insert1451 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK),
    .Y(CLK_hier0_bF$buf0)
);

CLKBUF1 CLKBUF1_insert1450 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK),
    .Y(CLK_hier0_bF$buf1)
);

CLKBUF1 CLKBUF1_insert1449 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK),
    .Y(CLK_hier0_bF$buf2)
);

CLKBUF1 CLKBUF1_insert1448 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK),
    .Y(CLK_hier0_bF$buf3)
);

CLKBUF1 CLKBUF1_insert1447 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK),
    .Y(CLK_hier0_bF$buf4)
);

CLKBUF1 CLKBUF1_insert1446 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK),
    .Y(CLK_hier0_bF$buf5)
);

CLKBUF1 CLKBUF1_insert1445 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK),
    .Y(CLK_hier0_bF$buf6)
);

CLKBUF1 CLKBUF1_insert1444 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK),
    .Y(CLK_hier0_bF$buf7)
);

CLKBUF1 CLKBUF1_insert1443 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK),
    .Y(CLK_hier0_bF$buf8)
);

CLKBUF1 CLKBUF1_insert1442 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK),
    .Y(CLK_hier0_bF$buf9)
);

CLKBUF1 CLKBUF1_insert1441 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK),
    .Y(CLK_hier0_bF$buf10)
);

CLKBUF1 CLKBUF1_insert1440 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK),
    .Y(CLK_hier0_bF$buf11)
);

BUFX2 BUFX2_insert1439 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_hier0_bF$buf0 )
);

BUFX2 BUFX2_insert1438 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_hier0_bF$buf1 )
);

BUFX2 BUFX2_insert1437 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_hier0_bF$buf2 )
);

BUFX2 BUFX2_insert1436 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_hier0_bF$buf3 )
);

BUFX2 BUFX2_insert1435 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_hier0_bF$buf4 )
);

BUFX2 BUFX2_insert1434 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [17]),
    .Y(\datapath.idinstr_17_hier0_bF$buf5 )
);

BUFX2 BUFX2_insert1433 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [20]),
    .Y(\datapath.idinstr_20_hier0_bF$buf0 )
);

BUFX2 BUFX2_insert1432 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [20]),
    .Y(\datapath.idinstr_20_hier0_bF$buf1 )
);

BUFX2 BUFX2_insert1431 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [20]),
    .Y(\datapath.idinstr_20_hier0_bF$buf2 )
);

BUFX2 BUFX2_insert1430 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [20]),
    .Y(\datapath.idinstr_20_hier0_bF$buf3 )
);

BUFX2 BUFX2_insert1429 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [20]),
    .Y(\datapath.idinstr_20_hier0_bF$buf4 )
);

BUFX2 BUFX2_insert1428 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [20]),
    .Y(\datapath.idinstr_20_hier0_bF$buf5 )
);

BUFX2 BUFX2_insert1427 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [20]),
    .Y(\datapath.idinstr_20_hier0_bF$buf6 )
);

BUFX2 BUFX2_insert1426 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [15]),
    .Y(\datapath.idinstr_15_hier0_bF$buf0 )
);

BUFX2 BUFX2_insert1425 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [15]),
    .Y(\datapath.idinstr_15_hier0_bF$buf1 )
);

BUFX2 BUFX2_insert1424 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [15]),
    .Y(\datapath.idinstr_15_hier0_bF$buf2 )
);

BUFX2 BUFX2_insert1423 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [15]),
    .Y(\datapath.idinstr_15_hier0_bF$buf3 )
);

BUFX2 BUFX2_insert1422 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [15]),
    .Y(\datapath.idinstr_15_hier0_bF$buf4 )
);

BUFX2 BUFX2_insert1421 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [15]),
    .Y(\datapath.idinstr_15_hier0_bF$buf5 )
);

BUFX2 BUFX2_insert1420 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [15]),
    .Y(\datapath.idinstr_15_hier0_bF$buf6 )
);

BUFX2 BUFX2_insert1419 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [21]),
    .Y(\datapath.idinstr_21_hier0_bF$buf0 )
);

BUFX2 BUFX2_insert1418 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [21]),
    .Y(\datapath.idinstr_21_hier0_bF$buf1 )
);

BUFX2 BUFX2_insert1417 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [21]),
    .Y(\datapath.idinstr_21_hier0_bF$buf2 )
);

BUFX2 BUFX2_insert1416 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [21]),
    .Y(\datapath.idinstr_21_hier0_bF$buf3 )
);

BUFX2 BUFX2_insert1415 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [21]),
    .Y(\datapath.idinstr_21_hier0_bF$buf4 )
);

BUFX2 BUFX2_insert1414 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [21]),
    .Y(\datapath.idinstr_21_hier0_bF$buf5 )
);

BUFX2 BUFX2_insert1413 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472_),
    .Y(_5472__bF$buf0)
);

BUFX2 BUFX2_insert1412 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472_),
    .Y(_5472__bF$buf1)
);

BUFX2 BUFX2_insert1411 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472_),
    .Y(_5472__bF$buf2)
);

BUFX2 BUFX2_insert1410 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472_),
    .Y(_5472__bF$buf3)
);

BUFX2 BUFX2_insert1409 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472_),
    .Y(_5472__bF$buf4)
);

BUFX2 BUFX2_insert1408 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_494_),
    .Y(_494__bF$buf0)
);

BUFX2 BUFX2_insert1407 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_494_),
    .Y(_494__bF$buf1)
);

BUFX2 BUFX2_insert1406 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_494_),
    .Y(_494__bF$buf2)
);

BUFX2 BUFX2_insert1405 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_494_),
    .Y(_494__bF$buf3)
);

BUFX2 BUFX2_insert1404 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_494_),
    .Y(_494__bF$buf4)
);

BUFX2 BUFX2_insert1403 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5434_),
    .Y(_5434__bF$buf0)
);

BUFX2 BUFX2_insert1402 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5434_),
    .Y(_5434__bF$buf1)
);

BUFX2 BUFX2_insert1401 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5434_),
    .Y(_5434__bF$buf2)
);

BUFX2 BUFX2_insert1400 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5434_),
    .Y(_5434__bF$buf3)
);

BUFX2 BUFX2_insert1399 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5434_),
    .Y(_5434__bF$buf4)
);

BUFX2 BUFX2_insert1398 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5434_),
    .Y(_5434__bF$buf5)
);

BUFX2 BUFX2_insert1397 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5434_),
    .Y(_5434__bF$buf6)
);

BUFX2 BUFX2_insert1396 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5434_),
    .Y(_5434__bF$buf7)
);

BUFX2 BUFX2_insert1395 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5434_),
    .Y(_5434__bF$buf8)
);

BUFX2 BUFX2_insert1394 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5434_),
    .Y(_5434__bF$buf9)
);

BUFX2 BUFX2_insert1393 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5434_),
    .Y(_5434__bF$buf10)
);

BUFX2 BUFX2_insert1392 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5434_),
    .Y(_5434__bF$buf11)
);

BUFX2 BUFX2_insert1391 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5434_),
    .Y(_5434__bF$buf12)
);

BUFX2 BUFX2_insert1390 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5434_),
    .Y(_5434__bF$buf13)
);

BUFX2 BUFX2_insert1389 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5434_),
    .Y(_5434__bF$buf14)
);

BUFX2 BUFX2_insert1388 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760_),
    .Y(_5760__bF$buf0)
);

BUFX2 BUFX2_insert1387 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760_),
    .Y(_5760__bF$buf1)
);

BUFX2 BUFX2_insert1386 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760_),
    .Y(_5760__bF$buf2)
);

BUFX2 BUFX2_insert1385 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760_),
    .Y(_5760__bF$buf3)
);

BUFX2 BUFX2_insert1384 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760_),
    .Y(_5760__bF$buf4)
);

BUFX2 BUFX2_insert1383 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760_),
    .Y(_5760__bF$buf5)
);

BUFX2 BUFX2_insert1382 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760_),
    .Y(_5760__bF$buf6)
);

BUFX2 BUFX2_insert1381 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760_),
    .Y(_5760__bF$buf7)
);

BUFX2 BUFX2_insert1380 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760_),
    .Y(_5760__bF$buf8)
);

BUFX2 BUFX2_insert1379 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_609_),
    .Y(_609__bF$buf0)
);

BUFX2 BUFX2_insert1378 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_609_),
    .Y(_609__bF$buf1)
);

BUFX2 BUFX2_insert1377 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_609_),
    .Y(_609__bF$buf2)
);

BUFX2 BUFX2_insert1376 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_609_),
    .Y(_609__bF$buf3)
);

BUFX2 BUFX2_insert1375 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_609_),
    .Y(_609__bF$buf4)
);

BUFX2 BUFX2_insert1374 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076_),
    .Y(_9076__bF$buf0)
);

BUFX2 BUFX2_insert1373 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076_),
    .Y(_9076__bF$buf1)
);

BUFX2 BUFX2_insert1372 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076_),
    .Y(_9076__bF$buf2)
);

BUFX2 BUFX2_insert1371 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076_),
    .Y(_9076__bF$buf3)
);

BUFX2 BUFX2_insert1370 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076_),
    .Y(_9076__bF$buf4)
);

BUFX2 BUFX2_insert1369 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076_),
    .Y(_9076__bF$buf5)
);

BUFX2 BUFX2_insert1368 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076_),
    .Y(_9076__bF$buf6)
);

BUFX2 BUFX2_insert1367 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076_),
    .Y(_9076__bF$buf7)
);

BUFX2 BUFX2_insert1366 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076_),
    .Y(_9076__bF$buf8)
);

BUFX2 BUFX2_insert1365 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_497_),
    .Y(_497__bF$buf0)
);

BUFX2 BUFX2_insert1364 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_497_),
    .Y(_497__bF$buf1)
);

BUFX2 BUFX2_insert1363 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_497_),
    .Y(_497__bF$buf2)
);

BUFX2 BUFX2_insert1362 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_497_),
    .Y(_497__bF$buf3)
);

BUFX2 BUFX2_insert1361 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_497_),
    .Y(_497__bF$buf4)
);

BUFX2 BUFX2_insert1360 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9041_),
    .Y(_9041__bF$buf0)
);

BUFX2 BUFX2_insert1359 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9041_),
    .Y(_9041__bF$buf1)
);

BUFX2 BUFX2_insert1358 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9041_),
    .Y(_9041__bF$buf2)
);

BUFX2 BUFX2_insert1357 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9041_),
    .Y(_9041__bF$buf3)
);

BUFX2 BUFX2_insert1356 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9041_),
    .Y(_9041__bF$buf4)
);

BUFX2 BUFX2_insert1355 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9041_),
    .Y(_9041__bF$buf5)
);

BUFX2 BUFX2_insert1354 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9041_),
    .Y(_9041__bF$buf6)
);

BUFX2 BUFX2_insert1353 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9041_),
    .Y(_9041__bF$buf7)
);

BUFX2 BUFX2_insert1352 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440_),
    .Y(_5440__bF$buf0)
);

BUFX2 BUFX2_insert1351 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440_),
    .Y(_5440__bF$buf1)
);

BUFX2 BUFX2_insert1350 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440_),
    .Y(_5440__bF$buf2)
);

BUFX2 BUFX2_insert1349 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440_),
    .Y(_5440__bF$buf3)
);

BUFX2 BUFX2_insert1348 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440_),
    .Y(_5440__bF$buf4)
);

BUFX2 BUFX2_insert1347 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478_),
    .Y(_5478__bF$buf0)
);

BUFX2 BUFX2_insert1346 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478_),
    .Y(_5478__bF$buf1)
);

BUFX2 BUFX2_insert1345 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478_),
    .Y(_5478__bF$buf2)
);

BUFX2 BUFX2_insert1344 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478_),
    .Y(_5478__bF$buf3)
);

BUFX2 BUFX2_insert1343 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478_),
    .Y(_5478__bF$buf4)
);

BUFX2 BUFX2_insert1342 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_597_),
    .Y(_597__bF$buf0)
);

BUFX2 BUFX2_insert1341 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_597_),
    .Y(_597__bF$buf1)
);

BUFX2 BUFX2_insert1340 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_597_),
    .Y(_597__bF$buf2)
);

BUFX2 BUFX2_insert1339 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_597_),
    .Y(_597__bF$buf3)
);

BUFX2 BUFX2_insert1338 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_597_),
    .Y(_597__bF$buf4)
);

BUFX2 BUFX2_insert1337 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_979_),
    .Y(_979__bF$buf0)
);

BUFX2 BUFX2_insert1336 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_979_),
    .Y(_979__bF$buf1)
);

BUFX2 BUFX2_insert1335 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_979_),
    .Y(_979__bF$buf2)
);

BUFX2 BUFX2_insert1334 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_979_),
    .Y(_979__bF$buf3)
);

BUFX2 BUFX2_insert1333 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_979_),
    .Y(_979__bF$buf4)
);

BUFX2 BUFX2_insert1332 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5960_),
    .Y(_5960__bF$buf0)
);

BUFX2 BUFX2_insert1331 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5960_),
    .Y(_5960__bF$buf1)
);

BUFX2 BUFX2_insert1330 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5960_),
    .Y(_5960__bF$buf2)
);

BUFX2 BUFX2_insert1329 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5960_),
    .Y(_5960__bF$buf3)
);

BUFX2 BUFX2_insert1328 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5960_),
    .Y(_5960__bF$buf4)
);

BUFX2 BUFX2_insert1327 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_982_),
    .Y(_982__bF$buf0)
);

BUFX2 BUFX2_insert1326 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_982_),
    .Y(_982__bF$buf1)
);

BUFX2 BUFX2_insert1325 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_982_),
    .Y(_982__bF$buf2)
);

BUFX2 BUFX2_insert1324 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_982_),
    .Y(_982__bF$buf3)
);

BUFX2 BUFX2_insert1323 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_982_),
    .Y(_982__bF$buf4)
);

BUFX2 BUFX2_insert1322 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040_),
    .Y(_6040__bF$buf0)
);

BUFX2 BUFX2_insert1321 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040_),
    .Y(_6040__bF$buf1)
);

BUFX2 BUFX2_insert1320 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040_),
    .Y(_6040__bF$buf2)
);

BUFX2 BUFX2_insert1319 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040_),
    .Y(_6040__bF$buf3)
);

BUFX2 BUFX2_insert1318 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040_),
    .Y(_6040__bF$buf4)
);

BUFX2 BUFX2_insert1317 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484_),
    .Y(_5484__bF$buf0)
);

BUFX2 BUFX2_insert1316 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484_),
    .Y(_5484__bF$buf1)
);

BUFX2 BUFX2_insert1315 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484_),
    .Y(_5484__bF$buf2)
);

BUFX2 BUFX2_insert1314 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484_),
    .Y(_5484__bF$buf3)
);

BUFX2 BUFX2_insert1313 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484_),
    .Y(_5484__bF$buf4)
);

BUFX2 BUFX2_insert1312 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446_),
    .Y(_5446__bF$buf0)
);

BUFX2 BUFX2_insert1311 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446_),
    .Y(_5446__bF$buf1)
);

BUFX2 BUFX2_insert1310 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446_),
    .Y(_5446__bF$buf2)
);

BUFX2 BUFX2_insert1309 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446_),
    .Y(_5446__bF$buf3)
);

BUFX2 BUFX2_insert1308 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446_),
    .Y(_5446__bF$buf4)
);

BUFX2 BUFX2_insert1307 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap ),
    .Y(\datapath.regcsrtrap_bF$buf0 )
);

BUFX2 BUFX2_insert1306 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap ),
    .Y(\datapath.regcsrtrap_bF$buf1 )
);

BUFX2 BUFX2_insert1305 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap ),
    .Y(\datapath.regcsrtrap_bF$buf2 )
);

BUFX2 BUFX2_insert1304 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap ),
    .Y(\datapath.regcsrtrap_bF$buf3 )
);

BUFX2 BUFX2_insert1303 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap ),
    .Y(\datapath.regcsrtrap_bF$buf4 )
);

BUFX2 BUFX2_insert1302 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap ),
    .Y(\datapath.regcsrtrap_bF$buf5 )
);

BUFX2 BUFX2_insert1301 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap ),
    .Y(\datapath.regcsrtrap_bF$buf6 )
);

BUFX2 BUFX2_insert1300 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap ),
    .Y(\datapath.regcsrtrap_bF$buf7 )
);

BUFX2 BUFX2_insert1299 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3800_),
    .Y(_3800__bF$buf0)
);

BUFX2 BUFX2_insert1298 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3800_),
    .Y(_3800__bF$buf1)
);

BUFX2 BUFX2_insert1297 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3800_),
    .Y(_3800__bF$buf2)
);

BUFX2 BUFX2_insert1296 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3800_),
    .Y(_3800__bF$buf3)
);

BUFX2 BUFX2_insert1295 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3800_),
    .Y(_3800__bF$buf4)
);

BUFX2 BUFX2_insert1294 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3800_),
    .Y(_3800__bF$buf5)
);

BUFX2 BUFX2_insert1293 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3800_),
    .Y(_3800__bF$buf6)
);

BUFX2 BUFX2_insert1292 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3800_),
    .Y(_3800__bF$buf7)
);

BUFX2 BUFX2_insert1291 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5505_),
    .Y(_5505__bF$buf0)
);

BUFX2 BUFX2_insert1290 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5505_),
    .Y(_5505__bF$buf1)
);

BUFX2 BUFX2_insert1289 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5505_),
    .Y(_5505__bF$buf2)
);

BUFX2 BUFX2_insert1288 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5505_),
    .Y(_5505__bF$buf3)
);

BUFX2 BUFX2_insert1287 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5505_),
    .Y(_5505__bF$buf4)
);

BUFX2 BUFX2_insert1286 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5505_),
    .Y(_5505__bF$buf5)
);

BUFX2 BUFX2_insert1285 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5505_),
    .Y(_5505__bF$buf6)
);

BUFX2 BUFX2_insert1284 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5505_),
    .Y(_5505__bF$buf7)
);

BUFX2 BUFX2_insert1283 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685_),
    .Y(_3685__bF$buf0)
);

BUFX2 BUFX2_insert1282 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685_),
    .Y(_3685__bF$buf1)
);

BUFX2 BUFX2_insert1281 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685_),
    .Y(_3685__bF$buf2)
);

BUFX2 BUFX2_insert1280 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685_),
    .Y(_3685__bF$buf3)
);

BUFX2 BUFX2_insert1279 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685_),
    .Y(_3685__bF$buf4)
);

BUFX2 BUFX2_insert1278 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480_),
    .Y(_2480__bF$buf0)
);

BUFX2 BUFX2_insert1277 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480_),
    .Y(_2480__bF$buf1)
);

BUFX2 BUFX2_insert1276 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480_),
    .Y(_2480__bF$buf2)
);

BUFX2 BUFX2_insert1275 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480_),
    .Y(_2480__bF$buf3)
);

BUFX2 BUFX2_insert1274 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480_),
    .Y(_2480__bF$buf4)
);

BUFX2 BUFX2_insert1273 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480_),
    .Y(_2480__bF$buf5)
);

BUFX2 BUFX2_insert1272 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6140_),
    .Y(_6140__bF$buf0)
);

BUFX2 BUFX2_insert1271 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6140_),
    .Y(_6140__bF$buf1)
);

BUFX2 BUFX2_insert1270 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6140_),
    .Y(_6140__bF$buf2)
);

BUFX2 BUFX2_insert1269 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6140_),
    .Y(_6140__bF$buf3)
);

BUFX2 BUFX2_insert1268 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6140_),
    .Y(_6140__bF$buf4)
);

BUFX2 BUFX2_insert1267 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_16_bF$buf0 )
);

BUFX2 BUFX2_insert1266 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_16_bF$buf1 )
);

BUFX2 BUFX2_insert1265 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_16_bF$buf2 )
);

BUFX2 BUFX2_insert1264 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_16_bF$buf3 )
);

BUFX2 BUFX2_insert1263 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_16_bF$buf4 )
);

BUFX2 BUFX2_insert1262 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_16_bF$buf5 )
);

BUFX2 BUFX2_insert1261 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_16_bF$buf6 )
);

BUFX2 BUFX2_insert1260 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_16_bF$buf7 )
);

BUFX2 BUFX2_insert1259 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_16_bF$buf8 )
);

BUFX2 BUFX2_insert1258 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_16_bF$buf9 )
);

BUFX2 BUFX2_insert1257 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_16_bF$buf10 )
);

BUFX2 BUFX2_insert1256 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_16_bF$buf11 )
);

BUFX2 BUFX2_insert1255 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_16_bF$buf12 )
);

BUFX2 BUFX2_insert1254 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_16_bF$buf13 )
);

BUFX2 BUFX2_insert1253 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_16_bF$buf14 )
);

BUFX2 BUFX2_insert1252 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_16_bF$buf15 )
);

BUFX2 BUFX2_insert1251 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_16_bF$buf16 )
);

BUFX2 BUFX2_insert1250 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_16_bF$buf17 )
);

BUFX2 BUFX2_insert1249 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_16_bF$buf18 )
);

BUFX2 BUFX2_insert1248 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_16_bF$buf19 )
);

BUFX2 BUFX2_insert1247 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_16_bF$buf20 )
);

BUFX2 BUFX2_insert1246 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_16_bF$buf21 )
);

BUFX2 BUFX2_insert1245 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_16_bF$buf22 )
);

BUFX2 BUFX2_insert1244 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_16_bF$buf23 )
);

BUFX2 BUFX2_insert1243 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_16_bF$buf24 )
);

BUFX2 BUFX2_insert1242 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_16_bF$buf25 )
);

BUFX2 BUFX2_insert1241 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_16_bF$buf26 )
);

BUFX2 BUFX2_insert1240 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_16_bF$buf27 )
);

BUFX2 BUFX2_insert1239 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_16_bF$buf28 )
);

BUFX2 BUFX2_insert1238 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_16_bF$buf29 )
);

BUFX2 BUFX2_insert1237 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_16_bF$buf30 )
);

BUFX2 BUFX2_insert1236 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_16_bF$buf31 )
);

BUFX2 BUFX2_insert1235 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_16_bF$buf32 )
);

BUFX2 BUFX2_insert1234 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_16_bF$buf33 )
);

BUFX2 BUFX2_insert1233 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_16_bF$buf34 )
);

BUFX2 BUFX2_insert1232 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_16_bF$buf35 )
);

BUFX2 BUFX2_insert1231 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_16_bF$buf36 )
);

BUFX2 BUFX2_insert1230 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_16_bF$buf37 )
);

BUFX2 BUFX2_insert1229 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_16_bF$buf38 )
);

BUFX2 BUFX2_insert1228 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_16_bF$buf39 )
);

BUFX2 BUFX2_insert1227 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_16_bF$buf40 )
);

BUFX2 BUFX2_insert1226 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_16_bF$buf41 )
);

BUFX2 BUFX2_insert1225 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_16_bF$buf42 )
);

BUFX2 BUFX2_insert1224 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_16_bF$buf43 )
);

BUFX2 BUFX2_insert1223 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_16_bF$buf44 )
);

BUFX2 BUFX2_insert1222 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_16_bF$buf45 )
);

BUFX2 BUFX2_insert1221 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9109_),
    .Y(_9109__bF$buf0)
);

BUFX2 BUFX2_insert1220 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9109_),
    .Y(_9109__bF$buf1)
);

BUFX2 BUFX2_insert1219 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9109_),
    .Y(_9109__bF$buf2)
);

BUFX2 BUFX2_insert1218 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9109_),
    .Y(_9109__bF$buf3)
);

BUFX2 BUFX2_insert1217 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9109_),
    .Y(_9109__bF$buf4)
);

BUFX2 BUFX2_insert1216 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9244_),
    .Y(_9244__bF$buf0)
);

BUFX2 BUFX2_insert1215 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9244_),
    .Y(_9244__bF$buf1)
);

BUFX2 BUFX2_insert1214 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9244_),
    .Y(_9244__bF$buf2)
);

BUFX2 BUFX2_insert1213 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9244_),
    .Y(_9244__bF$buf3)
);

BUFX2 BUFX2_insert1212 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9244_),
    .Y(_9244__bF$buf4)
);

BUFX2 BUFX2_insert1211 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546_),
    .Y(_5546__bF$buf0)
);

BUFX2 BUFX2_insert1210 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546_),
    .Y(_5546__bF$buf1)
);

BUFX2 BUFX2_insert1209 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546_),
    .Y(_5546__bF$buf2)
);

BUFX2 BUFX2_insert1208 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546_),
    .Y(_5546__bF$buf3)
);

BUFX2 BUFX2_insert1207 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546_),
    .Y(_5546__bF$buf4)
);

BUFX2 BUFX2_insert1206 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546_),
    .Y(_5546__bF$buf5)
);

BUFX2 BUFX2_insert1205 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546_),
    .Y(_5546__bF$buf6)
);

BUFX2 BUFX2_insert1204 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546_),
    .Y(_5546__bF$buf7)
);

BUFX2 BUFX2_insert1203 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546_),
    .Y(_5546__bF$buf8)
);

BUFX2 BUFX2_insert1202 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546_),
    .Y(_5546__bF$buf9)
);

BUFX2 BUFX2_insert1201 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546_),
    .Y(_5546__bF$buf10)
);

BUFX2 BUFX2_insert1200 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546_),
    .Y(_5546__bF$buf11)
);

BUFX2 BUFX2_insert1199 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546_),
    .Y(_5546__bF$buf12)
);

BUFX2 BUFX2_insert1198 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546_),
    .Y(_5546__bF$buf13)
);

BUFX2 BUFX2_insert1197 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546_),
    .Y(_5546__bF$buf14)
);

BUFX2 BUFX2_insert1196 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546_),
    .Y(_5546__bF$buf15)
);

BUFX2 BUFX2_insert1195 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490_),
    .Y(_5490__bF$buf0)
);

BUFX2 BUFX2_insert1194 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490_),
    .Y(_5490__bF$buf1)
);

BUFX2 BUFX2_insert1193 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490_),
    .Y(_5490__bF$buf2)
);

BUFX2 BUFX2_insert1192 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490_),
    .Y(_5490__bF$buf3)
);

BUFX2 BUFX2_insert1191 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490_),
    .Y(_5490__bF$buf4)
);

BUFX2 BUFX2_insert1190 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5681_),
    .Y(_5681__bF$buf0)
);

BUFX2 BUFX2_insert1189 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5681_),
    .Y(_5681__bF$buf1)
);

BUFX2 BUFX2_insert1188 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5681_),
    .Y(_5681__bF$buf2)
);

BUFX2 BUFX2_insert1187 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5681_),
    .Y(_5681__bF$buf3)
);

BUFX2 BUFX2_insert1186 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5681_),
    .Y(_5681__bF$buf4)
);

BUFX2 BUFX2_insert1185 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452_),
    .Y(_5452__bF$buf0)
);

BUFX2 BUFX2_insert1184 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452_),
    .Y(_5452__bF$buf1)
);

BUFX2 BUFX2_insert1183 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452_),
    .Y(_5452__bF$buf2)
);

BUFX2 BUFX2_insert1182 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452_),
    .Y(_5452__bF$buf3)
);

BUFX2 BUFX2_insert1181 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452_),
    .Y(_5452__bF$buf4)
);

BUFX2 BUFX2_insert1180 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[0]),
    .Y(_0__0_bF$buf0)
);

BUFX2 BUFX2_insert1179 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[0]),
    .Y(_0__0_bF$buf1)
);

BUFX2 BUFX2_insert1178 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[0]),
    .Y(_0__0_bF$buf2)
);

BUFX2 BUFX2_insert1177 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[0]),
    .Y(_0__0_bF$buf3)
);

BUFX2 BUFX2_insert1176 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[0]),
    .Y(_0__0_bF$buf4)
);

BUFX2 BUFX2_insert1175 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143_),
    .Y(_6143__bF$buf0)
);

BUFX2 BUFX2_insert1174 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143_),
    .Y(_6143__bF$buf1)
);

BUFX2 BUFX2_insert1173 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143_),
    .Y(_6143__bF$buf2)
);

BUFX2 BUFX2_insert1172 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143_),
    .Y(_6143__bF$buf3)
);

BUFX2 BUFX2_insert1171 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143_),
    .Y(_6143__bF$buf4)
);

BUFX2 BUFX2_insert1170 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2865_),
    .Y(_2865__bF$buf0)
);

BUFX2 BUFX2_insert1169 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2865_),
    .Y(_2865__bF$buf1)
);

BUFX2 BUFX2_insert1168 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2865_),
    .Y(_2865__bF$buf2)
);

BUFX2 BUFX2_insert1167 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2865_),
    .Y(_2865__bF$buf3)
);

BUFX2 BUFX2_insert1166 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1240_),
    .Y(_1240__bF$buf0)
);

BUFX2 BUFX2_insert1165 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1240_),
    .Y(_1240__bF$buf1)
);

BUFX2 BUFX2_insert1164 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1240_),
    .Y(_1240__bF$buf2)
);

BUFX2 BUFX2_insert1163 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1240_),
    .Y(_1240__bF$buf3)
);

BUFX2 BUFX2_insert1162 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1240_),
    .Y(_1240__bF$buf4)
);

BUFX2 BUFX2_insert1161 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [19]),
    .Y(\datapath.idinstr_19_bF$buf0 )
);

BUFX2 BUFX2_insert1160 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [19]),
    .Y(\datapath.idinstr_19_bF$buf1 )
);

BUFX2 BUFX2_insert1159 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [19]),
    .Y(\datapath.idinstr_19_bF$buf2 )
);

BUFX2 BUFX2_insert1158 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [19]),
    .Y(\datapath.idinstr_19_bF$buf3 )
);

BUFX2 BUFX2_insert1157 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [19]),
    .Y(\datapath.idinstr_19_bF$buf4 )
);

BUFX2 BUFX2_insert1156 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [19]),
    .Y(\datapath.idinstr_19_bF$buf5 )
);

BUFX2 BUFX2_insert1155 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_22_bF$buf0 )
);

BUFX2 BUFX2_insert1154 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_22_bF$buf1 )
);

BUFX2 BUFX2_insert1153 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_22_bF$buf2 )
);

BUFX2 BUFX2_insert1152 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_22_bF$buf3 )
);

BUFX2 BUFX2_insert1151 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_22_bF$buf4 )
);

BUFX2 BUFX2_insert1150 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_22_bF$buf5 )
);

BUFX2 BUFX2_insert1149 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_22_bF$buf6 )
);

BUFX2 BUFX2_insert1148 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_22_bF$buf7 )
);

BUFX2 BUFX2_insert1147 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_22_bF$buf8 )
);

BUFX2 BUFX2_insert1146 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_22_bF$buf9 )
);

BUFX2 BUFX2_insert1145 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_22_bF$buf10 )
);

BUFX2 BUFX2_insert1144 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_22_bF$buf11 )
);

BUFX2 BUFX2_insert1143 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_22_bF$buf12 )
);

BUFX2 BUFX2_insert1142 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_22_bF$buf13 )
);

BUFX2 BUFX2_insert1141 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_22_bF$buf14 )
);

BUFX2 BUFX2_insert1140 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_22_bF$buf15 )
);

BUFX2 BUFX2_insert1139 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_22_bF$buf16 )
);

BUFX2 BUFX2_insert1138 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_22_bF$buf17 )
);

BUFX2 BUFX2_insert1137 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_22_bF$buf18 )
);

BUFX2 BUFX2_insert1136 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_22_bF$buf19 )
);

BUFX2 BUFX2_insert1135 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_22_bF$buf20 )
);

BUFX2 BUFX2_insert1134 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_22_bF$buf21 )
);

BUFX2 BUFX2_insert1133 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_22_bF$buf22 )
);

BUFX2 BUFX2_insert1132 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_22_bF$buf23 )
);

BUFX2 BUFX2_insert1131 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_22_bF$buf24 )
);

BUFX2 BUFX2_insert1130 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_22_bF$buf25 )
);

BUFX2 BUFX2_insert1129 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_22_bF$buf26 )
);

BUFX2 BUFX2_insert1128 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_22_bF$buf27 )
);

BUFX2 BUFX2_insert1127 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_22_bF$buf28 )
);

BUFX2 BUFX2_insert1126 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_22_bF$buf29 )
);

BUFX2 BUFX2_insert1125 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_22_bF$buf30 )
);

BUFX2 BUFX2_insert1124 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_22_bF$buf31 )
);

BUFX2 BUFX2_insert1123 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_22_bF$buf32 )
);

BUFX2 BUFX2_insert1122 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_22_bF$buf33 )
);

BUFX2 BUFX2_insert1121 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_22_bF$buf34 )
);

BUFX2 BUFX2_insert1120 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_22_bF$buf35 )
);

BUFX2 BUFX2_insert1119 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_22_bF$buf36 )
);

BUFX2 BUFX2_insert1118 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_22_bF$buf37 )
);

BUFX2 BUFX2_insert1117 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_22_bF$buf38 )
);

BUFX2 BUFX2_insert1116 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_22_bF$buf39 )
);

BUFX2 BUFX2_insert1115 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_22_bF$buf40 )
);

BUFX2 BUFX2_insert1114 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_22_bF$buf41 )
);

BUFX2 BUFX2_insert1113 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_22_bF$buf42 )
);

BUFX2 BUFX2_insert1112 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_22_bF$buf43 )
);

BUFX2 BUFX2_insert1111 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall ),
    .Y(\datapath.pcstall_bF$buf0 )
);

BUFX2 BUFX2_insert1110 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall ),
    .Y(\datapath.pcstall_bF$buf1 )
);

BUFX2 BUFX2_insert1109 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall ),
    .Y(\datapath.pcstall_bF$buf2 )
);

BUFX2 BUFX2_insert1108 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall ),
    .Y(\datapath.pcstall_bF$buf3 )
);

BUFX2 BUFX2_insert1107 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall ),
    .Y(\datapath.pcstall_bF$buf4 )
);

BUFX2 BUFX2_insert1106 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall ),
    .Y(\datapath.pcstall_bF$buf5 )
);

BUFX2 BUFX2_insert1105 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall ),
    .Y(\datapath.pcstall_bF$buf6 )
);

BUFX2 BUFX2_insert1104 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall ),
    .Y(\datapath.pcstall_bF$buf7 )
);

BUFX2 BUFX2_insert1103 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2680_),
    .Y(_2680__bF$buf0)
);

BUFX2 BUFX2_insert1102 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2680_),
    .Y(_2680__bF$buf1)
);

BUFX2 BUFX2_insert1101 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2680_),
    .Y(_2680__bF$buf2)
);

BUFX2 BUFX2_insert1100 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2680_),
    .Y(_2680__bF$buf3)
);

BUFX2 BUFX2_insert1099 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret ),
    .Y(\datapath.regmret_bF$buf0 )
);

BUFX2 BUFX2_insert1098 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret ),
    .Y(\datapath.regmret_bF$buf1 )
);

BUFX2 BUFX2_insert1097 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret ),
    .Y(\datapath.regmret_bF$buf2 )
);

BUFX2 BUFX2_insert1096 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret ),
    .Y(\datapath.regmret_bF$buf3 )
);

BUFX2 BUFX2_insert1095 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret ),
    .Y(\datapath.regmret_bF$buf4 )
);

BUFX2 BUFX2_insert1094 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496_),
    .Y(_5496__bF$buf0)
);

BUFX2 BUFX2_insert1093 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496_),
    .Y(_5496__bF$buf1)
);

BUFX2 BUFX2_insert1092 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496_),
    .Y(_5496__bF$buf2)
);

BUFX2 BUFX2_insert1091 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496_),
    .Y(_5496__bF$buf3)
);

BUFX2 BUFX2_insert1090 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496_),
    .Y(_5496__bF$buf4)
);

BUFX2 BUFX2_insert1089 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458_),
    .Y(_5458__bF$buf0)
);

BUFX2 BUFX2_insert1088 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458_),
    .Y(_5458__bF$buf1)
);

BUFX2 BUFX2_insert1087 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458_),
    .Y(_5458__bF$buf2)
);

BUFX2 BUFX2_insert1086 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458_),
    .Y(_5458__bF$buf3)
);

BUFX2 BUFX2_insert1085 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458_),
    .Y(_5458__bF$buf4)
);

BUFX2 BUFX2_insert1084 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489_),
    .Y(_2489__bF$buf0)
);

BUFX2 BUFX2_insert1083 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489_),
    .Y(_2489__bF$buf1)
);

BUFX2 BUFX2_insert1082 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489_),
    .Y(_2489__bF$buf2)
);

BUFX2 BUFX2_insert1081 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489_),
    .Y(_2489__bF$buf3)
);

BUFX2 BUFX2_insert1080 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489_),
    .Y(_2489__bF$buf4)
);

BUFX2 BUFX2_insert1079 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489_),
    .Y(_2489__bF$buf5)
);

BUFX2 BUFX2_insert1078 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489_),
    .Y(_2489__bF$buf6)
);

BUFX2 BUFX2_insert1077 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489_),
    .Y(_2489__bF$buf7)
);

BUFX2 BUFX2_insert1076 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .Y(_254__bF$buf0)
);

BUFX2 BUFX2_insert1075 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .Y(_254__bF$buf1)
);

BUFX2 BUFX2_insert1074 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .Y(_254__bF$buf2)
);

BUFX2 BUFX2_insert1073 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .Y(_254__bF$buf3)
);

BUFX2 BUFX2_insert1072 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .Y(_254__bF$buf4)
);

BUFX2 BUFX2_insert1071 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614_),
    .Y(_5614__bF$buf0)
);

BUFX2 BUFX2_insert1070 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614_),
    .Y(_5614__bF$buf1)
);

BUFX2 BUFX2_insert1069 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614_),
    .Y(_5614__bF$buf2)
);

BUFX2 BUFX2_insert1068 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614_),
    .Y(_5614__bF$buf3)
);

BUFX2 BUFX2_insert1067 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614_),
    .Y(_5614__bF$buf4)
);

BUFX2 BUFX2_insert1066 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7607_),
    .Y(_7607__bF$buf0)
);

BUFX2 BUFX2_insert1065 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7607_),
    .Y(_7607__bF$buf1)
);

BUFX2 BUFX2_insert1064 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7607_),
    .Y(_7607__bF$buf2)
);

BUFX2 BUFX2_insert1063 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7607_),
    .Y(_7607__bF$buf3)
);

BUFX2 BUFX2_insert1062 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7607_),
    .Y(_7607__bF$buf4)
);

BUFX2 BUFX2_insert1061 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf0 )
);

BUFX2 BUFX2_insert1060 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf1 )
);

BUFX2 BUFX2_insert1059 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf2 )
);

BUFX2 BUFX2_insert1058 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf3 )
);

BUFX2 BUFX2_insert1057 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf4 )
);

BUFX2 BUFX2_insert1056 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf5 )
);

BUFX2 BUFX2_insert1055 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf6 )
);

BUFX2 BUFX2_insert1054 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf7 )
);

BUFX2 BUFX2_insert1053 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf8 )
);

BUFX2 BUFX2_insert1052 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf9 )
);

BUFX2 BUFX2_insert1051 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [0]),
    .Y(\datapath.alu.b_0_bF$buf10 )
);

BUFX2 BUFX2_insert1050 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610_),
    .Y(_7610__bF$buf0)
);

BUFX2 BUFX2_insert1049 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610_),
    .Y(_7610__bF$buf1)
);

BUFX2 BUFX2_insert1048 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610_),
    .Y(_7610__bF$buf2)
);

BUFX2 BUFX2_insert1047 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610_),
    .Y(_7610__bF$buf3)
);

BUFX2 BUFX2_insert1046 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610_),
    .Y(_7610__bF$buf4)
);

BUFX2 BUFX2_insert1045 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464_),
    .Y(_5464__bF$buf0)
);

BUFX2 BUFX2_insert1044 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464_),
    .Y(_5464__bF$buf1)
);

BUFX2 BUFX2_insert1043 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464_),
    .Y(_5464__bF$buf2)
);

BUFX2 BUFX2_insert1042 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464_),
    .Y(_5464__bF$buf3)
);

BUFX2 BUFX2_insert1041 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464_),
    .Y(_5464__bF$buf4)
);

BUFX2 BUFX2_insert1040 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_),
    .Y(_486__bF$buf0)
);

BUFX2 BUFX2_insert1039 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_),
    .Y(_486__bF$buf1)
);

BUFX2 BUFX2_insert1038 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_),
    .Y(_486__bF$buf2)
);

BUFX2 BUFX2_insert1037 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_),
    .Y(_486__bF$buf3)
);

BUFX2 BUFX2_insert1036 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_),
    .Y(_486__bF$buf4)
);

BUFX2 BUFX2_insert1035 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495_),
    .Y(_2495__bF$buf0)
);

BUFX2 BUFX2_insert1034 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495_),
    .Y(_2495__bF$buf1)
);

BUFX2 BUFX2_insert1033 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495_),
    .Y(_2495__bF$buf2)
);

BUFX2 BUFX2_insert1032 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495_),
    .Y(_2495__bF$buf3)
);

BUFX2 BUFX2_insert1031 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495_),
    .Y(_2495__bF$buf4)
);

BUFX2 BUFX2_insert1030 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495_),
    .Y(_2495__bF$buf5)
);

BUFX2 BUFX2_insert1029 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495_),
    .Y(_2495__bF$buf6)
);

BUFX2 BUFX2_insert1028 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_965_),
    .Y(_965__bF$buf0)
);

BUFX2 BUFX2_insert1027 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_965_),
    .Y(_965__bF$buf1)
);

BUFX2 BUFX2_insert1026 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_965_),
    .Y(_965__bF$buf2)
);

BUFX2 BUFX2_insert1025 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_965_),
    .Y(_965__bF$buf3)
);

BUFX2 BUFX2_insert1024 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_965_),
    .Y(_965__bF$buf4)
);

BUFX2 BUFX2_insert1023 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3339_),
    .Y(_3339__bF$buf0)
);

BUFX2 BUFX2_insert1022 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3339_),
    .Y(_3339__bF$buf1)
);

BUFX2 BUFX2_insert1021 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3339_),
    .Y(_3339__bF$buf2)
);

BUFX2 BUFX2_insert1020 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3339_),
    .Y(_3339__bF$buf3)
);

BUFX2 BUFX2_insert1019 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3339_),
    .Y(_3339__bF$buf4)
);

BUFX2 BUFX2_insert1018 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3339_),
    .Y(_3339__bF$buf5)
);

BUFX2 BUFX2_insert1017 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3339_),
    .Y(_3339__bF$buf6)
);

BUFX2 BUFX2_insert1016 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_604_),
    .Y(_604__bF$buf0)
);

BUFX2 BUFX2_insert1015 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_604_),
    .Y(_604__bF$buf1)
);

BUFX2 BUFX2_insert1014 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_604_),
    .Y(_604__bF$buf2)
);

BUFX2 BUFX2_insert1013 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_604_),
    .Y(_604__bF$buf3)
);

BUFX2 BUFX2_insert1012 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_604_),
    .Y(_604__bF$buf4)
);

BUFX2 BUFX2_insert1011 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [3]),
    .Y(\datapath.alu.b_3_bF$buf0 )
);

BUFX2 BUFX2_insert1010 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [3]),
    .Y(\datapath.alu.b_3_bF$buf1 )
);

BUFX2 BUFX2_insert1009 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [3]),
    .Y(\datapath.alu.b_3_bF$buf2 )
);

BUFX2 BUFX2_insert1008 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [3]),
    .Y(\datapath.alu.b_3_bF$buf3 )
);

BUFX2 BUFX2_insert1007 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [3]),
    .Y(\datapath.alu.b_3_bF$buf4 )
);

BUFX2 BUFX2_insert1006 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [3]),
    .Y(\datapath.alu.b_3_bF$buf5 )
);

BUFX2 BUFX2_insert1005 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [3]),
    .Y(\datapath.alu.b_3_bF$buf6 )
);

BUFX2 BUFX2_insert1004 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_298_),
    .Y(_298__bF$buf0)
);

BUFX2 BUFX2_insert1003 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_298_),
    .Y(_298__bF$buf1)
);

BUFX2 BUFX2_insert1002 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_298_),
    .Y(_298__bF$buf2)
);

BUFX2 BUFX2_insert1001 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_298_),
    .Y(_298__bF$buf3)
);

BUFX2 BUFX2_insert1000 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_298_),
    .Y(_298__bF$buf4)
);

BUFX2 BUFX2_insert999 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429_),
    .Y(_5429__bF$buf0)
);

BUFX2 BUFX2_insert998 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429_),
    .Y(_5429__bF$buf1)
);

BUFX2 BUFX2_insert997 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429_),
    .Y(_5429__bF$buf2)
);

BUFX2 BUFX2_insert996 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429_),
    .Y(_5429__bF$buf3)
);

BUFX2 BUFX2_insert995 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429_),
    .Y(_5429__bF$buf4)
);

BUFX2 BUFX2_insert994 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5793_),
    .Y(_5793__bF$buf0)
);

BUFX2 BUFX2_insert993 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5793_),
    .Y(_5793__bF$buf1)
);

BUFX2 BUFX2_insert992 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5793_),
    .Y(_5793__bF$buf2)
);

BUFX2 BUFX2_insert991 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5793_),
    .Y(_5793__bF$buf3)
);

BUFX2 BUFX2_insert990 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5793_),
    .Y(_5793__bF$buf4)
);

BUFX2 BUFX2_insert989 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470_),
    .Y(_5470__bF$buf0)
);

BUFX2 BUFX2_insert988 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470_),
    .Y(_5470__bF$buf1)
);

BUFX2 BUFX2_insert987 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470_),
    .Y(_5470__bF$buf2)
);

BUFX2 BUFX2_insert986 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470_),
    .Y(_5470__bF$buf3)
);

BUFX2 BUFX2_insert985 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470_),
    .Y(_5470__bF$buf4)
);

BUFX2 BUFX2_insert984 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432_),
    .Y(_5432__bF$buf0)
);

BUFX2 BUFX2_insert983 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432_),
    .Y(_5432__bF$buf1)
);

BUFX2 BUFX2_insert982 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432_),
    .Y(_5432__bF$buf2)
);

BUFX2 BUFX2_insert981 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432_),
    .Y(_5432__bF$buf3)
);

BUFX2 BUFX2_insert980 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432_),
    .Y(_5432__bF$buf4)
);

BUFX2 BUFX2_insert979 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432_),
    .Y(_5432__bF$buf5)
);

BUFX2 BUFX2_insert978 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432_),
    .Y(_5432__bF$buf6)
);

BUFX2 BUFX2_insert977 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432_),
    .Y(_5432__bF$buf7)
);

BUFX2 BUFX2_insert976 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432_),
    .Y(_5432__bF$buf8)
);

BUFX2 BUFX2_insert975 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432_),
    .Y(_5432__bF$buf9)
);

BUFX2 BUFX2_insert974 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432_),
    .Y(_5432__bF$buf10)
);

BUFX2 BUFX2_insert973 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893_),
    .Y(_5893__bF$buf0)
);

BUFX2 BUFX2_insert972 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893_),
    .Y(_5893__bF$buf1)
);

BUFX2 BUFX2_insert971 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893_),
    .Y(_5893__bF$buf2)
);

BUFX2 BUFX2_insert970 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893_),
    .Y(_5893__bF$buf3)
);

BUFX2 BUFX2_insert969 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893_),
    .Y(_5893__bF$buf4)
);

BUFX2 BUFX2_insert968 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_495_),
    .Y(_495__bF$buf0)
);

BUFX2 BUFX2_insert967 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_495_),
    .Y(_495__bF$buf1)
);

BUFX2 BUFX2_insert966 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_495_),
    .Y(_495__bF$buf2)
);

BUFX2 BUFX2_insert965 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_495_),
    .Y(_495__bF$buf3)
);

BUFX2 BUFX2_insert964 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_495_),
    .Y(_495__bF$buf4)
);

CLKBUF1 CLKBUF1_insert963 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf0)
);

CLKBUF1 CLKBUF1_insert962 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf1)
);

CLKBUF1 CLKBUF1_insert961 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf2)
);

CLKBUF1 CLKBUF1_insert960 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf3)
);

CLKBUF1 CLKBUF1_insert959 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf4)
);

CLKBUF1 CLKBUF1_insert958 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf5)
);

CLKBUF1 CLKBUF1_insert957 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf6)
);

CLKBUF1 CLKBUF1_insert956 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf7)
);

CLKBUF1 CLKBUF1_insert955 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf8)
);

CLKBUF1 CLKBUF1_insert954 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf9)
);

CLKBUF1 CLKBUF1_insert953 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf10)
);

CLKBUF1 CLKBUF1_insert952 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf11)
);

CLKBUF1 CLKBUF1_insert951 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf12)
);

CLKBUF1 CLKBUF1_insert950 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf13)
);

CLKBUF1 CLKBUF1_insert949 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf14)
);

CLKBUF1 CLKBUF1_insert948 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf15)
);

CLKBUF1 CLKBUF1_insert947 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf16)
);

CLKBUF1 CLKBUF1_insert946 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf17)
);

CLKBUF1 CLKBUF1_insert945 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf18)
);

CLKBUF1 CLKBUF1_insert944 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf19)
);

CLKBUF1 CLKBUF1_insert943 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf20)
);

CLKBUF1 CLKBUF1_insert942 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf21)
);

CLKBUF1 CLKBUF1_insert941 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf22)
);

CLKBUF1 CLKBUF1_insert940 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf23)
);

CLKBUF1 CLKBUF1_insert939 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf24)
);

CLKBUF1 CLKBUF1_insert938 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf25)
);

CLKBUF1 CLKBUF1_insert937 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf26)
);

CLKBUF1 CLKBUF1_insert936 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf27)
);

CLKBUF1 CLKBUF1_insert935 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf28)
);

CLKBUF1 CLKBUF1_insert934 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf29)
);

CLKBUF1 CLKBUF1_insert933 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf30)
);

CLKBUF1 CLKBUF1_insert932 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf31)
);

CLKBUF1 CLKBUF1_insert931 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf32)
);

CLKBUF1 CLKBUF1_insert930 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf33)
);

CLKBUF1 CLKBUF1_insert929 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf34)
);

CLKBUF1 CLKBUF1_insert928 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf35)
);

CLKBUF1 CLKBUF1_insert927 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf36)
);

CLKBUF1 CLKBUF1_insert926 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf37)
);

CLKBUF1 CLKBUF1_insert925 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf38)
);

CLKBUF1 CLKBUF1_insert924 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf39)
);

CLKBUF1 CLKBUF1_insert923 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf40)
);

CLKBUF1 CLKBUF1_insert922 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf41)
);

CLKBUF1 CLKBUF1_insert921 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf42)
);

CLKBUF1 CLKBUF1_insert920 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf43)
);

CLKBUF1 CLKBUF1_insert919 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf44)
);

CLKBUF1 CLKBUF1_insert918 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf45)
);

CLKBUF1 CLKBUF1_insert917 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf46)
);

CLKBUF1 CLKBUF1_insert916 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf47)
);

CLKBUF1 CLKBUF1_insert915 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf48)
);

CLKBUF1 CLKBUF1_insert914 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf49)
);

CLKBUF1 CLKBUF1_insert913 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf50)
);

CLKBUF1 CLKBUF1_insert912 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf51)
);

CLKBUF1 CLKBUF1_insert911 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf52)
);

CLKBUF1 CLKBUF1_insert910 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf53)
);

CLKBUF1 CLKBUF1_insert909 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf54)
);

CLKBUF1 CLKBUF1_insert908 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf55)
);

CLKBUF1 CLKBUF1_insert907 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf56)
);

CLKBUF1 CLKBUF1_insert906 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf57)
);

CLKBUF1 CLKBUF1_insert905 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf58)
);

CLKBUF1 CLKBUF1_insert904 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf59)
);

CLKBUF1 CLKBUF1_insert903 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf60)
);

CLKBUF1 CLKBUF1_insert902 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf61)
);

CLKBUF1 CLKBUF1_insert901 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf62)
);

CLKBUF1 CLKBUF1_insert900 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf63)
);

CLKBUF1 CLKBUF1_insert899 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf64)
);

CLKBUF1 CLKBUF1_insert898 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf65)
);

CLKBUF1 CLKBUF1_insert897 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf66)
);

CLKBUF1 CLKBUF1_insert896 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf67)
);

CLKBUF1 CLKBUF1_insert895 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf68)
);

CLKBUF1 CLKBUF1_insert894 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf69)
);

CLKBUF1 CLKBUF1_insert893 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf70)
);

CLKBUF1 CLKBUF1_insert892 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf71)
);

CLKBUF1 CLKBUF1_insert891 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf72)
);

CLKBUF1 CLKBUF1_insert890 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf73)
);

CLKBUF1 CLKBUF1_insert889 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf74)
);

CLKBUF1 CLKBUF1_insert888 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf75)
);

CLKBUF1 CLKBUF1_insert887 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf76)
);

CLKBUF1 CLKBUF1_insert886 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf77)
);

CLKBUF1 CLKBUF1_insert885 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf78)
);

CLKBUF1 CLKBUF1_insert884 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf79)
);

CLKBUF1 CLKBUF1_insert883 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf80)
);

CLKBUF1 CLKBUF1_insert882 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf81)
);

CLKBUF1 CLKBUF1_insert881 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf82)
);

CLKBUF1 CLKBUF1_insert880 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf83)
);

CLKBUF1 CLKBUF1_insert879 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf84)
);

CLKBUF1 CLKBUF1_insert878 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf85)
);

CLKBUF1 CLKBUF1_insert877 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf86)
);

CLKBUF1 CLKBUF1_insert876 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf87)
);

CLKBUF1 CLKBUF1_insert875 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf88)
);

CLKBUF1 CLKBUF1_insert874 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf89)
);

CLKBUF1 CLKBUF1_insert873 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf90)
);

CLKBUF1 CLKBUF1_insert872 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf91)
);

CLKBUF1 CLKBUF1_insert871 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf92)
);

CLKBUF1 CLKBUF1_insert870 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf93)
);

CLKBUF1 CLKBUF1_insert869 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf94)
);

CLKBUF1 CLKBUF1_insert868 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf95)
);

CLKBUF1 CLKBUF1_insert867 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf96)
);

CLKBUF1 CLKBUF1_insert866 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf97)
);

CLKBUF1 CLKBUF1_insert865 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf98)
);

CLKBUF1 CLKBUF1_insert864 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf99)
);

CLKBUF1 CLKBUF1_insert863 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf100)
);

CLKBUF1 CLKBUF1_insert862 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf101)
);

CLKBUF1 CLKBUF1_insert861 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf102)
);

CLKBUF1 CLKBUF1_insert860 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf103)
);

CLKBUF1 CLKBUF1_insert859 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf104)
);

CLKBUF1 CLKBUF1_insert858 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf105)
);

CLKBUF1 CLKBUF1_insert857 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf106)
);

CLKBUF1 CLKBUF1_insert856 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf107)
);

CLKBUF1 CLKBUF1_insert855 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf108)
);

CLKBUF1 CLKBUF1_insert854 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf109)
);

CLKBUF1 CLKBUF1_insert853 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf110)
);

CLKBUF1 CLKBUF1_insert852 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf111)
);

CLKBUF1 CLKBUF1_insert851 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf112)
);

CLKBUF1 CLKBUF1_insert850 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf113)
);

CLKBUF1 CLKBUF1_insert849 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf114)
);

CLKBUF1 CLKBUF1_insert848 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf115)
);

CLKBUF1 CLKBUF1_insert847 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf116)
);

CLKBUF1 CLKBUF1_insert846 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf117)
);

CLKBUF1 CLKBUF1_insert845 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf118)
);

CLKBUF1 CLKBUF1_insert844 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf119)
);

CLKBUF1 CLKBUF1_insert843 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf120)
);

CLKBUF1 CLKBUF1_insert842 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf121)
);

CLKBUF1 CLKBUF1_insert841 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf122)
);

CLKBUF1 CLKBUF1_insert840 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf123)
);

CLKBUF1 CLKBUF1_insert839 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf124)
);

CLKBUF1 CLKBUF1_insert838 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf125)
);

CLKBUF1 CLKBUF1_insert837 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf126)
);

CLKBUF1 CLKBUF1_insert836 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf127)
);

CLKBUF1 CLKBUF1_insert835 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf128)
);

CLKBUF1 CLKBUF1_insert834 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf129)
);

CLKBUF1 CLKBUF1_insert833 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf130)
);

CLKBUF1 CLKBUF1_insert832 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf131)
);

CLKBUF1 CLKBUF1_insert831 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf132)
);

CLKBUF1 CLKBUF1_insert830 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf133)
);

CLKBUF1 CLKBUF1_insert829 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf134)
);

CLKBUF1 CLKBUF1_insert828 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf135)
);

CLKBUF1 CLKBUF1_insert827 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf136)
);

CLKBUF1 CLKBUF1_insert826 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf137)
);

CLKBUF1 CLKBUF1_insert825 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf138)
);

CLKBUF1 CLKBUF1_insert824 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf139)
);

CLKBUF1 CLKBUF1_insert823 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf140)
);

CLKBUF1 CLKBUF1_insert822 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf141)
);

CLKBUF1 CLKBUF1_insert821 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf1),
    .Y(CLK_bF$buf142)
);

CLKBUF1 CLKBUF1_insert820 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf0),
    .Y(CLK_bF$buf143)
);

CLKBUF1 CLKBUF1_insert819 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf11),
    .Y(CLK_bF$buf144)
);

CLKBUF1 CLKBUF1_insert818 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf10),
    .Y(CLK_bF$buf145)
);

CLKBUF1 CLKBUF1_insert817 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf9),
    .Y(CLK_bF$buf146)
);

CLKBUF1 CLKBUF1_insert816 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf8),
    .Y(CLK_bF$buf147)
);

CLKBUF1 CLKBUF1_insert815 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf7),
    .Y(CLK_bF$buf148)
);

CLKBUF1 CLKBUF1_insert814 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf6),
    .Y(CLK_bF$buf149)
);

CLKBUF1 CLKBUF1_insert813 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf5),
    .Y(CLK_bF$buf150)
);

CLKBUF1 CLKBUF1_insert812 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf4),
    .Y(CLK_bF$buf151)
);

CLKBUF1 CLKBUF1_insert811 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf3),
    .Y(CLK_bF$buf152)
);

CLKBUF1 CLKBUF1_insert810 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CLK_hier0_bF$buf2),
    .Y(CLK_bF$buf153)
);

BUFX2 BUFX2_insert809 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_974_),
    .Y(_974__bF$buf0)
);

BUFX2 BUFX2_insert808 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_974_),
    .Y(_974__bF$buf1)
);

BUFX2 BUFX2_insert807 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_974_),
    .Y(_974__bF$buf2)
);

BUFX2 BUFX2_insert806 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_974_),
    .Y(_974__bF$buf3)
);

BUFX2 BUFX2_insert805 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_974_),
    .Y(_974__bF$buf4)
);

BUFX2 BUFX2_insert804 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476_),
    .Y(_5476__bF$buf0)
);

BUFX2 BUFX2_insert803 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476_),
    .Y(_5476__bF$buf1)
);

BUFX2 BUFX2_insert802 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476_),
    .Y(_5476__bF$buf2)
);

BUFX2 BUFX2_insert801 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476_),
    .Y(_5476__bF$buf3)
);

BUFX2 BUFX2_insert800 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476_),
    .Y(_5476__bF$buf4)
);

BUFX2 BUFX2_insert799 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .Y(_498__bF$buf0)
);

BUFX2 BUFX2_insert798 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .Y(_498__bF$buf1)
);

BUFX2 BUFX2_insert797 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .Y(_498__bF$buf2)
);

BUFX2 BUFX2_insert796 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .Y(_498__bF$buf3)
);

BUFX2 BUFX2_insert795 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .Y(_498__bF$buf4)
);

BUFX2 BUFX2_insert794 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438_),
    .Y(_5438__bF$buf0)
);

BUFX2 BUFX2_insert793 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438_),
    .Y(_5438__bF$buf1)
);

BUFX2 BUFX2_insert792 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438_),
    .Y(_5438__bF$buf2)
);

BUFX2 BUFX2_insert791 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438_),
    .Y(_5438__bF$buf3)
);

BUFX2 BUFX2_insert790 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438_),
    .Y(_5438__bF$buf4)
);

BUFX2 BUFX2_insert789 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5993_),
    .Y(_5993__bF$buf0)
);

BUFX2 BUFX2_insert788 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5993_),
    .Y(_5993__bF$buf1)
);

BUFX2 BUFX2_insert787 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5993_),
    .Y(_5993__bF$buf2)
);

BUFX2 BUFX2_insert786 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5993_),
    .Y(_5993__bF$buf3)
);

BUFX2 BUFX2_insert785 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5993_),
    .Y(_5993__bF$buf4)
);

BUFX2 BUFX2_insert784 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5993_),
    .Y(_5993__bF$buf5)
);

BUFX2 BUFX2_insert783 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5993_),
    .Y(_5993__bF$buf6)
);

BUFX2 BUFX2_insert782 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5993_),
    .Y(_5993__bF$buf7)
);

BUFX2 BUFX2_insert781 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_595_),
    .Y(_595__bF$buf0)
);

BUFX2 BUFX2_insert780 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_595_),
    .Y(_595__bF$buf1)
);

BUFX2 BUFX2_insert779 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_595_),
    .Y(_595__bF$buf2)
);

BUFX2 BUFX2_insert778 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_595_),
    .Y(_595__bF$buf3)
);

BUFX2 BUFX2_insert777 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_595_),
    .Y(_595__bF$buf4)
);

BUFX2 BUFX2_insert776 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_977_),
    .Y(_977__bF$buf0)
);

BUFX2 BUFX2_insert775 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_977_),
    .Y(_977__bF$buf1)
);

BUFX2 BUFX2_insert774 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_977_),
    .Y(_977__bF$buf2)
);

BUFX2 BUFX2_insert773 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_977_),
    .Y(_977__bF$buf3)
);

BUFX2 BUFX2_insert772 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_977_),
    .Y(_977__bF$buf4)
);

BUFX2 BUFX2_insert771 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3448_),
    .Y(_3448__bF$buf0)
);

BUFX2 BUFX2_insert770 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3448_),
    .Y(_3448__bF$buf1)
);

BUFX2 BUFX2_insert769 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3448_),
    .Y(_3448__bF$buf2)
);

BUFX2 BUFX2_insert768 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3448_),
    .Y(_3448__bF$buf3)
);

BUFX2 BUFX2_insert767 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3448_),
    .Y(_3448__bF$buf4)
);

BUFX2 BUFX2_insert766 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482_),
    .Y(_5482__bF$buf0)
);

BUFX2 BUFX2_insert765 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482_),
    .Y(_5482__bF$buf1)
);

BUFX2 BUFX2_insert764 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482_),
    .Y(_5482__bF$buf2)
);

BUFX2 BUFX2_insert763 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482_),
    .Y(_5482__bF$buf3)
);

BUFX2 BUFX2_insert762 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482_),
    .Y(_5482__bF$buf4)
);

BUFX2 BUFX2_insert761 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9142_),
    .Y(_9142__bF$buf0)
);

BUFX2 BUFX2_insert760 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9142_),
    .Y(_9142__bF$buf1)
);

BUFX2 BUFX2_insert759 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9142_),
    .Y(_9142__bF$buf2)
);

BUFX2 BUFX2_insert758 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9142_),
    .Y(_9142__bF$buf3)
);

BUFX2 BUFX2_insert757 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9142_),
    .Y(_9142__bF$buf4)
);

BUFX2 BUFX2_insert756 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444_),
    .Y(_5444__bF$buf0)
);

BUFX2 BUFX2_insert755 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444_),
    .Y(_5444__bF$buf1)
);

BUFX2 BUFX2_insert754 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444_),
    .Y(_5444__bF$buf2)
);

BUFX2 BUFX2_insert753 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444_),
    .Y(_5444__bF$buf3)
);

BUFX2 BUFX2_insert752 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444_),
    .Y(_5444__bF$buf4)
);

BUFX2 BUFX2_insert751 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5826_),
    .Y(_5826__bF$buf0)
);

BUFX2 BUFX2_insert750 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5826_),
    .Y(_5826__bF$buf1)
);

BUFX2 BUFX2_insert749 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5826_),
    .Y(_5826__bF$buf2)
);

BUFX2 BUFX2_insert748 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5826_),
    .Y(_5826__bF$buf3)
);

BUFX2 BUFX2_insert747 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5826_),
    .Y(_5826__bF$buf4)
);

BUFX2 BUFX2_insert746 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041_),
    .Y(_6041__bF$buf0)
);

BUFX2 BUFX2_insert745 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041_),
    .Y(_6041__bF$buf1)
);

BUFX2 BUFX2_insert744 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041_),
    .Y(_6041__bF$buf2)
);

BUFX2 BUFX2_insert743 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041_),
    .Y(_6041__bF$buf3)
);

BUFX2 BUFX2_insert742 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041_),
    .Y(_6041__bF$buf4)
);

BUFX2 BUFX2_insert741 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041_),
    .Y(_6041__bF$buf5)
);

BUFX2 BUFX2_insert740 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041_),
    .Y(_6041__bF$buf6)
);

BUFX2 BUFX2_insert739 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041_),
    .Y(_6041__bF$buf7)
);

BUFX2 BUFX2_insert738 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041_),
    .Y(_6041__bF$buf8)
);

BUFX2 BUFX2_insert737 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9277_),
    .Y(_9277__bF$buf0)
);

BUFX2 BUFX2_insert736 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9277_),
    .Y(_9277__bF$buf1)
);

BUFX2 BUFX2_insert735 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9277_),
    .Y(_9277__bF$buf2)
);

BUFX2 BUFX2_insert734 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9277_),
    .Y(_9277__bF$buf3)
);

BUFX2 BUFX2_insert733 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9277_),
    .Y(_9277__bF$buf4)
);

BUFX2 BUFX2_insert732 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579_),
    .Y(_5579__bF$buf0)
);

BUFX2 BUFX2_insert731 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579_),
    .Y(_5579__bF$buf1)
);

BUFX2 BUFX2_insert730 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579_),
    .Y(_5579__bF$buf2)
);

BUFX2 BUFX2_insert729 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579_),
    .Y(_5579__bF$buf3)
);

BUFX2 BUFX2_insert728 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579_),
    .Y(_5579__bF$buf4)
);

BUFX2 BUFX2_insert727 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579_),
    .Y(_5579__bF$buf5)
);

BUFX2 BUFX2_insert726 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450_),
    .Y(_5450__bF$buf0)
);

BUFX2 BUFX2_insert725 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450_),
    .Y(_5450__bF$buf1)
);

BUFX2 BUFX2_insert724 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450_),
    .Y(_5450__bF$buf2)
);

BUFX2 BUFX2_insert723 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450_),
    .Y(_5450__bF$buf3)
);

BUFX2 BUFX2_insert722 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450_),
    .Y(_5450__bF$buf4)
);

BUFX2 BUFX2_insert721 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141_),
    .Y(_6141__bF$buf0)
);

BUFX2 BUFX2_insert720 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141_),
    .Y(_6141__bF$buf1)
);

BUFX2 BUFX2_insert719 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141_),
    .Y(_6141__bF$buf2)
);

BUFX2 BUFX2_insert718 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141_),
    .Y(_6141__bF$buf3)
);

BUFX2 BUFX2_insert717 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141_),
    .Y(_6141__bF$buf4)
);

BUFX2 BUFX2_insert716 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141_),
    .Y(_6141__bF$buf5)
);

BUFX2 BUFX2_insert715 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141_),
    .Y(_6141__bF$buf6)
);

BUFX2 BUFX2_insert714 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141_),
    .Y(_6141__bF$buf7)
);

BUFX2 BUFX2_insert713 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141_),
    .Y(_6141__bF$buf8)
);

BUFX2 BUFX2_insert712 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141_),
    .Y(_6141__bF$buf9)
);

BUFX2 BUFX2_insert711 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141_),
    .Y(_6141__bF$buf10)
);

BUFX2 BUFX2_insert710 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9377_),
    .Y(_9377__bF$buf0)
);

BUFX2 BUFX2_insert709 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9377_),
    .Y(_9377__bF$buf1)
);

BUFX2 BUFX2_insert708 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9377_),
    .Y(_9377__bF$buf2)
);

BUFX2 BUFX2_insert707 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9377_),
    .Y(_9377__bF$buf3)
);

BUFX2 BUFX2_insert706 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9377_),
    .Y(_9377__bF$buf4)
);

BUFX2 BUFX2_insert705 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_17_bF$buf0 )
);

BUFX2 BUFX2_insert704 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_17_bF$buf1 )
);

BUFX2 BUFX2_insert703 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_17_bF$buf2 )
);

BUFX2 BUFX2_insert702 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_17_bF$buf3 )
);

BUFX2 BUFX2_insert701 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_17_bF$buf4 )
);

BUFX2 BUFX2_insert700 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_17_bF$buf5 )
);

BUFX2 BUFX2_insert699 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_17_bF$buf6 )
);

BUFX2 BUFX2_insert698 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_17_bF$buf7 )
);

BUFX2 BUFX2_insert697 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_17_bF$buf8 )
);

BUFX2 BUFX2_insert696 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_17_bF$buf9 )
);

BUFX2 BUFX2_insert695 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_17_bF$buf10 )
);

BUFX2 BUFX2_insert694 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_17_bF$buf11 )
);

BUFX2 BUFX2_insert693 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_17_bF$buf12 )
);

BUFX2 BUFX2_insert692 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_17_bF$buf13 )
);

BUFX2 BUFX2_insert691 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_17_bF$buf14 )
);

BUFX2 BUFX2_insert690 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_17_bF$buf15 )
);

BUFX2 BUFX2_insert689 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_17_bF$buf16 )
);

BUFX2 BUFX2_insert688 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_17_bF$buf17 )
);

BUFX2 BUFX2_insert687 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_17_bF$buf18 )
);

BUFX2 BUFX2_insert686 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_17_bF$buf19 )
);

BUFX2 BUFX2_insert685 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_17_bF$buf20 )
);

BUFX2 BUFX2_insert684 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_17_bF$buf21 )
);

BUFX2 BUFX2_insert683 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_17_bF$buf22 )
);

BUFX2 BUFX2_insert682 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_17_bF$buf23 )
);

BUFX2 BUFX2_insert681 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_17_bF$buf24 )
);

BUFX2 BUFX2_insert680 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_17_bF$buf25 )
);

BUFX2 BUFX2_insert679 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_17_bF$buf26 )
);

BUFX2 BUFX2_insert678 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_17_bF$buf27 )
);

BUFX2 BUFX2_insert677 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_17_bF$buf28 )
);

BUFX2 BUFX2_insert676 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_17_bF$buf29 )
);

BUFX2 BUFX2_insert675 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_17_bF$buf30 )
);

BUFX2 BUFX2_insert674 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_17_bF$buf31 )
);

BUFX2 BUFX2_insert673 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_17_bF$buf32 )
);

BUFX2 BUFX2_insert672 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_17_bF$buf33 )
);

BUFX2 BUFX2_insert671 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_17_bF$buf34 )
);

BUFX2 BUFX2_insert670 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_17_bF$buf35 )
);

BUFX2 BUFX2_insert669 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_17_bF$buf36 )
);

BUFX2 BUFX2_insert668 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_17_bF$buf37 )
);

BUFX2 BUFX2_insert667 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_17_bF$buf38 )
);

BUFX2 BUFX2_insert666 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_17_bF$buf39 )
);

BUFX2 BUFX2_insert665 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_17_bF$buf40 )
);

BUFX2 BUFX2_insert664 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_17_bF$buf41 )
);

BUFX2 BUFX2_insert663 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488_),
    .Y(_5488__bF$buf0)
);

BUFX2 BUFX2_insert662 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488_),
    .Y(_5488__bF$buf1)
);

BUFX2 BUFX2_insert661 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488_),
    .Y(_5488__bF$buf2)
);

BUFX2 BUFX2_insert660 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488_),
    .Y(_5488__bF$buf3)
);

BUFX2 BUFX2_insert659 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488_),
    .Y(_5488__bF$buf4)
);

BUFX2 BUFX2_insert658 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_20_bF$buf0 )
);

BUFX2 BUFX2_insert657 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_20_bF$buf1 )
);

BUFX2 BUFX2_insert656 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_20_bF$buf2 )
);

BUFX2 BUFX2_insert655 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_20_bF$buf3 )
);

BUFX2 BUFX2_insert654 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_20_bF$buf4 )
);

BUFX2 BUFX2_insert653 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_20_bF$buf5 )
);

BUFX2 BUFX2_insert652 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_20_bF$buf6 )
);

BUFX2 BUFX2_insert651 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_20_bF$buf7 )
);

BUFX2 BUFX2_insert650 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_20_bF$buf8 )
);

BUFX2 BUFX2_insert649 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_20_bF$buf9 )
);

BUFX2 BUFX2_insert648 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_20_bF$buf10 )
);

BUFX2 BUFX2_insert647 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_20_bF$buf11 )
);

BUFX2 BUFX2_insert646 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_20_bF$buf12 )
);

BUFX2 BUFX2_insert645 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_20_bF$buf13 )
);

BUFX2 BUFX2_insert644 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_20_bF$buf14 )
);

BUFX2 BUFX2_insert643 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_20_bF$buf15 )
);

BUFX2 BUFX2_insert642 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_20_bF$buf16 )
);

BUFX2 BUFX2_insert641 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_20_bF$buf17 )
);

BUFX2 BUFX2_insert640 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_20_bF$buf18 )
);

BUFX2 BUFX2_insert639 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_20_bF$buf19 )
);

BUFX2 BUFX2_insert638 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_20_bF$buf20 )
);

BUFX2 BUFX2_insert637 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_20_bF$buf21 )
);

BUFX2 BUFX2_insert636 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_20_bF$buf22 )
);

BUFX2 BUFX2_insert635 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_20_bF$buf23 )
);

BUFX2 BUFX2_insert634 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_20_bF$buf24 )
);

BUFX2 BUFX2_insert633 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_20_bF$buf25 )
);

BUFX2 BUFX2_insert632 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_20_bF$buf26 )
);

BUFX2 BUFX2_insert631 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_20_bF$buf27 )
);

BUFX2 BUFX2_insert630 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_20_bF$buf28 )
);

BUFX2 BUFX2_insert629 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_20_bF$buf29 )
);

BUFX2 BUFX2_insert628 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_20_bF$buf30 )
);

BUFX2 BUFX2_insert627 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_20_bF$buf31 )
);

BUFX2 BUFX2_insert626 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_20_bF$buf32 )
);

BUFX2 BUFX2_insert625 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_20_bF$buf33 )
);

BUFX2 BUFX2_insert624 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_20_bF$buf34 )
);

BUFX2 BUFX2_insert623 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_20_bF$buf35 )
);

BUFX2 BUFX2_insert622 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_20_bF$buf36 )
);

BUFX2 BUFX2_insert621 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_20_bF$buf37 )
);

BUFX2 BUFX2_insert620 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_20_bF$buf38 )
);

BUFX2 BUFX2_insert619 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_20_bF$buf39 )
);

BUFX2 BUFX2_insert618 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_20_bF$buf40 )
);

BUFX2 BUFX2_insert617 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_20_bF$buf41 )
);

BUFX2 BUFX2_insert616 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_20_bF$buf42 )
);

BUFX2 BUFX2_insert615 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_20_bF$buf43 )
);

BUFX2 BUFX2_insert614 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_20_bF$buf44 )
);

BUFX2 BUFX2_insert613 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_20_bF$buf45 )
);

BUFX2 BUFX2_insert612 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_20_bF$buf46 )
);

BUFX2 BUFX2_insert611 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_20_bF$buf47 )
);

BUFX2 BUFX2_insert610 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_20_bF$buf48 )
);

BUFX2 BUFX2_insert609 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_20_bF$buf49 )
);

BUFX2 BUFX2_insert608 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_20_bF$buf50 )
);

BUFX2 BUFX2_insert607 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_20_bF$buf51 )
);

BUFX2 BUFX2_insert606 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_20_bF$buf52 )
);

BUFX2 BUFX2_insert605 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_20_bF$buf53 )
);

BUFX2 BUFX2_insert604 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_20_bF$buf54 )
);

BUFX2 BUFX2_insert603 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_20_bF$buf55 )
);

BUFX2 BUFX2_insert602 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1238_),
    .Y(_1238__bF$buf0)
);

BUFX2 BUFX2_insert601 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1238_),
    .Y(_1238__bF$buf1)
);

BUFX2 BUFX2_insert600 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1238_),
    .Y(_1238__bF$buf2)
);

BUFX2 BUFX2_insert599 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1238_),
    .Y(_1238__bF$buf3)
);

BUFX2 BUFX2_insert598 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1238_),
    .Y(_1238__bF$buf4)
);

BUFX2 BUFX2_insert597 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5509_),
    .Y(_5509__bF$buf0)
);

BUFX2 BUFX2_insert596 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5509_),
    .Y(_5509__bF$buf1)
);

BUFX2 BUFX2_insert595 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5509_),
    .Y(_5509__bF$buf2)
);

BUFX2 BUFX2_insert594 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5509_),
    .Y(_5509__bF$buf3)
);

BUFX2 BUFX2_insert593 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5509_),
    .Y(_5509__bF$buf4)
);

BUFX2 BUFX2_insert592 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[1]),
    .Y(_0__1_bF$buf0)
);

BUFX2 BUFX2_insert591 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[1]),
    .Y(_0__1_bF$buf1)
);

BUFX2 BUFX2_insert590 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[1]),
    .Y(_0__1_bF$buf2)
);

BUFX2 BUFX2_insert589 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[1]),
    .Y(_0__1_bF$buf3)
);

BUFX2 BUFX2_insert588 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[1]),
    .Y(_0__1_bF$buf4)
);

BUFX2 BUFX2_insert587 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[1]),
    .Y(_0__1_bF$buf5)
);

BUFX2 BUFX2_insert586 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[1]),
    .Y(_0__1_bF$buf6)
);

BUFX2 BUFX2_insert585 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[1]),
    .Y(_0__1_bF$buf7)
);

BUFX2 BUFX2_insert584 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[1]),
    .Y(_0__1_bF$buf8)
);

BUFX2 BUFX2_insert583 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[1]),
    .Y(_0__1_bF$buf9)
);

BUFX2 BUFX2_insert582 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144_),
    .Y(_6144__bF$buf0)
);

BUFX2 BUFX2_insert581 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144_),
    .Y(_6144__bF$buf1)
);

BUFX2 BUFX2_insert580 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144_),
    .Y(_6144__bF$buf2)
);

BUFX2 BUFX2_insert579 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144_),
    .Y(_6144__bF$buf3)
);

BUFX2 BUFX2_insert578 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144_),
    .Y(_6144__bF$buf4)
);

BUFX2 BUFX2_insert577 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144_),
    .Y(_6144__bF$buf5)
);

BUFX2 BUFX2_insert576 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144_),
    .Y(_6144__bF$buf6)
);

BUFX2 BUFX2_insert575 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144_),
    .Y(_6144__bF$buf7)
);

BUFX2 BUFX2_insert574 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144_),
    .Y(_6144__bF$buf8)
);

BUFX2 BUFX2_insert573 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144_),
    .Y(_6144__bF$buf9)
);

BUFX2 BUFX2_insert572 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144_),
    .Y(_6144__bF$buf10)
);

BUFX2 BUFX2_insert571 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210_),
    .Y(_9210__bF$buf0)
);

BUFX2 BUFX2_insert570 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210_),
    .Y(_9210__bF$buf1)
);

BUFX2 BUFX2_insert569 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210_),
    .Y(_9210__bF$buf2)
);

BUFX2 BUFX2_insert568 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210_),
    .Y(_9210__bF$buf3)
);

BUFX2 BUFX2_insert567 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210_),
    .Y(_9210__bF$buf4)
);

BUFX2 BUFX2_insert566 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463_),
    .Y(_3463__bF$buf0)
);

BUFX2 BUFX2_insert565 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463_),
    .Y(_3463__bF$buf1)
);

BUFX2 BUFX2_insert564 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463_),
    .Y(_3463__bF$buf2)
);

BUFX2 BUFX2_insert563 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463_),
    .Y(_3463__bF$buf3)
);

BUFX2 BUFX2_insert562 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463_),
    .Y(_3463__bF$buf4)
);

BUFX2 BUFX2_insert561 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463_),
    .Y(_3463__bF$buf5)
);

BUFX2 BUFX2_insert560 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463_),
    .Y(_3463__bF$buf6)
);

BUFX2 BUFX2_insert559 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192_),
    .Y(_4192__bF$buf0)
);

BUFX2 BUFX2_insert558 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192_),
    .Y(_4192__bF$buf1)
);

BUFX2 BUFX2_insert557 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192_),
    .Y(_4192__bF$buf2)
);

BUFX2 BUFX2_insert556 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192_),
    .Y(_4192__bF$buf3)
);

BUFX2 BUFX2_insert555 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192_),
    .Y(_4192__bF$buf4)
);

BUFX2 BUFX2_insert554 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [23]),
    .Y(\datapath.idinstr_23_bF$buf0 )
);

BUFX2 BUFX2_insert553 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [23]),
    .Y(\datapath.idinstr_23_bF$buf1 )
);

BUFX2 BUFX2_insert552 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [23]),
    .Y(\datapath.idinstr_23_bF$buf2 )
);

BUFX2 BUFX2_insert551 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [23]),
    .Y(\datapath.idinstr_23_bF$buf3 )
);

BUFX2 BUFX2_insert550 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [23]),
    .Y(\datapath.idinstr_23_bF$buf4 )
);

BUFX2 BUFX2_insert549 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [23]),
    .Y(\datapath.idinstr_23_bF$buf5 )
);

BUFX2 BUFX2_insert548 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [23]),
    .Y(\datapath.idinstr_23_bF$buf6 )
);

BUFX2 BUFX2_insert547 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [23]),
    .Y(\datapath.idinstr_23_bF$buf7 )
);

BUFX2 BUFX2_insert546 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494_),
    .Y(_5494__bF$buf0)
);

BUFX2 BUFX2_insert545 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494_),
    .Y(_5494__bF$buf1)
);

BUFX2 BUFX2_insert544 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494_),
    .Y(_5494__bF$buf2)
);

BUFX2 BUFX2_insert543 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494_),
    .Y(_5494__bF$buf3)
);

BUFX2 BUFX2_insert542 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494_),
    .Y(_5494__bF$buf4)
);

BUFX2 BUFX2_insert541 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060_),
    .Y(_4060__bF$buf0)
);

BUFX2 BUFX2_insert540 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060_),
    .Y(_4060__bF$buf1)
);

BUFX2 BUFX2_insert539 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060_),
    .Y(_4060__bF$buf2)
);

BUFX2 BUFX2_insert538 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060_),
    .Y(_4060__bF$buf3)
);

BUFX2 BUFX2_insert537 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456_),
    .Y(_5456__bF$buf0)
);

BUFX2 BUFX2_insert536 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456_),
    .Y(_5456__bF$buf1)
);

BUFX2 BUFX2_insert535 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456_),
    .Y(_5456__bF$buf2)
);

BUFX2 BUFX2_insert534 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456_),
    .Y(_5456__bF$buf3)
);

BUFX2 BUFX2_insert533 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456_),
    .Y(_5456__bF$buf4)
);

BUFX2 BUFX2_insert532 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6147_),
    .Y(_6147__bF$buf0)
);

BUFX2 BUFX2_insert531 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6147_),
    .Y(_6147__bF$buf1)
);

BUFX2 BUFX2_insert530 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6147_),
    .Y(_6147__bF$buf2)
);

BUFX2 BUFX2_insert529 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6147_),
    .Y(_6147__bF$buf3)
);

BUFX2 BUFX2_insert528 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6147_),
    .Y(_6147__bF$buf4)
);

BUFX2 BUFX2_insert527 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2869_),
    .Y(_2869__bF$buf0)
);

BUFX2 BUFX2_insert526 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2869_),
    .Y(_2869__bF$buf1)
);

BUFX2 BUFX2_insert525 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2869_),
    .Y(_2869__bF$buf2)
);

BUFX2 BUFX2_insert524 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2869_),
    .Y(_2869__bF$buf3)
);

BUFX2 BUFX2_insert523 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9310_),
    .Y(_9310__bF$buf0)
);

BUFX2 BUFX2_insert522 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9310_),
    .Y(_9310__bF$buf1)
);

BUFX2 BUFX2_insert521 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9310_),
    .Y(_9310__bF$buf2)
);

BUFX2 BUFX2_insert520 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9310_),
    .Y(_9310__bF$buf3)
);

BUFX2 BUFX2_insert519 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9310_),
    .Y(_9310__bF$buf4)
);

BUFX2 BUFX2_insert518 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9310_),
    .Y(_9310__bF$buf5)
);

BUFX2 BUFX2_insert517 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9310_),
    .Y(_9310__bF$buf6)
);

BUFX2 BUFX2_insert516 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9310_),
    .Y(_9310__bF$buf7)
);

BUFX2 BUFX2_insert515 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462_),
    .Y(_5462__bF$buf0)
);

BUFX2 BUFX2_insert514 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462_),
    .Y(_5462__bF$buf1)
);

BUFX2 BUFX2_insert513 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462_),
    .Y(_5462__bF$buf2)
);

BUFX2 BUFX2_insert512 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462_),
    .Y(_5462__bF$buf3)
);

BUFX2 BUFX2_insert511 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462_),
    .Y(_5462__bF$buf4)
);

BUFX2 BUFX2_insert510 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615_),
    .Y(_5615__bF$buf0)
);

BUFX2 BUFX2_insert509 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615_),
    .Y(_5615__bF$buf1)
);

BUFX2 BUFX2_insert508 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615_),
    .Y(_5615__bF$buf2)
);

BUFX2 BUFX2_insert507 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615_),
    .Y(_5615__bF$buf3)
);

BUFX2 BUFX2_insert506 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615_),
    .Y(_5615__bF$buf4)
);

BUFX2 BUFX2_insert505 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615_),
    .Y(_5615__bF$buf5)
);

BUFX2 BUFX2_insert504 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615_),
    .Y(_5615__bF$buf6)
);

BUFX2 BUFX2_insert503 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615_),
    .Y(_5615__bF$buf7)
);

BUFX2 BUFX2_insert502 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615_),
    .Y(_5615__bF$buf8)
);

BUFX2 BUFX2_insert501 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4198_),
    .Y(_4198__bF$buf0)
);

BUFX2 BUFX2_insert500 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4198_),
    .Y(_4198__bF$buf1)
);

BUFX2 BUFX2_insert499 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4198_),
    .Y(_4198__bF$buf2)
);

BUFX2 BUFX2_insert498 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4198_),
    .Y(_4198__bF$buf3)
);

BUFX2 BUFX2_insert497 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4198_),
    .Y(_4198__bF$buf4)
);

BUFX2 BUFX2_insert496 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9410_),
    .Y(_9410__bF$buf0)
);

BUFX2 BUFX2_insert495 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9410_),
    .Y(_9410__bF$buf1)
);

BUFX2 BUFX2_insert494 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9410_),
    .Y(_9410__bF$buf2)
);

BUFX2 BUFX2_insert493 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9410_),
    .Y(_9410__bF$buf3)
);

BUFX2 BUFX2_insert492 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9410_),
    .Y(_9410__bF$buf4)
);

BUFX2 BUFX2_insert491 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_963_),
    .Y(_963__bF$buf0)
);

BUFX2 BUFX2_insert490 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_963_),
    .Y(_963__bF$buf1)
);

BUFX2 BUFX2_insert489 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_963_),
    .Y(_963__bF$buf2)
);

BUFX2 BUFX2_insert488 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_963_),
    .Y(_963__bF$buf3)
);

BUFX2 BUFX2_insert487 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_963_),
    .Y(_963__bF$buf4)
);

BUFX2 BUFX2_insert486 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608_),
    .Y(_7608__bF$buf0)
);

BUFX2 BUFX2_insert485 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608_),
    .Y(_7608__bF$buf1)
);

BUFX2 BUFX2_insert484 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608_),
    .Y(_7608__bF$buf2)
);

BUFX2 BUFX2_insert483 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608_),
    .Y(_7608__bF$buf3)
);

BUFX2 BUFX2_insert482 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608_),
    .Y(_7608__bF$buf4)
);

BUFX2 BUFX2_insert481 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608_),
    .Y(_7608__bF$buf5)
);

BUFX2 BUFX2_insert480 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608_),
    .Y(_7608__bF$buf6)
);

BUFX2 BUFX2_insert479 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608_),
    .Y(_7608__bF$buf7)
);

BUFX2 BUFX2_insert478 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608_),
    .Y(_7608__bF$buf8)
);

BUFX2 BUFX2_insert477 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608_),
    .Y(_7608__bF$buf9)
);

BUFX2 BUFX2_insert476 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608_),
    .Y(_7608__bF$buf10)
);

BUFX2 BUFX2_insert475 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [1]),
    .Y(\datapath.alu.b_1_bF$buf0 )
);

BUFX2 BUFX2_insert474 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [1]),
    .Y(\datapath.alu.b_1_bF$buf1 )
);

BUFX2 BUFX2_insert473 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [1]),
    .Y(\datapath.alu.b_1_bF$buf2 )
);

BUFX2 BUFX2_insert472 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [1]),
    .Y(\datapath.alu.b_1_bF$buf3 )
);

BUFX2 BUFX2_insert471 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [1]),
    .Y(\datapath.alu.b_1_bF$buf4 )
);

BUFX2 BUFX2_insert470 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [1]),
    .Y(\datapath.alu.b_1_bF$buf5 )
);

BUFX2 BUFX2_insert469 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [1]),
    .Y(\datapath.alu.b_1_bF$buf6 )
);

BUFX2 BUFX2_insert468 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611_),
    .Y(_7611__bF$buf0)
);

BUFX2 BUFX2_insert467 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611_),
    .Y(_7611__bF$buf1)
);

BUFX2 BUFX2_insert466 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611_),
    .Y(_7611__bF$buf2)
);

BUFX2 BUFX2_insert465 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611_),
    .Y(_7611__bF$buf3)
);

BUFX2 BUFX2_insert464 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611_),
    .Y(_7611__bF$buf4)
);

BUFX2 BUFX2_insert463 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611_),
    .Y(_7611__bF$buf5)
);

BUFX2 BUFX2_insert462 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611_),
    .Y(_7611__bF$buf6)
);

BUFX2 BUFX2_insert461 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611_),
    .Y(_7611__bF$buf7)
);

BUFX2 BUFX2_insert460 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611_),
    .Y(_7611__bF$buf8)
);

BUFX2 BUFX2_insert459 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611_),
    .Y(_7611__bF$buf9)
);

BUFX2 BUFX2_insert458 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611_),
    .Y(_7611__bF$buf10)
);

BUFX2 BUFX2_insert457 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3798_),
    .Y(_3798__bF$buf0)
);

BUFX2 BUFX2_insert456 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3798_),
    .Y(_3798__bF$buf1)
);

BUFX2 BUFX2_insert455 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3798_),
    .Y(_3798__bF$buf2)
);

BUFX2 BUFX2_insert454 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3798_),
    .Y(_3798__bF$buf3)
);

BUFX2 BUFX2_insert453 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3798_),
    .Y(_3798__bF$buf4)
);

BUFX2 BUFX2_insert452 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5715_),
    .Y(_5715__bF$buf0)
);

BUFX2 BUFX2_insert451 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5715_),
    .Y(_5715__bF$buf1)
);

BUFX2 BUFX2_insert450 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5715_),
    .Y(_5715__bF$buf2)
);

BUFX2 BUFX2_insert449 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5715_),
    .Y(_5715__bF$buf3)
);

BUFX2 BUFX2_insert448 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5715_),
    .Y(_5715__bF$buf4)
);

BUFX2 BUFX2_insert447 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5715_),
    .Y(_5715__bF$buf5)
);

BUFX2 BUFX2_insert446 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5715_),
    .Y(_5715__bF$buf6)
);

BUFX2 BUFX2_insert445 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5715_),
    .Y(_5715__bF$buf7)
);

BUFX2 BUFX2_insert444 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_490_),
    .Y(_490__bF$buf0)
);

BUFX2 BUFX2_insert443 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_490_),
    .Y(_490__bF$buf1)
);

BUFX2 BUFX2_insert442 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_490_),
    .Y(_490__bF$buf2)
);

BUFX2 BUFX2_insert441 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_490_),
    .Y(_490__bF$buf3)
);

BUFX2 BUFX2_insert440 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_490_),
    .Y(_490__bF$buf4)
);

BUFX2 BUFX2_insert439 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2708_),
    .Y(_2708__bF$buf0)
);

BUFX2 BUFX2_insert438 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2708_),
    .Y(_2708__bF$buf1)
);

BUFX2 BUFX2_insert437 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2708_),
    .Y(_2708__bF$buf2)
);

BUFX2 BUFX2_insert436 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2708_),
    .Y(_2708__bF$buf3)
);

BUFX2 BUFX2_insert435 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [4]),
    .Y(\datapath.alu.b_4_bF$buf0 )
);

BUFX2 BUFX2_insert434 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [4]),
    .Y(\datapath.alu.b_4_bF$buf1 )
);

BUFX2 BUFX2_insert433 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [4]),
    .Y(\datapath.alu.b_4_bF$buf2 )
);

BUFX2 BUFX2_insert432 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [4]),
    .Y(\datapath.alu.b_4_bF$buf3 )
);

BUFX2 BUFX2_insert431 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [4]),
    .Y(\datapath.alu.b_4_bF$buf4 )
);

BUFX2 BUFX2_insert430 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7614_),
    .Y(_7614__bF$buf0)
);

BUFX2 BUFX2_insert429 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7614_),
    .Y(_7614__bF$buf1)
);

BUFX2 BUFX2_insert428 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7614_),
    .Y(_7614__bF$buf2)
);

BUFX2 BUFX2_insert427 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7614_),
    .Y(_7614__bF$buf3)
);

BUFX2 BUFX2_insert426 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7614_),
    .Y(_7614__bF$buf4)
);

BUFX2 BUFX2_insert425 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468_),
    .Y(_5468__bF$buf0)
);

BUFX2 BUFX2_insert424 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468_),
    .Y(_5468__bF$buf1)
);

BUFX2 BUFX2_insert423 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468_),
    .Y(_5468__bF$buf2)
);

BUFX2 BUFX2_insert422 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468_),
    .Y(_5468__bF$buf3)
);

BUFX2 BUFX2_insert421 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468_),
    .Y(_5468__bF$buf4)
);

BUFX2 BUFX2_insert420 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075_),
    .Y(_9075__bF$buf0)
);

BUFX2 BUFX2_insert419 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075_),
    .Y(_9075__bF$buf1)
);

BUFX2 BUFX2_insert418 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075_),
    .Y(_9075__bF$buf2)
);

BUFX2 BUFX2_insert417 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075_),
    .Y(_9075__bF$buf3)
);

BUFX2 BUFX2_insert416 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075_),
    .Y(_9075__bF$buf4)
);

BUFX2 BUFX2_insert415 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .Y(_611__bF$buf0)
);

BUFX2 BUFX2_insert414 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .Y(_611__bF$buf1)
);

BUFX2 BUFX2_insert413 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .Y(_611__bF$buf2)
);

BUFX2 BUFX2_insert412 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .Y(_611__bF$buf3)
);

BUFX2 BUFX2_insert411 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .Y(_611__bF$buf4)
);

BUFX2 BUFX2_insert410 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759_),
    .Y(_5759__bF$buf0)
);

BUFX2 BUFX2_insert409 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759_),
    .Y(_5759__bF$buf1)
);

BUFX2 BUFX2_insert408 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759_),
    .Y(_5759__bF$buf2)
);

BUFX2 BUFX2_insert407 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759_),
    .Y(_5759__bF$buf3)
);

BUFX2 BUFX2_insert406 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759_),
    .Y(_5759__bF$buf4)
);

BUFX2 BUFX2_insert405 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474_),
    .Y(_5474__bF$buf0)
);

BUFX2 BUFX2_insert404 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474_),
    .Y(_5474__bF$buf1)
);

BUFX2 BUFX2_insert403 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474_),
    .Y(_5474__bF$buf2)
);

BUFX2 BUFX2_insert402 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474_),
    .Y(_5474__bF$buf3)
);

BUFX2 BUFX2_insert401 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474_),
    .Y(_5474__bF$buf4)
);

BUFX2 BUFX2_insert400 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894_),
    .Y(_5894__bF$buf0)
);

BUFX2 BUFX2_insert399 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894_),
    .Y(_5894__bF$buf1)
);

BUFX2 BUFX2_insert398 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894_),
    .Y(_5894__bF$buf2)
);

BUFX2 BUFX2_insert397 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894_),
    .Y(_5894__bF$buf3)
);

BUFX2 BUFX2_insert396 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894_),
    .Y(_5894__bF$buf4)
);

BUFX2 BUFX2_insert395 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894_),
    .Y(_5894__bF$buf5)
);

BUFX2 BUFX2_insert394 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894_),
    .Y(_5894__bF$buf6)
);

BUFX2 BUFX2_insert393 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894_),
    .Y(_5894__bF$buf7)
);

BUFX2 BUFX2_insert392 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894_),
    .Y(_5894__bF$buf8)
);

BUFX2 BUFX2_insert391 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436_),
    .Y(_5436__bF$buf0)
);

BUFX2 BUFX2_insert390 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436_),
    .Y(_5436__bF$buf1)
);

BUFX2 BUFX2_insert389 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436_),
    .Y(_5436__bF$buf2)
);

BUFX2 BUFX2_insert388 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436_),
    .Y(_5436__bF$buf3)
);

BUFX2 BUFX2_insert387 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436_),
    .Y(_5436__bF$buf4)
);

BUFX2 BUFX2_insert386 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3675_),
    .Y(_3675__bF$buf0)
);

BUFX2 BUFX2_insert385 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3675_),
    .Y(_3675__bF$buf1)
);

BUFX2 BUFX2_insert384 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3675_),
    .Y(_3675__bF$buf2)
);

BUFX2 BUFX2_insert383 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3675_),
    .Y(_3675__bF$buf3)
);

BUFX2 BUFX2_insert382 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3675_),
    .Y(_3675__bF$buf4)
);

BUFX2 BUFX2_insert381 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_614_),
    .Y(_614__bF$buf0)
);

BUFX2 BUFX2_insert380 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_614_),
    .Y(_614__bF$buf1)
);

BUFX2 BUFX2_insert379 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_614_),
    .Y(_614__bF$buf2)
);

BUFX2 BUFX2_insert378 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_614_),
    .Y(_614__bF$buf3)
);

BUFX2 BUFX2_insert377 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_614_),
    .Y(_614__bF$buf4)
);

BUFX2 BUFX2_insert376 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9175_),
    .Y(_9175__bF$buf0)
);

BUFX2 BUFX2_insert375 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9175_),
    .Y(_9175__bF$buf1)
);

BUFX2 BUFX2_insert374 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9175_),
    .Y(_9175__bF$buf2)
);

BUFX2 BUFX2_insert373 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9175_),
    .Y(_9175__bF$buf3)
);

BUFX2 BUFX2_insert372 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9175_),
    .Y(_9175__bF$buf4)
);

BUFX2 BUFX2_insert371 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9175_),
    .Y(_9175__bF$buf5)
);

BUFX2 BUFX2_insert370 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9175_),
    .Y(_9175__bF$buf6)
);

BUFX2 BUFX2_insert369 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9175_),
    .Y(_9175__bF$buf7)
);

BUFX2 BUFX2_insert368 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5859_),
    .Y(_5859__bF$buf0)
);

BUFX2 BUFX2_insert367 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5859_),
    .Y(_5859__bF$buf1)
);

BUFX2 BUFX2_insert366 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5859_),
    .Y(_5859__bF$buf2)
);

BUFX2 BUFX2_insert365 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5859_),
    .Y(_5859__bF$buf3)
);

BUFX2 BUFX2_insert364 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5859_),
    .Y(_5859__bF$buf4)
);

BUFX2 BUFX2_insert363 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5859_),
    .Y(_5859__bF$buf5)
);

BUFX2 BUFX2_insert362 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5859_),
    .Y(_5859__bF$buf6)
);

BUFX2 BUFX2_insert361 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5859_),
    .Y(_5859__bF$buf7)
);

BUFX2 BUFX2_insert360 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_596_),
    .Y(_596__bF$buf0)
);

BUFX2 BUFX2_insert359 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_596_),
    .Y(_596__bF$buf1)
);

BUFX2 BUFX2_insert358 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_596_),
    .Y(_596__bF$buf2)
);

BUFX2 BUFX2_insert357 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_596_),
    .Y(_596__bF$buf3)
);

BUFX2 BUFX2_insert356 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_596_),
    .Y(_596__bF$buf4)
);

BUFX2 BUFX2_insert355 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6074_),
    .Y(_6074__bF$buf0)
);

BUFX2 BUFX2_insert354 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6074_),
    .Y(_6074__bF$buf1)
);

BUFX2 BUFX2_insert353 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6074_),
    .Y(_6074__bF$buf2)
);

BUFX2 BUFX2_insert352 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6074_),
    .Y(_6074__bF$buf3)
);

BUFX2 BUFX2_insert351 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6074_),
    .Y(_6074__bF$buf4)
);

BUFX2 BUFX2_insert350 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480_),
    .Y(_5480__bF$buf0)
);

BUFX2 BUFX2_insert349 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480_),
    .Y(_5480__bF$buf1)
);

BUFX2 BUFX2_insert348 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480_),
    .Y(_5480__bF$buf2)
);

BUFX2 BUFX2_insert347 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480_),
    .Y(_5480__bF$buf3)
);

BUFX2 BUFX2_insert346 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480_),
    .Y(_5480__bF$buf4)
);

BUFX2 BUFX2_insert345 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442_),
    .Y(_5442__bF$buf0)
);

BUFX2 BUFX2_insert344 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442_),
    .Y(_5442__bF$buf1)
);

BUFX2 BUFX2_insert343 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442_),
    .Y(_5442__bF$buf2)
);

BUFX2 BUFX2_insert342 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442_),
    .Y(_5442__bF$buf3)
);

BUFX2 BUFX2_insert341 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442_),
    .Y(_5442__bF$buf4)
);

BUFX2 BUFX2_insert340 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_617_),
    .Y(_617__bF$buf0)
);

BUFX2 BUFX2_insert339 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_617_),
    .Y(_617__bF$buf1)
);

BUFX2 BUFX2_insert338 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_617_),
    .Y(_617__bF$buf2)
);

BUFX2 BUFX2_insert337 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_617_),
    .Y(_617__bF$buf3)
);

BUFX2 BUFX2_insert336 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_617_),
    .Y(_617__bF$buf4)
);

BUFX2 BUFX2_insert335 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall ),
    .Y(\bypassandflushunit.stall_bF$buf0 )
);

BUFX2 BUFX2_insert334 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall ),
    .Y(\bypassandflushunit.stall_bF$buf1 )
);

BUFX2 BUFX2_insert333 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall ),
    .Y(\bypassandflushunit.stall_bF$buf2 )
);

BUFX2 BUFX2_insert332 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall ),
    .Y(\bypassandflushunit.stall_bF$buf3 )
);

BUFX2 BUFX2_insert331 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall ),
    .Y(\bypassandflushunit.stall_bF$buf4 )
);

BUFX2 BUFX2_insert330 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall ),
    .Y(\bypassandflushunit.stall_bF$buf5 )
);

BUFX2 BUFX2_insert329 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall ),
    .Y(\bypassandflushunit.stall_bF$buf6 )
);

BUFX2 BUFX2_insert328 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall ),
    .Y(\bypassandflushunit.stall_bF$buf7 )
);

BUFX2 BUFX2_insert327 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall ),
    .Y(\bypassandflushunit.stall_bF$buf8 )
);

BUFX2 BUFX2_insert326 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall ),
    .Y(\bypassandflushunit.stall_bF$buf9 )
);

BUFX2 BUFX2_insert325 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4008_),
    .Y(_4008__bF$buf0)
);

BUFX2 BUFX2_insert324 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4008_),
    .Y(_4008__bF$buf1)
);

BUFX2 BUFX2_insert323 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4008_),
    .Y(_4008__bF$buf2)
);

BUFX2 BUFX2_insert322 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4008_),
    .Y(_4008__bF$buf3)
);

BUFX2 BUFX2_insert321 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2799_),
    .Y(_2799__bF$buf0)
);

BUFX2 BUFX2_insert320 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2799_),
    .Y(_2799__bF$buf1)
);

BUFX2 BUFX2_insert319 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2799_),
    .Y(_2799__bF$buf2)
);

BUFX2 BUFX2_insert318 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2799_),
    .Y(_2799__bF$buf3)
);

BUFX2 BUFX2_insert317 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580_),
    .Y(_5580__bF$buf0)
);

BUFX2 BUFX2_insert316 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580_),
    .Y(_5580__bF$buf1)
);

BUFX2 BUFX2_insert315 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580_),
    .Y(_5580__bF$buf2)
);

BUFX2 BUFX2_insert314 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580_),
    .Y(_5580__bF$buf3)
);

BUFX2 BUFX2_insert313 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580_),
    .Y(_5580__bF$buf4)
);

BUFX2 BUFX2_insert312 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_15_bF$buf0 )
);

BUFX2 BUFX2_insert311 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_15_bF$buf1 )
);

BUFX2 BUFX2_insert310 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_15_bF$buf2 )
);

BUFX2 BUFX2_insert309 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_15_bF$buf3 )
);

BUFX2 BUFX2_insert308 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_15_bF$buf4 )
);

BUFX2 BUFX2_insert307 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_15_bF$buf5 )
);

BUFX2 BUFX2_insert306 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_15_bF$buf6 )
);

BUFX2 BUFX2_insert305 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_15_bF$buf7 )
);

BUFX2 BUFX2_insert304 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_15_bF$buf8 )
);

BUFX2 BUFX2_insert303 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_15_bF$buf9 )
);

BUFX2 BUFX2_insert302 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_15_bF$buf10 )
);

BUFX2 BUFX2_insert301 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_15_bF$buf11 )
);

BUFX2 BUFX2_insert300 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_15_bF$buf12 )
);

BUFX2 BUFX2_insert299 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_15_bF$buf13 )
);

BUFX2 BUFX2_insert298 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_15_bF$buf14 )
);

BUFX2 BUFX2_insert297 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_15_bF$buf15 )
);

BUFX2 BUFX2_insert296 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_15_bF$buf16 )
);

BUFX2 BUFX2_insert295 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_15_bF$buf17 )
);

BUFX2 BUFX2_insert294 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_15_bF$buf18 )
);

BUFX2 BUFX2_insert293 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_15_bF$buf19 )
);

BUFX2 BUFX2_insert292 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_15_bF$buf20 )
);

BUFX2 BUFX2_insert291 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_15_bF$buf21 )
);

BUFX2 BUFX2_insert290 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_15_bF$buf22 )
);

BUFX2 BUFX2_insert289 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_15_bF$buf23 )
);

BUFX2 BUFX2_insert288 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_15_bF$buf24 )
);

BUFX2 BUFX2_insert287 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_15_bF$buf25 )
);

BUFX2 BUFX2_insert286 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_15_bF$buf26 )
);

BUFX2 BUFX2_insert285 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_15_bF$buf27 )
);

BUFX2 BUFX2_insert284 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_15_bF$buf28 )
);

BUFX2 BUFX2_insert283 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_15_bF$buf29 )
);

BUFX2 BUFX2_insert282 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_15_bF$buf30 )
);

BUFX2 BUFX2_insert281 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_15_bF$buf31 )
);

BUFX2 BUFX2_insert280 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_15_bF$buf32 )
);

BUFX2 BUFX2_insert279 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_15_bF$buf33 )
);

BUFX2 BUFX2_insert278 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_15_bF$buf34 )
);

BUFX2 BUFX2_insert277 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_15_bF$buf35 )
);

BUFX2 BUFX2_insert276 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_15_bF$buf36 )
);

BUFX2 BUFX2_insert275 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_15_bF$buf37 )
);

BUFX2 BUFX2_insert274 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_15_bF$buf38 )
);

BUFX2 BUFX2_insert273 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_15_bF$buf39 )
);

BUFX2 BUFX2_insert272 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_15_bF$buf40 )
);

BUFX2 BUFX2_insert271 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_15_bF$buf41 )
);

BUFX2 BUFX2_insert270 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_15_bF$buf42 )
);

BUFX2 BUFX2_insert269 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_15_bF$buf43 )
);

BUFX2 BUFX2_insert268 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_15_bF$buf44 )
);

BUFX2 BUFX2_insert267 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_15_bF$buf45 )
);

BUFX2 BUFX2_insert266 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_15_bF$buf46 )
);

BUFX2 BUFX2_insert265 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_15_bF$buf47 )
);

BUFX2 BUFX2_insert264 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_15_bF$buf48 )
);

BUFX2 BUFX2_insert263 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf6 ),
    .Y(\datapath.idinstr_15_bF$buf49 )
);

BUFX2 BUFX2_insert262 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_15_bF$buf50 )
);

BUFX2 BUFX2_insert261 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_15_bF$buf51 )
);

BUFX2 BUFX2_insert260 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_15_bF$buf52 )
);

BUFX2 BUFX2_insert259 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_15_bF$buf53 )
);

BUFX2 BUFX2_insert258 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486_),
    .Y(_5486__bF$buf0)
);

BUFX2 BUFX2_insert257 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486_),
    .Y(_5486__bF$buf1)
);

BUFX2 BUFX2_insert256 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486_),
    .Y(_5486__bF$buf2)
);

BUFX2 BUFX2_insert255 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486_),
    .Y(_5486__bF$buf3)
);

BUFX2 BUFX2_insert254 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486_),
    .Y(_5486__bF$buf4)
);

BUFX2 BUFX2_insert253 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448_),
    .Y(_5448__bF$buf0)
);

BUFX2 BUFX2_insert252 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448_),
    .Y(_5448__bF$buf1)
);

BUFX2 BUFX2_insert251 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448_),
    .Y(_5448__bF$buf2)
);

BUFX2 BUFX2_insert250 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448_),
    .Y(_5448__bF$buf3)
);

BUFX2 BUFX2_insert249 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448_),
    .Y(_5448__bF$buf4)
);

BUFX2 BUFX2_insert248 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545_),
    .Y(_5545__bF$buf0)
);

BUFX2 BUFX2_insert247 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545_),
    .Y(_5545__bF$buf1)
);

BUFX2 BUFX2_insert246 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545_),
    .Y(_5545__bF$buf2)
);

BUFX2 BUFX2_insert245 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545_),
    .Y(_5545__bF$buf3)
);

BUFX2 BUFX2_insert244 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545_),
    .Y(_5545__bF$buf4)
);

BUFX2 BUFX2_insert243 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802_),
    .Y(_3802__bF$buf0)
);

BUFX2 BUFX2_insert242 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802_),
    .Y(_3802__bF$buf1)
);

BUFX2 BUFX2_insert241 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802_),
    .Y(_3802__bF$buf2)
);

BUFX2 BUFX2_insert240 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802_),
    .Y(_3802__bF$buf3)
);

BUFX2 BUFX2_insert239 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802_),
    .Y(_3802__bF$buf4)
);

BUFX2 BUFX2_insert238 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802_),
    .Y(_3802__bF$buf5)
);

BUFX2 BUFX2_insert237 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802_),
    .Y(_3802__bF$buf6)
);

BUFX2 BUFX2_insert236 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236_),
    .Y(_1236__bF$buf0)
);

BUFX2 BUFX2_insert235 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236_),
    .Y(_1236__bF$buf1)
);

BUFX2 BUFX2_insert234 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236_),
    .Y(_1236__bF$buf2)
);

BUFX2 BUFX2_insert233 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236_),
    .Y(_1236__bF$buf3)
);

BUFX2 BUFX2_insert232 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236_),
    .Y(_1236__bF$buf4)
);

BUFX2 BUFX2_insert231 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5927_),
    .Y(_5927__bF$buf0)
);

BUFX2 BUFX2_insert230 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5927_),
    .Y(_5927__bF$buf1)
);

BUFX2 BUFX2_insert229 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5927_),
    .Y(_5927__bF$buf2)
);

BUFX2 BUFX2_insert228 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5927_),
    .Y(_5927__bF$buf3)
);

BUFX2 BUFX2_insert227 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5927_),
    .Y(_5927__bF$buf4)
);

BUFX2 BUFX2_insert226 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3267_),
    .Y(_3267__bF$buf0)
);

BUFX2 BUFX2_insert225 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3267_),
    .Y(_3267__bF$buf1)
);

BUFX2 BUFX2_insert224 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3267_),
    .Y(_3267__bF$buf2)
);

BUFX2 BUFX2_insert223 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3267_),
    .Y(_3267__bF$buf3)
);

BUFX2 BUFX2_insert222 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3267_),
    .Y(_3267__bF$buf4)
);

BUFX2 BUFX2_insert221 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3267_),
    .Y(_3267__bF$buf5)
);

BUFX2 BUFX2_insert220 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3267_),
    .Y(_3267__bF$buf6)
);

BUFX2 BUFX2_insert219 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .Y(_5510__bF$buf0)
);

BUFX2 BUFX2_insert218 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .Y(_5510__bF$buf1)
);

BUFX2 BUFX2_insert217 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .Y(_5510__bF$buf2)
);

BUFX2 BUFX2_insert216 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .Y(_5510__bF$buf3)
);

BUFX2 BUFX2_insert215 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .Y(_5510__bF$buf4)
);

BUFX2 BUFX2_insert214 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .Y(_5510__bF$buf5)
);

BUFX2 BUFX2_insert213 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .Y(_5510__bF$buf6)
);

BUFX2 BUFX2_insert212 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .Y(_5510__bF$buf7)
);

BUFX2 BUFX2_insert211 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .Y(_5510__bF$buf8)
);

BUFX2 BUFX2_insert210 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .Y(_5510__bF$buf9)
);

BUFX2 BUFX2_insert209 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .Y(_5510__bF$buf10)
);

BUFX2 BUFX2_insert208 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .Y(_5510__bF$buf11)
);

BUFX2 BUFX2_insert207 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .Y(_5510__bF$buf12)
);

BUFX2 BUFX2_insert206 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .Y(_5510__bF$buf13)
);

BUFX2 BUFX2_insert205 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .Y(_5510__bF$buf14)
);

BUFX2 BUFX2_insert204 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .Y(_5510__bF$buf15)
);

BUFX2 BUFX2_insert203 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [18]),
    .Y(\datapath.idinstr_18_bF$buf0 )
);

BUFX2 BUFX2_insert202 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [18]),
    .Y(\datapath.idinstr_18_bF$buf1 )
);

BUFX2 BUFX2_insert201 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [18]),
    .Y(\datapath.idinstr_18_bF$buf2 )
);

BUFX2 BUFX2_insert200 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [18]),
    .Y(\datapath.idinstr_18_bF$buf3 )
);

BUFX2 BUFX2_insert199 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [18]),
    .Y(\datapath.idinstr_18_bF$buf4 )
);

BUFX2 BUFX2_insert198 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [18]),
    .Y(\datapath.idinstr_18_bF$buf5 )
);

BUFX2 BUFX2_insert197 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [18]),
    .Y(\datapath.idinstr_18_bF$buf6 )
);

BUFX2 BUFX2_insert196 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [18]),
    .Y(\datapath.idinstr_18_bF$buf7 )
);

BUFX2 BUFX2_insert195 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3690_),
    .Y(_3690__bF$buf0)
);

BUFX2 BUFX2_insert194 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3690_),
    .Y(_3690__bF$buf1)
);

BUFX2 BUFX2_insert193 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3690_),
    .Y(_3690__bF$buf2)
);

BUFX2 BUFX2_insert192 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3690_),
    .Y(_3690__bF$buf3)
);

BUFX2 BUFX2_insert191 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3690_),
    .Y(_3690__bF$buf4)
);

BUFX2 BUFX2_insert190 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_21_bF$buf0 )
);

BUFX2 BUFX2_insert189 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_21_bF$buf1 )
);

BUFX2 BUFX2_insert188 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_21_bF$buf2 )
);

BUFX2 BUFX2_insert187 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_21_bF$buf3 )
);

BUFX2 BUFX2_insert186 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_21_bF$buf4 )
);

BUFX2 BUFX2_insert185 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_21_bF$buf5 )
);

BUFX2 BUFX2_insert184 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_21_bF$buf6 )
);

BUFX2 BUFX2_insert183 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_21_bF$buf7 )
);

BUFX2 BUFX2_insert182 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_21_bF$buf8 )
);

BUFX2 BUFX2_insert181 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_21_bF$buf9 )
);

BUFX2 BUFX2_insert180 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_21_bF$buf10 )
);

BUFX2 BUFX2_insert179 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_21_bF$buf11 )
);

BUFX2 BUFX2_insert178 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_21_bF$buf12 )
);

BUFX2 BUFX2_insert177 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_21_bF$buf13 )
);

BUFX2 BUFX2_insert176 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_21_bF$buf14 )
);

BUFX2 BUFX2_insert175 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_21_bF$buf15 )
);

BUFX2 BUFX2_insert174 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_21_bF$buf16 )
);

BUFX2 BUFX2_insert173 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_21_bF$buf17 )
);

BUFX2 BUFX2_insert172 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_21_bF$buf18 )
);

BUFX2 BUFX2_insert171 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_21_bF$buf19 )
);

BUFX2 BUFX2_insert170 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_21_bF$buf20 )
);

BUFX2 BUFX2_insert169 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_21_bF$buf21 )
);

BUFX2 BUFX2_insert168 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_21_bF$buf22 )
);

BUFX2 BUFX2_insert167 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_21_bF$buf23 )
);

BUFX2 BUFX2_insert166 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_21_bF$buf24 )
);

BUFX2 BUFX2_insert165 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_21_bF$buf25 )
);

BUFX2 BUFX2_insert164 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_21_bF$buf26 )
);

BUFX2 BUFX2_insert163 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_21_bF$buf27 )
);

BUFX2 BUFX2_insert162 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_21_bF$buf28 )
);

BUFX2 BUFX2_insert161 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_21_bF$buf29 )
);

BUFX2 BUFX2_insert160 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_21_bF$buf30 )
);

BUFX2 BUFX2_insert159 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_21_bF$buf31 )
);

BUFX2 BUFX2_insert158 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_21_bF$buf32 )
);

BUFX2 BUFX2_insert157 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_21_bF$buf33 )
);

BUFX2 BUFX2_insert156 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_21_bF$buf34 )
);

BUFX2 BUFX2_insert155 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_21_bF$buf35 )
);

BUFX2 BUFX2_insert154 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_21_bF$buf36 )
);

BUFX2 BUFX2_insert153 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_21_bF$buf37 )
);

BUFX2 BUFX2_insert152 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_21_bF$buf38 )
);

BUFX2 BUFX2_insert151 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf2 ),
    .Y(\datapath.idinstr_21_bF$buf39 )
);

BUFX2 BUFX2_insert150 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf1 ),
    .Y(\datapath.idinstr_21_bF$buf40 )
);

BUFX2 BUFX2_insert149 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf0 ),
    .Y(\datapath.idinstr_21_bF$buf41 )
);

BUFX2 BUFX2_insert148 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf5 ),
    .Y(\datapath.idinstr_21_bF$buf42 )
);

BUFX2 BUFX2_insert147 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf4 ),
    .Y(\datapath.idinstr_21_bF$buf43 )
);

BUFX2 BUFX2_insert146 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_hier0_bF$buf3 ),
    .Y(\datapath.idinstr_21_bF$buf44 )
);

BUFX2 BUFX2_insert145 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492_),
    .Y(_5492__bF$buf0)
);

BUFX2 BUFX2_insert144 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492_),
    .Y(_5492__bF$buf1)
);

BUFX2 BUFX2_insert143 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492_),
    .Y(_5492__bF$buf2)
);

BUFX2 BUFX2_insert142 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492_),
    .Y(_5492__bF$buf3)
);

BUFX2 BUFX2_insert141 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492_),
    .Y(_5492__bF$buf4)
);

BUFX2 BUFX2_insert140 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9343_),
    .Y(_9343__bF$buf0)
);

BUFX2 BUFX2_insert139 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9343_),
    .Y(_9343__bF$buf1)
);

BUFX2 BUFX2_insert138 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9343_),
    .Y(_9343__bF$buf2)
);

BUFX2 BUFX2_insert137 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9343_),
    .Y(_9343__bF$buf3)
);

BUFX2 BUFX2_insert136 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9343_),
    .Y(_9343__bF$buf4)
);

BUFX2 BUFX2_insert135 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9343_),
    .Y(_9343__bF$buf5)
);

BUFX2 BUFX2_insert134 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9343_),
    .Y(_9343__bF$buf6)
);

BUFX2 BUFX2_insert133 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9343_),
    .Y(_9343__bF$buf7)
);

BUFX2 BUFX2_insert132 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454_),
    .Y(_5454__bF$buf0)
);

BUFX2 BUFX2_insert131 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454_),
    .Y(_5454__bF$buf1)
);

BUFX2 BUFX2_insert130 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454_),
    .Y(_5454__bF$buf2)
);

BUFX2 BUFX2_insert129 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454_),
    .Y(_5454__bF$buf3)
);

BUFX2 BUFX2_insert128 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454_),
    .Y(_5454__bF$buf4)
);

BUFX2 BUFX2_insert127 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6145_),
    .Y(_6145__bF$buf0)
);

BUFX2 BUFX2_insert126 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6145_),
    .Y(_6145__bF$buf1)
);

BUFX2 BUFX2_insert125 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6145_),
    .Y(_6145__bF$buf2)
);

BUFX2 BUFX2_insert124 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6145_),
    .Y(_6145__bF$buf3)
);

BUFX2 BUFX2_insert123 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6145_),
    .Y(_6145__bF$buf4)
);

BUFX2 BUFX2_insert122 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6145_),
    .Y(_6145__bF$buf5)
);

BUFX2 BUFX2_insert121 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6145_),
    .Y(_6145__bF$buf6)
);

BUFX2 BUFX2_insert120 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6145_),
    .Y(_6145__bF$buf7)
);

BUFX2 BUFX2_insert119 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211_),
    .Y(_9211__bF$buf0)
);

BUFX2 BUFX2_insert118 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211_),
    .Y(_9211__bF$buf1)
);

BUFX2 BUFX2_insert117 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211_),
    .Y(_9211__bF$buf2)
);

BUFX2 BUFX2_insert116 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211_),
    .Y(_9211__bF$buf3)
);

BUFX2 BUFX2_insert115 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211_),
    .Y(_9211__bF$buf4)
);

BUFX2 BUFX2_insert114 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211_),
    .Y(_9211__bF$buf5)
);

BUFX2 BUFX2_insert113 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211_),
    .Y(_9211__bF$buf6)
);

BUFX2 BUFX2_insert112 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211_),
    .Y(_9211__bF$buf7)
);

BUFX2 BUFX2_insert111 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211_),
    .Y(_9211__bF$buf8)
);

BUFX2 BUFX2_insert110 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1242_),
    .Y(_1242__bF$buf0)
);

BUFX2 BUFX2_insert109 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1242_),
    .Y(_1242__bF$buf1)
);

BUFX2 BUFX2_insert108 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1242_),
    .Y(_1242__bF$buf2)
);

BUFX2 BUFX2_insert107 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1242_),
    .Y(_1242__bF$buf3)
);

BUFX2 BUFX2_insert106 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1242_),
    .Y(_1242__bF$buf4)
);

BUFX2 BUFX2_insert105 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6107_),
    .Y(_6107__bF$buf0)
);

BUFX2 BUFX2_insert104 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6107_),
    .Y(_6107__bF$buf1)
);

BUFX2 BUFX2_insert103 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6107_),
    .Y(_6107__bF$buf2)
);

BUFX2 BUFX2_insert102 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6107_),
    .Y(_6107__bF$buf3)
);

BUFX2 BUFX2_insert101 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6107_),
    .Y(_6107__bF$buf4)
);

BUFX2 BUFX2_insert100 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193_),
    .Y(_4193__bF$buf0)
);

BUFX2 BUFX2_insert99 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193_),
    .Y(_4193__bF$buf1)
);

BUFX2 BUFX2_insert98 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193_),
    .Y(_4193__bF$buf2)
);

BUFX2 BUFX2_insert97 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193_),
    .Y(_4193__bF$buf3)
);

BUFX2 BUFX2_insert96 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193_),
    .Y(_4193__bF$buf4)
);

BUFX2 BUFX2_insert95 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [24]),
    .Y(\datapath.idinstr_24_bF$buf0 )
);

BUFX2 BUFX2_insert94 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [24]),
    .Y(\datapath.idinstr_24_bF$buf1 )
);

BUFX2 BUFX2_insert93 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [24]),
    .Y(\datapath.idinstr_24_bF$buf2 )
);

BUFX2 BUFX2_insert92 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [24]),
    .Y(\datapath.idinstr_24_bF$buf3 )
);

BUFX2 BUFX2_insert91 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [24]),
    .Y(\datapath.idinstr_24_bF$buf4 )
);

BUFX2 BUFX2_insert90 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [24]),
    .Y(\datapath.idinstr_24_bF$buf5 )
);

BUFX2 BUFX2_insert89 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5648_),
    .Y(_5648__bF$buf0)
);

BUFX2 BUFX2_insert88 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5648_),
    .Y(_5648__bF$buf1)
);

BUFX2 BUFX2_insert87 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5648_),
    .Y(_5648__bF$buf2)
);

BUFX2 BUFX2_insert86 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5648_),
    .Y(_5648__bF$buf3)
);

BUFX2 BUFX2_insert85 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5648_),
    .Y(_5648__bF$buf4)
);

BUFX2 BUFX2_insert84 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460_),
    .Y(_5460__bF$buf0)
);

BUFX2 BUFX2_insert83 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460_),
    .Y(_5460__bF$buf1)
);

BUFX2 BUFX2_insert82 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460_),
    .Y(_5460__bF$buf2)
);

BUFX2 BUFX2_insert81 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460_),
    .Y(_5460__bF$buf3)
);

BUFX2 BUFX2_insert80 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460_),
    .Y(_5460__bF$buf4)
);

BUFX2 BUFX2_insert79 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4196_),
    .Y(_4196__bF$buf0)
);

BUFX2 BUFX2_insert78 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4196_),
    .Y(_4196__bF$buf1)
);

BUFX2 BUFX2_insert77 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4196_),
    .Y(_4196__bF$buf2)
);

BUFX2 BUFX2_insert76 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4196_),
    .Y(_4196__bF$buf3)
);

BUFX2 BUFX2_insert75 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4196_),
    .Y(_4196__bF$buf4)
);

BUFX2 BUFX2_insert74 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498_),
    .Y(_5498__bF$buf0)
);

BUFX2 BUFX2_insert73 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498_),
    .Y(_5498__bF$buf1)
);

BUFX2 BUFX2_insert72 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498_),
    .Y(_5498__bF$buf2)
);

BUFX2 BUFX2_insert71 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498_),
    .Y(_5498__bF$buf3)
);

BUFX2 BUFX2_insert70 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498_),
    .Y(_5498__bF$buf4)
);

BUFX2 BUFX2_insert69 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2703_),
    .Y(_2703__bF$buf0)
);

BUFX2 BUFX2_insert68 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2703_),
    .Y(_2703__bF$buf1)
);

BUFX2 BUFX2_insert67 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2703_),
    .Y(_2703__bF$buf2)
);

BUFX2 BUFX2_insert66 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2703_),
    .Y(_2703__bF$buf3)
);

BUFX2 BUFX2_insert65 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3796_),
    .Y(_3796__bF$buf0)
);

BUFX2 BUFX2_insert64 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3796_),
    .Y(_3796__bF$buf1)
);

BUFX2 BUFX2_insert63 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3796_),
    .Y(_3796__bF$buf2)
);

BUFX2 BUFX2_insert62 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3796_),
    .Y(_3796__bF$buf3)
);

BUFX2 BUFX2_insert61 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3796_),
    .Y(_3796__bF$buf4)
);

BUFX2 BUFX2_insert60 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_964_),
    .Y(_964__bF$buf0)
);

BUFX2 BUFX2_insert59 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_964_),
    .Y(_964__bF$buf1)
);

BUFX2 BUFX2_insert58 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_964_),
    .Y(_964__bF$buf2)
);

BUFX2 BUFX2_insert57 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_964_),
    .Y(_964__bF$buf3)
);

BUFX2 BUFX2_insert56 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_964_),
    .Y(_964__bF$buf4)
);

BUFX2 BUFX2_insert55 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2706_),
    .Y(_2706__bF$buf0)
);

BUFX2 BUFX2_insert54 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2706_),
    .Y(_2706__bF$buf1)
);

BUFX2 BUFX2_insert53 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2706_),
    .Y(_2706__bF$buf2)
);

BUFX2 BUFX2_insert52 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2706_),
    .Y(_2706__bF$buf3)
);

BUFX2 BUFX2_insert51 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [2]),
    .Y(\datapath.alu.b_2_bF$buf0 )
);

BUFX2 BUFX2_insert50 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [2]),
    .Y(\datapath.alu.b_2_bF$buf1 )
);

BUFX2 BUFX2_insert49 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [2]),
    .Y(\datapath.alu.b_2_bF$buf2 )
);

BUFX2 BUFX2_insert48 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [2]),
    .Y(\datapath.alu.b_2_bF$buf3 )
);

BUFX2 BUFX2_insert47 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [2]),
    .Y(\datapath.alu.b_2_bF$buf4 )
);

BUFX2 BUFX2_insert46 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [2]),
    .Y(\datapath.alu.b_2_bF$buf5 )
);

BUFX2 BUFX2_insert45 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [2]),
    .Y(\datapath.alu.b_2_bF$buf6 )
);

BUFX2 BUFX2_insert44 (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [2]),
    .Y(\datapath.alu.b_2_bF$buf7 )
);

BUFX2 BUFX2_insert43 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .Y(_297__bF$buf0)
);

BUFX2 BUFX2_insert42 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .Y(_297__bF$buf1)
);

BUFX2 BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .Y(_297__bF$buf2)
);

BUFX2 BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .Y(_297__bF$buf3)
);

BUFX2 BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .Y(_297__bF$buf4)
);

BUFX2 BUFX2_insert38 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .Y(_297__bF$buf5)
);

BUFX2 BUFX2_insert37 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .Y(_297__bF$buf6)
);

BUFX2 BUFX2_insert36 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .Y(_297__bF$buf7)
);

BUFX2 BUFX2_insert35 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .Y(_297__bF$buf8)
);

BUFX2 BUFX2_insert34 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7612_),
    .Y(_7612__bF$buf0)
);

BUFX2 BUFX2_insert33 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7612_),
    .Y(_7612__bF$buf1)
);

BUFX2 BUFX2_insert32 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7612_),
    .Y(_7612__bF$buf2)
);

BUFX2 BUFX2_insert31 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7612_),
    .Y(_7612__bF$buf3)
);

BUFX2 BUFX2_insert30 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7612_),
    .Y(_7612__bF$buf4)
);

BUFX2 BUFX2_insert29 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7612_),
    .Y(_7612__bF$buf5)
);

BUFX2 BUFX2_insert28 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7612_),
    .Y(_7612__bF$buf6)
);

BUFX2 BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7612_),
    .Y(_7612__bF$buf7)
);

BUFX2 BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466_),
    .Y(_5466__bF$buf0)
);

BUFX2 BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466_),
    .Y(_5466__bF$buf1)
);

BUFX2 BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466_),
    .Y(_5466__bF$buf2)
);

BUFX2 BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466_),
    .Y(_5466__bF$buf3)
);

BUFX2 BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466_),
    .Y(_5466__bF$buf4)
);

BUFX2 BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497_),
    .Y(_2497__bF$buf0)
);

BUFX2 BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497_),
    .Y(_2497__bF$buf1)
);

BUFX2 BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497_),
    .Y(_2497__bF$buf2)
);

BUFX2 BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497_),
    .Y(_2497__bF$buf3)
);

BUFX2 BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497_),
    .Y(_2497__bF$buf4)
);

BUFX2 BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497_),
    .Y(_2497__bF$buf5)
);

BUFX2 BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497_),
    .Y(_2497__bF$buf6)
);

BUFX2 BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2688_),
    .Y(_2688__bF$buf0)
);

BUFX2 BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2688_),
    .Y(_2688__bF$buf1)
);

BUFX2 BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2688_),
    .Y(_2688__bF$buf2)
);

BUFX2 BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2688_),
    .Y(_2688__bF$buf3)
);

BUFX2 BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_970_),
    .Y(_970__bF$buf0)
);

BUFX2 BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_970_),
    .Y(_970__bF$buf1)
);

BUFX2 BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_970_),
    .Y(_970__bF$buf2)
);

BUFX2 BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_970_),
    .Y(_970__bF$buf3)
);

BUFX2 BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_970_),
    .Y(_970__bF$buf4)
);

BUFX2 BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250_),
    .Y(_3250__bF$buf0)
);

BUFX2 BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250_),
    .Y(_3250__bF$buf1)
);

BUFX2 BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250_),
    .Y(_3250__bF$buf2)
);

BUFX2 BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250_),
    .Y(_3250__bF$buf3)
);

BUFX2 BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250_),
    .Y(_3250__bF$buf4)
);

BUFX2 BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250_),
    .Y(_3250__bF$buf5)
);

INVX1 _10000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [6]),
    .Y(_370_)
);

NAND2X1 _10001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [6]),
    .B(_297__bF$buf8),
    .Y(_371_)
);

OAI21X1 _10002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf7),
    .B(_370_),
    .C(_371_),
    .Y(\datapath._05_ [6])
);

INVX1 _10003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [7]),
    .Y(_372_)
);

NAND2X1 _10004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [7]),
    .B(_297__bF$buf6),
    .Y(_373_)
);

OAI21X1 _10005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf5),
    .B(_372_),
    .C(_373_),
    .Y(\datapath._05_ [7])
);

INVX1 _10006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [8]),
    .Y(_374_)
);

NAND2X1 _10007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [8]),
    .B(_297__bF$buf4),
    .Y(_375_)
);

OAI21X1 _10008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf3),
    .B(_374_),
    .C(_375_),
    .Y(\datapath._05_ [8])
);

INVX1 _10009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [9]),
    .Y(_376_)
);

NAND2X1 _10010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [9]),
    .B(_297__bF$buf2),
    .Y(_377_)
);

OAI21X1 _10011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf1),
    .B(_376_),
    .C(_377_),
    .Y(\datapath._05_ [9])
);

INVX1 _10012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [10]),
    .Y(_378_)
);

NAND2X1 _10013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [10]),
    .B(_297__bF$buf0),
    .Y(_379_)
);

OAI21X1 _10014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf8),
    .B(_378_),
    .C(_379_),
    .Y(\datapath._05_ [10])
);

INVX1 _10015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [11]),
    .Y(_380_)
);

NAND2X1 _10016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [11]),
    .B(_297__bF$buf7),
    .Y(_381_)
);

OAI21X1 _10017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf6),
    .B(_380_),
    .C(_381_),
    .Y(\datapath._05_ [11])
);

INVX1 _10018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [12]),
    .Y(_382_)
);

NAND2X1 _10019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [12]),
    .B(_297__bF$buf5),
    .Y(_383_)
);

OAI21X1 _10020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf4),
    .B(_382_),
    .C(_383_),
    .Y(\datapath._05_ [12])
);

INVX1 _10021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [13]),
    .Y(_384_)
);

NAND2X1 _10022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [13]),
    .B(_297__bF$buf3),
    .Y(_385_)
);

OAI21X1 _10023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf2),
    .B(_384_),
    .C(_385_),
    .Y(\datapath._05_ [13])
);

INVX1 _10024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [14]),
    .Y(_386_)
);

NAND2X1 _10025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [14]),
    .B(_297__bF$buf1),
    .Y(_387_)
);

OAI21X1 _10026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf0),
    .B(_386_),
    .C(_387_),
    .Y(\datapath._05_ [14])
);

INVX1 _10027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [15]),
    .Y(_388_)
);

NAND2X1 _10028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [15]),
    .B(_297__bF$buf8),
    .Y(_389_)
);

OAI21X1 _10029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf7),
    .B(_388_),
    .C(_389_),
    .Y(\datapath._05_ [15])
);

INVX1 _10030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [16]),
    .Y(_390_)
);

NAND2X1 _10031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [16]),
    .B(_297__bF$buf6),
    .Y(_391_)
);

OAI21X1 _10032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf5),
    .B(_390_),
    .C(_391_),
    .Y(\datapath._05_ [16])
);

INVX1 _10033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [17]),
    .Y(_392_)
);

NAND2X1 _10034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [17]),
    .B(_297__bF$buf4),
    .Y(_393_)
);

OAI21X1 _10035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf3),
    .B(_392_),
    .C(_393_),
    .Y(\datapath._05_ [17])
);

INVX1 _10036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [18]),
    .Y(_394_)
);

NAND2X1 _10037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [18]),
    .B(_297__bF$buf2),
    .Y(_395_)
);

OAI21X1 _10038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf1),
    .B(_394_),
    .C(_395_),
    .Y(\datapath._05_ [18])
);

INVX1 _10039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [19]),
    .Y(_396_)
);

NAND2X1 _10040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [19]),
    .B(_297__bF$buf0),
    .Y(_397_)
);

OAI21X1 _10041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf8),
    .B(_396_),
    .C(_397_),
    .Y(\datapath._05_ [19])
);

INVX1 _10042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [20]),
    .Y(_398_)
);

NAND2X1 _10043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [20]),
    .B(_297__bF$buf7),
    .Y(_399_)
);

OAI21X1 _10044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf6),
    .B(_398_),
    .C(_399_),
    .Y(\datapath._05_ [20])
);

INVX1 _10045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [21]),
    .Y(_400_)
);

NAND2X1 _10046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [21]),
    .B(_297__bF$buf5),
    .Y(_401_)
);

OAI21X1 _10047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf4),
    .B(_400_),
    .C(_401_),
    .Y(\datapath._05_ [21])
);

INVX1 _10048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [22]),
    .Y(_402_)
);

NAND2X1 _10049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [22]),
    .B(_297__bF$buf3),
    .Y(_403_)
);

OAI21X1 _10050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf2),
    .B(_402_),
    .C(_403_),
    .Y(\datapath._05_ [22])
);

INVX1 _10051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [23]),
    .Y(_404_)
);

NAND2X1 _10052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [23]),
    .B(_297__bF$buf1),
    .Y(_405_)
);

OAI21X1 _10053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf0),
    .B(_404_),
    .C(_405_),
    .Y(\datapath._05_ [23])
);

INVX1 _10054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [24]),
    .Y(_406_)
);

NAND2X1 _10055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [24]),
    .B(_297__bF$buf8),
    .Y(_407_)
);

OAI21X1 _10056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf7),
    .B(_406_),
    .C(_407_),
    .Y(\datapath._05_ [24])
);

INVX1 _10057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [25]),
    .Y(_408_)
);

NAND2X1 _10058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [25]),
    .B(_297__bF$buf6),
    .Y(_409_)
);

OAI21X1 _10059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf5),
    .B(_408_),
    .C(_409_),
    .Y(\datapath._05_ [25])
);

INVX1 _10060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [26]),
    .Y(_410_)
);

NAND2X1 _10061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [26]),
    .B(_297__bF$buf4),
    .Y(_411_)
);

OAI21X1 _10062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf3),
    .B(_410_),
    .C(_411_),
    .Y(\datapath._05_ [26])
);

INVX1 _10063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [27]),
    .Y(_412_)
);

NAND2X1 _10064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [27]),
    .B(_297__bF$buf2),
    .Y(_413_)
);

OAI21X1 _10065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf1),
    .B(_412_),
    .C(_413_),
    .Y(\datapath._05_ [27])
);

INVX1 _10066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [28]),
    .Y(_414_)
);

NAND2X1 _10067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [28]),
    .B(_297__bF$buf0),
    .Y(_415_)
);

OAI21X1 _10068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf8),
    .B(_414_),
    .C(_415_),
    .Y(\datapath._05_ [28])
);

INVX1 _10069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [29]),
    .Y(_416_)
);

NAND2X1 _10070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [29]),
    .B(_297__bF$buf7),
    .Y(_417_)
);

OAI21X1 _10071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf6),
    .B(_416_),
    .C(_417_),
    .Y(\datapath._05_ [29])
);

INVX1 _10072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [30]),
    .Y(_418_)
);

NAND2X1 _10073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [30]),
    .B(_297__bF$buf5),
    .Y(_419_)
);

OAI21X1 _10074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf4),
    .B(_418_),
    .C(_419_),
    .Y(\datapath._05_ [30])
);

INVX1 _10075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [31]),
    .Y(_420_)
);

NAND2X1 _10076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [31]),
    .B(_297__bF$buf3),
    .Y(_421_)
);

OAI21X1 _10077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf2),
    .B(_420_),
    .C(_421_),
    .Y(\datapath._05_ [31])
);

INVX1 _10078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [0]),
    .Y(_422_)
);

NAND2X1 _10079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf9 ),
    .B(\datapath.idpc_4 [0]),
    .Y(_423_)
);

OAI21X1 _10080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_422_),
    .B(\bypassandflushunit.stall_bF$buf8 ),
    .C(_423_),
    .Y(\datapath._06_ [0])
);

INVX1 _10081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [1]),
    .Y(_424_)
);

NAND2X1 _10082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf7 ),
    .B(\datapath.idpc_4 [1]),
    .Y(_425_)
);

OAI21X1 _10083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_424_),
    .B(\bypassandflushunit.stall_bF$buf6 ),
    .C(_425_),
    .Y(\datapath._06_ [1])
);

INVX1 _10084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [2]),
    .Y(_426_)
);

NAND2X1 _10085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf5 ),
    .B(\datapath.idpc_4 [2]),
    .Y(_427_)
);

OAI21X1 _10086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_426_),
    .B(\bypassandflushunit.stall_bF$buf4 ),
    .C(_427_),
    .Y(\datapath._06_ [2])
);

INVX1 _10087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [3]),
    .Y(_428_)
);

NAND2X1 _10088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf3 ),
    .B(\datapath.idpc_4 [3]),
    .Y(_429_)
);

OAI21X1 _10089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_428_),
    .B(\bypassandflushunit.stall_bF$buf2 ),
    .C(_429_),
    .Y(\datapath._06_ [3])
);

INVX1 _10090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [4]),
    .Y(_430_)
);

NAND2X1 _10091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf1 ),
    .B(\datapath.idpc_4 [4]),
    .Y(_431_)
);

OAI21X1 _10092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_430_),
    .B(\bypassandflushunit.stall_bF$buf0 ),
    .C(_431_),
    .Y(\datapath._06_ [4])
);

INVX1 _10093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [5]),
    .Y(_432_)
);

NAND2X1 _10094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf9 ),
    .B(\datapath.idpc_4 [5]),
    .Y(_433_)
);

OAI21X1 _10095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_432_),
    .B(\bypassandflushunit.stall_bF$buf8 ),
    .C(_433_),
    .Y(\datapath._06_ [5])
);

INVX1 _10096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [6]),
    .Y(_434_)
);

NAND2X1 _10097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf7 ),
    .B(\datapath.idpc_4 [6]),
    .Y(_435_)
);

OAI21X1 _10098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_434_),
    .B(\bypassandflushunit.stall_bF$buf6 ),
    .C(_435_),
    .Y(\datapath._06_ [6])
);

INVX1 _10099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [7]),
    .Y(_436_)
);

NAND2X1 _10100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf5 ),
    .B(\datapath.idpc_4 [7]),
    .Y(_437_)
);

OAI21X1 _10101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_436_),
    .B(\bypassandflushunit.stall_bF$buf4 ),
    .C(_437_),
    .Y(\datapath._06_ [7])
);

INVX1 _10102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [8]),
    .Y(_438_)
);

NAND2X1 _10103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf3 ),
    .B(\datapath.idpc_4 [8]),
    .Y(_439_)
);

OAI21X1 _10104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_438_),
    .B(\bypassandflushunit.stall_bF$buf2 ),
    .C(_439_),
    .Y(\datapath._06_ [8])
);

INVX1 _10105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [9]),
    .Y(_440_)
);

NAND2X1 _10106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf1 ),
    .B(\datapath.idpc_4 [9]),
    .Y(_441_)
);

OAI21X1 _10107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_440_),
    .B(\bypassandflushunit.stall_bF$buf0 ),
    .C(_441_),
    .Y(\datapath._06_ [9])
);

INVX1 _10108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [10]),
    .Y(_442_)
);

NAND2X1 _10109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf9 ),
    .B(\datapath.idpc_4 [10]),
    .Y(_443_)
);

OAI21X1 _10110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_442_),
    .B(\bypassandflushunit.stall_bF$buf8 ),
    .C(_443_),
    .Y(\datapath._06_ [10])
);

INVX1 _10111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [11]),
    .Y(_444_)
);

NAND2X1 _10112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf7 ),
    .B(\datapath.idpc_4 [11]),
    .Y(_445_)
);

OAI21X1 _10113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_444_),
    .B(\bypassandflushunit.stall_bF$buf6 ),
    .C(_445_),
    .Y(\datapath._06_ [11])
);

INVX1 _10114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [12]),
    .Y(_446_)
);

NAND2X1 _10115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf5 ),
    .B(\datapath.idpc_4 [12]),
    .Y(_447_)
);

OAI21X1 _10116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_446_),
    .B(\bypassandflushunit.stall_bF$buf4 ),
    .C(_447_),
    .Y(\datapath._06_ [12])
);

INVX1 _10117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [13]),
    .Y(_448_)
);

NAND2X1 _10118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf3 ),
    .B(\datapath.idpc_4 [13]),
    .Y(_449_)
);

OAI21X1 _10119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_448_),
    .B(\bypassandflushunit.stall_bF$buf2 ),
    .C(_449_),
    .Y(\datapath._06_ [13])
);

INVX1 _10120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [14]),
    .Y(_450_)
);

NAND2X1 _10121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf1 ),
    .B(\datapath.idpc_4 [14]),
    .Y(_451_)
);

OAI21X1 _10122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_450_),
    .B(\bypassandflushunit.stall_bF$buf0 ),
    .C(_451_),
    .Y(\datapath._06_ [14])
);

INVX1 _10123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [15]),
    .Y(_452_)
);

NAND2X1 _10124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf9 ),
    .B(\datapath.idpc_4 [15]),
    .Y(_453_)
);

OAI21X1 _10125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_452_),
    .B(\bypassandflushunit.stall_bF$buf8 ),
    .C(_453_),
    .Y(\datapath._06_ [15])
);

INVX1 _10126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [16]),
    .Y(_454_)
);

NAND2X1 _10127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf7 ),
    .B(\datapath.idpc_4 [16]),
    .Y(_455_)
);

OAI21X1 _10128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_454_),
    .B(\bypassandflushunit.stall_bF$buf6 ),
    .C(_455_),
    .Y(\datapath._06_ [16])
);

INVX1 _10129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [17]),
    .Y(_456_)
);

NAND2X1 _10130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf5 ),
    .B(\datapath.idpc_4 [17]),
    .Y(_457_)
);

OAI21X1 _10131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_456_),
    .B(\bypassandflushunit.stall_bF$buf4 ),
    .C(_457_),
    .Y(\datapath._06_ [17])
);

INVX1 _10132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [18]),
    .Y(_458_)
);

NAND2X1 _10133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf3 ),
    .B(\datapath.idpc_4 [18]),
    .Y(_459_)
);

OAI21X1 _10134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_458_),
    .B(\bypassandflushunit.stall_bF$buf2 ),
    .C(_459_),
    .Y(\datapath._06_ [18])
);

INVX1 _10135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [19]),
    .Y(_460_)
);

NAND2X1 _10136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf1 ),
    .B(\datapath.idpc_4 [19]),
    .Y(_461_)
);

OAI21X1 _10137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_460_),
    .B(\bypassandflushunit.stall_bF$buf0 ),
    .C(_461_),
    .Y(\datapath._06_ [19])
);

INVX1 _10138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [20]),
    .Y(_462_)
);

NAND2X1 _10139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf9 ),
    .B(\datapath.idpc_4 [20]),
    .Y(_463_)
);

OAI21X1 _10140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_462_),
    .B(\bypassandflushunit.stall_bF$buf8 ),
    .C(_463_),
    .Y(\datapath._06_ [20])
);

INVX1 _10141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [21]),
    .Y(_464_)
);

NAND2X1 _10142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf7 ),
    .B(\datapath.idpc_4 [21]),
    .Y(_465_)
);

OAI21X1 _10143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_464_),
    .B(\bypassandflushunit.stall_bF$buf6 ),
    .C(_465_),
    .Y(\datapath._06_ [21])
);

INVX1 _10144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [22]),
    .Y(_466_)
);

NAND2X1 _10145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf5 ),
    .B(\datapath.idpc_4 [22]),
    .Y(_467_)
);

OAI21X1 _10146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_466_),
    .B(\bypassandflushunit.stall_bF$buf4 ),
    .C(_467_),
    .Y(\datapath._06_ [22])
);

INVX1 _10147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [23]),
    .Y(_468_)
);

NAND2X1 _10148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf3 ),
    .B(\datapath.idpc_4 [23]),
    .Y(_469_)
);

OAI21X1 _10149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_468_),
    .B(\bypassandflushunit.stall_bF$buf2 ),
    .C(_469_),
    .Y(\datapath._06_ [23])
);

INVX1 _10150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [24]),
    .Y(_470_)
);

NAND2X1 _10151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf1 ),
    .B(\datapath.idpc_4 [24]),
    .Y(_471_)
);

OAI21X1 _10152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470_),
    .B(\bypassandflushunit.stall_bF$buf0 ),
    .C(_471_),
    .Y(\datapath._06_ [24])
);

INVX1 _10153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [25]),
    .Y(_472_)
);

NAND2X1 _10154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf9 ),
    .B(\datapath.idpc_4 [25]),
    .Y(_473_)
);

OAI21X1 _10155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_472_),
    .B(\bypassandflushunit.stall_bF$buf8 ),
    .C(_473_),
    .Y(\datapath._06_ [25])
);

INVX1 _10156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [26]),
    .Y(_474_)
);

NAND2X1 _10157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf7 ),
    .B(\datapath.idpc_4 [26]),
    .Y(_475_)
);

OAI21X1 _10158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_474_),
    .B(\bypassandflushunit.stall_bF$buf6 ),
    .C(_475_),
    .Y(\datapath._06_ [26])
);

INVX1 _10159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [27]),
    .Y(_476_)
);

NAND2X1 _10160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf5 ),
    .B(\datapath.idpc_4 [27]),
    .Y(_477_)
);

OAI21X1 _10161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_476_),
    .B(\bypassandflushunit.stall_bF$buf4 ),
    .C(_477_),
    .Y(\datapath._06_ [27])
);

INVX1 _10162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [28]),
    .Y(_478_)
);

NAND2X1 _10163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf3 ),
    .B(\datapath.idpc_4 [28]),
    .Y(_479_)
);

OAI21X1 _10164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_478_),
    .B(\bypassandflushunit.stall_bF$buf2 ),
    .C(_479_),
    .Y(\datapath._06_ [28])
);

INVX1 _10165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [29]),
    .Y(_480_)
);

NAND2X1 _10166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf1 ),
    .B(\datapath.idpc_4 [29]),
    .Y(_481_)
);

OAI21X1 _10167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_480_),
    .B(\bypassandflushunit.stall_bF$buf0 ),
    .C(_481_),
    .Y(\datapath._06_ [29])
);

INVX1 _10168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [30]),
    .Y(_482_)
);

NAND2X1 _10169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf9 ),
    .B(\datapath.idpc_4 [30]),
    .Y(_483_)
);

OAI21X1 _10170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_482_),
    .B(\bypassandflushunit.stall_bF$buf8 ),
    .C(_483_),
    .Y(\datapath._06_ [30])
);

INVX1 _10171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [31]),
    .Y(_484_)
);

NAND2X1 _10172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf7 ),
    .B(\datapath.idpc_4 [31]),
    .Y(_485_)
);

OAI21X1 _10173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_484_),
    .B(\bypassandflushunit.stall_bF$buf6 ),
    .C(_485_),
    .Y(\datapath._06_ [31])
);

OR2X2 _10174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [0]),
    .B(\bypassandflushunit.flushalu ),
    .Y(\datapath._28_ [0])
);

OR2X2 _10175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [1]),
    .B(\bypassandflushunit.flushalu ),
    .Y(\datapath._28_ [1])
);

INVX8 _10176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.flushalu ),
    .Y(_486_)
);

AND2X2 _10177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf4),
    .B(\datapath.idinstr [2]),
    .Y(\datapath._28_ [2])
);

AND2X2 _10178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf3),
    .B(\datapath.idinstr [3]),
    .Y(\datapath._28_ [3])
);

OR2X2 _10179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [4]),
    .B(\bypassandflushunit.flushalu ),
    .Y(\datapath._28_ [4])
);

AND2X2 _10180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf2),
    .B(\datapath.idinstr [5]),
    .Y(\datapath._28_ [5])
);

AND2X2 _10181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf1),
    .B(\datapath.idinstr [6]),
    .Y(\datapath._28_ [6])
);

AND2X2 _10182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf0),
    .B(\datapath.idinstr [7]),
    .Y(\datapath._28_ [7])
);

AND2X2 _10183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf4),
    .B(\datapath.idinstr [8]),
    .Y(\datapath._28_ [8])
);

AND2X2 _10184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf3),
    .B(\datapath.idinstr [9]),
    .Y(\datapath._28_ [9])
);

AND2X2 _10185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf2),
    .B(\datapath.idinstr [10]),
    .Y(\datapath._28_ [10])
);

AND2X2 _10186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf1),
    .B(\datapath.idinstr [11]),
    .Y(\datapath._28_ [11])
);

AND2X2 _10187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf0),
    .B(\datapath.idinstr [12]),
    .Y(\datapath._28_ [12])
);

AND2X2 _10188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf4),
    .B(\datapath.idinstr [13]),
    .Y(\datapath._28_ [13])
);

AND2X2 _10189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf3),
    .B(\datapath.idinstr [14]),
    .Y(\datapath._28_ [14])
);

AND2X2 _10190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf2),
    .B(\datapath.idinstr_15_bF$buf53 ),
    .Y(\datapath._28_ [15])
);

AND2X2 _10191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf1),
    .B(\datapath.idinstr_16_bF$buf45 ),
    .Y(\datapath._28_ [16])
);

AND2X2 _10192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf0),
    .B(\datapath.idinstr_17_bF$buf41 ),
    .Y(\datapath._28_ [17])
);

AND2X2 _10193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf4),
    .B(\datapath.idinstr_18_bF$buf7 ),
    .Y(\datapath._28_ [18])
);

AND2X2 _10194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf3),
    .B(\datapath.idinstr_19_bF$buf5 ),
    .Y(\datapath._28_ [19])
);

AND2X2 _10195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf2),
    .B(\datapath.idinstr_20_bF$buf55 ),
    .Y(\datapath._28_ [20])
);

AND2X2 _10196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf1),
    .B(\datapath.idinstr_21_bF$buf44 ),
    .Y(\datapath._28_ [21])
);

AND2X2 _10197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf0),
    .B(\datapath.idinstr_22_bF$buf43 ),
    .Y(\datapath._28_ [22])
);

AND2X2 _10198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf4),
    .B(\datapath.idinstr_23_bF$buf7 ),
    .Y(\datapath._28_ [23])
);

AND2X2 _10199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf3),
    .B(\datapath.idinstr_24_bF$buf5 ),
    .Y(\datapath._28_ [24])
);

AND2X2 _10200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf2),
    .B(\datapath.idinstr [25]),
    .Y(\datapath._28_ [25])
);

AND2X2 _10201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf1),
    .B(\datapath.idinstr [26]),
    .Y(\datapath._28_ [26])
);

AND2X2 _10202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf0),
    .B(\datapath.idinstr [27]),
    .Y(\datapath._28_ [27])
);

AND2X2 _10203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf4),
    .B(\datapath.idinstr [28]),
    .Y(\datapath._28_ [28])
);

AND2X2 _10204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf3),
    .B(\datapath.idinstr [29]),
    .Y(\datapath._28_ [29])
);

AND2X2 _10205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf2),
    .B(\datapath.idinstr [30]),
    .Y(\datapath._28_ [30])
);

AND2X2 _10206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf1),
    .B(\datapath.idinstr [31]),
    .Y(\datapath._28_ [31])
);

AND2X2 _10207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf0),
    .B(\controlunit.ill_op ),
    .Y(\datapath._29_ [0])
);

AND2X2 _10208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf4),
    .B(\controlunit.ebreak ),
    .Y(\datapath._29_ [1])
);

AND2X2 _10209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486__bF$buf3),
    .B(\controlunit.ecall ),
    .Y(\datapath._29_ [2])
);

OR2X2 _10210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.flushid ),
    .B(\datapath.aluinstr [0]),
    .Y(\datapath._30_ [0])
);

OR2X2 _10211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.flushid ),
    .B(\datapath.aluinstr [1]),
    .Y(\datapath._30_ [1])
);

AND2X2 _10212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf4),
    .B(\datapath.aluinstr [2]),
    .Y(\datapath._30_ [2])
);

AND2X2 _10213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf3),
    .B(\datapath.aluinstr [3]),
    .Y(\datapath._30_ [3])
);

OR2X2 _10214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.flushid ),
    .B(\datapath.aluinstr [4]),
    .Y(\datapath._30_ [4])
);

AND2X2 _10215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf2),
    .B(\datapath.aluinstr [5]),
    .Y(\datapath._30_ [5])
);

AND2X2 _10216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf1),
    .B(\datapath.aluinstr [6]),
    .Y(\datapath._30_ [6])
);

AND2X2 _10217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf0),
    .B(\datapath.aluinstr [7]),
    .Y(\datapath._30_ [7])
);

AND2X2 _10218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf4),
    .B(\datapath.aluinstr [8]),
    .Y(\datapath._30_ [8])
);

AND2X2 _10219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf3),
    .B(\datapath.aluinstr [9]),
    .Y(\datapath._30_ [9])
);

AND2X2 _10220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf2),
    .B(\datapath.aluinstr [10]),
    .Y(\datapath._30_ [10])
);

AND2X2 _10221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf1),
    .B(\datapath.aluinstr [11]),
    .Y(\datapath._30_ [11])
);

AND2X2 _10222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf0),
    .B(\datapath.aluinstr [12]),
    .Y(\datapath._30_ [12])
);

AND2X2 _10223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf4),
    .B(\datapath.aluinstr [13]),
    .Y(\datapath._30_ [13])
);

AND2X2 _10224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf3),
    .B(\datapath.aluinstr [14]),
    .Y(\datapath._30_ [14])
);

AND2X2 _10225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf2),
    .B(\datapath.aluinstr [15]),
    .Y(\datapath._30_ [15])
);

AND2X2 _10226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf1),
    .B(\datapath.aluinstr [16]),
    .Y(\datapath._30_ [16])
);

AND2X2 _10227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf0),
    .B(\datapath.aluinstr [17]),
    .Y(\datapath._30_ [17])
);

AND2X2 _10228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf4),
    .B(\datapath.aluinstr [18]),
    .Y(\datapath._30_ [18])
);

AND2X2 _10229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf3),
    .B(\datapath.aluinstr [19]),
    .Y(\datapath._30_ [19])
);

AND2X2 _10230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf2),
    .B(\datapath.aluinstr [20]),
    .Y(\datapath._30_ [20])
);

AND2X2 _10231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf1),
    .B(\datapath.aluinstr [21]),
    .Y(\datapath._30_ [21])
);

AND2X2 _10232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf0),
    .B(\datapath.aluinstr [22]),
    .Y(\datapath._30_ [22])
);

AND2X2 _10233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf4),
    .B(\datapath.aluinstr [23]),
    .Y(\datapath._30_ [23])
);

AND2X2 _10234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf3),
    .B(\datapath.aluinstr [24]),
    .Y(\datapath._30_ [24])
);

AND2X2 _10235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf2),
    .B(\datapath.aluinstr [25]),
    .Y(\datapath._30_ [25])
);

AND2X2 _10236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf1),
    .B(\datapath.aluinstr [26]),
    .Y(\datapath._30_ [26])
);

AND2X2 _10237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf0),
    .B(\datapath.aluinstr [27]),
    .Y(\datapath._30_ [27])
);

AND2X2 _10238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf4),
    .B(\datapath.aluinstr [28]),
    .Y(\datapath._30_ [28])
);

AND2X2 _10239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf3),
    .B(\datapath.aluinstr [29]),
    .Y(\datapath._30_ [29])
);

AND2X2 _10240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf2),
    .B(\datapath.aluinstr [30]),
    .Y(\datapath._30_ [30])
);

AND2X2 _10241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf1),
    .B(\datapath.aluinstr [31]),
    .Y(\datapath._30_ [31])
);

AND2X2 _10242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf0),
    .B(\datapath.aluexecptions [0]),
    .Y(\datapath._31_ [0])
);

AND2X2 _10243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf4),
    .B(\datapath.aluexecptions [1]),
    .Y(\datapath._31_ [1])
);

AND2X2 _10244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf3),
    .B(\datapath.aluexecptions [2]),
    .Y(\datapath._31_ [2])
);

INVX2 _10245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.rs2_bypass_sel [2]),
    .Y(_487_)
);

NOR2X1 _10246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.rs2_bypass_sel [0]),
    .B(\bypassandflushunit.rs2_bypass_sel [1]),
    .Y(_488_)
);

INVX1 _10247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_488_),
    .Y(_489_)
);

NOR2X1 _10248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_),
    .B(_489_),
    .Y(_490_)
);

NAND2X1 _10249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [0]),
    .B(_490__bF$buf4),
    .Y(_491_)
);

INVX1 _10250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.rs2_bypass_sel [0]),
    .Y(_492_)
);

NAND2X1 _10251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.rs2_bypass_sel [1]),
    .B(_487_),
    .Y(_493_)
);

NOR2X1 _10252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_492_),
    .B(_493_),
    .Y(_494_)
);

AOI21X1 _10253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_),
    .B(\bypassandflushunit.rs2_bypass_sel [1]),
    .C(_488_),
    .Y(_495_)
);

AOI22X1 _10254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [0]),
    .B(_495__bF$buf4),
    .C(_494__bF$buf4),
    .D(_0__0_bF$buf4),
    .Y(_496_)
);

NOR2X1 _10255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.rs2_bypass_sel [2]),
    .B(_489_),
    .Y(_497_)
);

NOR2X1 _10256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.rs2_bypass_sel [0]),
    .B(_493_),
    .Y(_498_)
);

AOI22X1 _10257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.condtrue ),
    .B(_498__bF$buf4),
    .C(_497__bF$buf4),
    .D(\datapath.registers.regb_data [0]),
    .Y(_499_)
);

NAND3X1 _10258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_491_),
    .B(_496_),
    .C(_499_),
    .Y(_250_[0])
);

NAND2X1 _10259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [1]),
    .B(_490__bF$buf3),
    .Y(_500_)
);

AOI22X1 _10260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [1]),
    .B(_495__bF$buf3),
    .C(_494__bF$buf3),
    .D(_0__1_bF$buf9),
    .Y(_501_)
);

AOI22X1 _10261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [1]),
    .B(_498__bF$buf3),
    .C(_497__bF$buf3),
    .D(\datapath.registers.regb_data [1]),
    .Y(_502_)
);

NAND3X1 _10262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_500_),
    .B(_501_),
    .C(_502_),
    .Y(_250_[1])
);

NAND2X1 _10263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [2]),
    .B(_490__bF$buf2),
    .Y(_503_)
);

AOI22X1 _10264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [2]),
    .B(_495__bF$buf2),
    .C(_494__bF$buf2),
    .D(_0_[2]),
    .Y(_504_)
);

AOI22X1 _10265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [2]),
    .B(_498__bF$buf2),
    .C(_497__bF$buf2),
    .D(\datapath.registers.regb_data [2]),
    .Y(_505_)
);

NAND3X1 _10266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_503_),
    .B(_504_),
    .C(_505_),
    .Y(_250_[2])
);

NAND2X1 _10267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [3]),
    .B(_490__bF$buf1),
    .Y(_506_)
);

AOI22X1 _10268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [3]),
    .B(_495__bF$buf1),
    .C(_494__bF$buf1),
    .D(_0_[3]),
    .Y(_507_)
);

AOI22X1 _10269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [3]),
    .B(_498__bF$buf1),
    .C(_497__bF$buf1),
    .D(\datapath.registers.regb_data [3]),
    .Y(_508_)
);

NAND3X1 _10270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_506_),
    .B(_507_),
    .C(_508_),
    .Y(_250_[3])
);

NAND2X1 _10271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [4]),
    .B(_490__bF$buf0),
    .Y(_509_)
);

AOI22X1 _10272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [4]),
    .B(_495__bF$buf0),
    .C(_494__bF$buf0),
    .D(_0_[4]),
    .Y(_510_)
);

AOI22X1 _10273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [4]),
    .B(_498__bF$buf0),
    .C(_497__bF$buf0),
    .D(\datapath.registers.regb_data [4]),
    .Y(_511_)
);

NAND3X1 _10274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_509_),
    .B(_510_),
    .C(_511_),
    .Y(_250_[4])
);

NAND2X1 _10275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [5]),
    .B(_490__bF$buf4),
    .Y(_512_)
);

AOI22X1 _10276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [5]),
    .B(_495__bF$buf4),
    .C(_494__bF$buf4),
    .D(_0_[5]),
    .Y(_513_)
);

AOI22X1 _10277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [5]),
    .B(_498__bF$buf4),
    .C(_497__bF$buf4),
    .D(\datapath.registers.regb_data [5]),
    .Y(_514_)
);

NAND3X1 _10278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_512_),
    .B(_513_),
    .C(_514_),
    .Y(_250_[5])
);

NAND2X1 _10279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [6]),
    .B(_490__bF$buf3),
    .Y(_515_)
);

AOI22X1 _10280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [6]),
    .B(_495__bF$buf3),
    .C(_494__bF$buf3),
    .D(_0_[6]),
    .Y(_516_)
);

AOI22X1 _10281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [6]),
    .B(_498__bF$buf3),
    .C(_497__bF$buf3),
    .D(\datapath.registers.regb_data [6]),
    .Y(_517_)
);

NAND3X1 _10282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_515_),
    .B(_516_),
    .C(_517_),
    .Y(_250_[6])
);

NAND2X1 _10283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [7]),
    .B(_490__bF$buf2),
    .Y(_518_)
);

AOI22X1 _10284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [7]),
    .B(_495__bF$buf2),
    .C(_494__bF$buf2),
    .D(_0_[7]),
    .Y(_519_)
);

AOI22X1 _10285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [7]),
    .B(_498__bF$buf2),
    .C(_497__bF$buf2),
    .D(\datapath.registers.regb_data [7]),
    .Y(_520_)
);

NAND3X1 _10286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_518_),
    .B(_519_),
    .C(_520_),
    .Y(_250_[7])
);

NAND2X1 _10287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [8]),
    .B(_490__bF$buf1),
    .Y(_521_)
);

AOI22X1 _10288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [8]),
    .B(_495__bF$buf1),
    .C(_494__bF$buf1),
    .D(_0_[8]),
    .Y(_522_)
);

AOI22X1 _10289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [8]),
    .B(_498__bF$buf1),
    .C(_497__bF$buf1),
    .D(\datapath.registers.regb_data [8]),
    .Y(_523_)
);

NAND3X1 _10290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_521_),
    .B(_522_),
    .C(_523_),
    .Y(_250_[8])
);

NAND2X1 _10291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [9]),
    .B(_490__bF$buf0),
    .Y(_524_)
);

AOI22X1 _10292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [9]),
    .B(_495__bF$buf0),
    .C(_494__bF$buf0),
    .D(_0_[9]),
    .Y(_525_)
);

AOI22X1 _10293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [9]),
    .B(_498__bF$buf0),
    .C(_497__bF$buf0),
    .D(\datapath.registers.regb_data [9]),
    .Y(_526_)
);

NAND3X1 _10294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_524_),
    .B(_525_),
    .C(_526_),
    .Y(_250_[9])
);

NAND2X1 _10295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [10]),
    .B(_490__bF$buf4),
    .Y(_527_)
);

AOI22X1 _10296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [10]),
    .B(_495__bF$buf4),
    .C(_494__bF$buf4),
    .D(_0_[10]),
    .Y(_528_)
);

AOI22X1 _10297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [10]),
    .B(_498__bF$buf4),
    .C(_497__bF$buf4),
    .D(\datapath.registers.regb_data [10]),
    .Y(_529_)
);

NAND3X1 _10298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_527_),
    .B(_528_),
    .C(_529_),
    .Y(_250_[10])
);

NAND2X1 _10299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [11]),
    .B(_490__bF$buf3),
    .Y(_530_)
);

AOI22X1 _10300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [11]),
    .B(_495__bF$buf3),
    .C(_494__bF$buf3),
    .D(_0_[11]),
    .Y(_531_)
);

AOI22X1 _10301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [11]),
    .B(_498__bF$buf3),
    .C(_497__bF$buf3),
    .D(\datapath.registers.regb_data [11]),
    .Y(_532_)
);

NAND3X1 _10302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_530_),
    .B(_531_),
    .C(_532_),
    .Y(_250_[11])
);

NAND2X1 _10303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [12]),
    .B(_490__bF$buf2),
    .Y(_533_)
);

AOI22X1 _10304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [12]),
    .B(_495__bF$buf2),
    .C(_494__bF$buf2),
    .D(_0_[12]),
    .Y(_534_)
);

AOI22X1 _10305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [12]),
    .B(_498__bF$buf2),
    .C(_497__bF$buf2),
    .D(\datapath.registers.regb_data [12]),
    .Y(_535_)
);

NAND3X1 _10306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_533_),
    .B(_534_),
    .C(_535_),
    .Y(_250_[12])
);

NAND2X1 _10307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [13]),
    .B(_490__bF$buf1),
    .Y(_536_)
);

AOI22X1 _10308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [13]),
    .B(_495__bF$buf1),
    .C(_494__bF$buf1),
    .D(_0_[13]),
    .Y(_537_)
);

AOI22X1 _10309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [13]),
    .B(_498__bF$buf1),
    .C(_497__bF$buf1),
    .D(\datapath.registers.regb_data [13]),
    .Y(_538_)
);

NAND3X1 _10310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_536_),
    .B(_537_),
    .C(_538_),
    .Y(_250_[13])
);

NAND2X1 _10311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [14]),
    .B(_490__bF$buf0),
    .Y(_539_)
);

AOI22X1 _10312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [14]),
    .B(_495__bF$buf0),
    .C(_494__bF$buf0),
    .D(_0_[14]),
    .Y(_540_)
);

AOI22X1 _10313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [14]),
    .B(_498__bF$buf0),
    .C(_497__bF$buf0),
    .D(\datapath.registers.regb_data [14]),
    .Y(_541_)
);

NAND3X1 _10314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_539_),
    .B(_540_),
    .C(_541_),
    .Y(_250_[14])
);

NAND2X1 _10315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [15]),
    .B(_490__bF$buf4),
    .Y(_542_)
);

AOI22X1 _10316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [15]),
    .B(_495__bF$buf4),
    .C(_494__bF$buf4),
    .D(_0_[15]),
    .Y(_543_)
);

AOI22X1 _10317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [15]),
    .B(_498__bF$buf4),
    .C(_497__bF$buf4),
    .D(\datapath.registers.regb_data [15]),
    .Y(_544_)
);

NAND3X1 _10318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_542_),
    .B(_543_),
    .C(_544_),
    .Y(_250_[15])
);

NAND2X1 _10319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [16]),
    .B(_490__bF$buf3),
    .Y(_545_)
);

AOI22X1 _10320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [16]),
    .B(_495__bF$buf3),
    .C(_494__bF$buf3),
    .D(_0_[16]),
    .Y(_546_)
);

AOI22X1 _10321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [16]),
    .B(_498__bF$buf3),
    .C(_497__bF$buf3),
    .D(\datapath.registers.regb_data [16]),
    .Y(_547_)
);

NAND3X1 _10322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_545_),
    .B(_546_),
    .C(_547_),
    .Y(_250_[16])
);

NAND2X1 _10323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [17]),
    .B(_490__bF$buf2),
    .Y(_548_)
);

AOI22X1 _10324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [17]),
    .B(_495__bF$buf2),
    .C(_494__bF$buf2),
    .D(_0_[17]),
    .Y(_549_)
);

AOI22X1 _10325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [17]),
    .B(_498__bF$buf2),
    .C(_497__bF$buf2),
    .D(\datapath.registers.regb_data [17]),
    .Y(_550_)
);

NAND3X1 _10326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_548_),
    .B(_549_),
    .C(_550_),
    .Y(_250_[17])
);

NAND2X1 _10327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [18]),
    .B(_490__bF$buf1),
    .Y(_551_)
);

AOI22X1 _10328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [18]),
    .B(_495__bF$buf1),
    .C(_494__bF$buf1),
    .D(_0_[18]),
    .Y(_552_)
);

AOI22X1 _10329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [18]),
    .B(_498__bF$buf1),
    .C(_497__bF$buf1),
    .D(\datapath.registers.regb_data [18]),
    .Y(_553_)
);

NAND3X1 _10330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_551_),
    .B(_552_),
    .C(_553_),
    .Y(_250_[18])
);

NAND2X1 _10331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [19]),
    .B(_490__bF$buf0),
    .Y(_554_)
);

AOI22X1 _10332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [19]),
    .B(_495__bF$buf0),
    .C(_494__bF$buf0),
    .D(_0_[19]),
    .Y(_555_)
);

AOI22X1 _10333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [19]),
    .B(_498__bF$buf0),
    .C(_497__bF$buf0),
    .D(\datapath.registers.regb_data [19]),
    .Y(_556_)
);

NAND3X1 _10334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_554_),
    .B(_555_),
    .C(_556_),
    .Y(_250_[19])
);

NAND2X1 _10335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [20]),
    .B(_490__bF$buf4),
    .Y(_557_)
);

AOI22X1 _10336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [20]),
    .B(_495__bF$buf4),
    .C(_494__bF$buf4),
    .D(_0_[20]),
    .Y(_558_)
);

AOI22X1 _10337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [20]),
    .B(_498__bF$buf4),
    .C(_497__bF$buf4),
    .D(\datapath.registers.regb_data [20]),
    .Y(_559_)
);

NAND3X1 _10338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_557_),
    .B(_558_),
    .C(_559_),
    .Y(_250_[20])
);

NAND2X1 _10339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [21]),
    .B(_490__bF$buf3),
    .Y(_560_)
);

AOI22X1 _10340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [21]),
    .B(_495__bF$buf3),
    .C(_494__bF$buf3),
    .D(_0_[21]),
    .Y(_561_)
);

AOI22X1 _10341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [21]),
    .B(_498__bF$buf3),
    .C(_497__bF$buf3),
    .D(\datapath.registers.regb_data [21]),
    .Y(_562_)
);

NAND3X1 _10342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_560_),
    .B(_561_),
    .C(_562_),
    .Y(_250_[21])
);

NAND2X1 _10343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [22]),
    .B(_490__bF$buf2),
    .Y(_563_)
);

AOI22X1 _10344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [22]),
    .B(_495__bF$buf2),
    .C(_494__bF$buf2),
    .D(_0_[22]),
    .Y(_564_)
);

AOI22X1 _10345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [22]),
    .B(_498__bF$buf2),
    .C(_497__bF$buf2),
    .D(\datapath.registers.regb_data [22]),
    .Y(_565_)
);

NAND3X1 _10346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_563_),
    .B(_564_),
    .C(_565_),
    .Y(_250_[22])
);

NAND2X1 _10347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [23]),
    .B(_490__bF$buf1),
    .Y(_566_)
);

AOI22X1 _10348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [23]),
    .B(_495__bF$buf1),
    .C(_494__bF$buf1),
    .D(_0_[23]),
    .Y(_567_)
);

AOI22X1 _10349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [23]),
    .B(_498__bF$buf1),
    .C(_497__bF$buf1),
    .D(\datapath.registers.regb_data [23]),
    .Y(_568_)
);

NAND3X1 _10350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_566_),
    .B(_567_),
    .C(_568_),
    .Y(_250_[23])
);

NAND2X1 _10351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [24]),
    .B(_490__bF$buf0),
    .Y(_569_)
);

AOI22X1 _10352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [24]),
    .B(_495__bF$buf0),
    .C(_494__bF$buf0),
    .D(_0_[24]),
    .Y(_570_)
);

AOI22X1 _10353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [24]),
    .B(_498__bF$buf0),
    .C(_497__bF$buf0),
    .D(\datapath.registers.regb_data [24]),
    .Y(_571_)
);

NAND3X1 _10354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_569_),
    .B(_570_),
    .C(_571_),
    .Y(_250_[24])
);

NAND2X1 _10355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [25]),
    .B(_490__bF$buf4),
    .Y(_572_)
);

AOI22X1 _10356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [25]),
    .B(_495__bF$buf4),
    .C(_494__bF$buf4),
    .D(_0_[25]),
    .Y(_573_)
);

AOI22X1 _10357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [25]),
    .B(_498__bF$buf4),
    .C(_497__bF$buf4),
    .D(\datapath.registers.regb_data [25]),
    .Y(_574_)
);

NAND3X1 _10358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_572_),
    .B(_573_),
    .C(_574_),
    .Y(_250_[25])
);

NAND2X1 _10359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [26]),
    .B(_490__bF$buf3),
    .Y(_575_)
);

AOI22X1 _10360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [26]),
    .B(_495__bF$buf3),
    .C(_494__bF$buf3),
    .D(_0_[26]),
    .Y(_576_)
);

AOI22X1 _10361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [26]),
    .B(_498__bF$buf3),
    .C(_497__bF$buf3),
    .D(\datapath.registers.regb_data [26]),
    .Y(_577_)
);

NAND3X1 _10362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_575_),
    .B(_576_),
    .C(_577_),
    .Y(_250_[26])
);

NAND2X1 _10363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [27]),
    .B(_490__bF$buf2),
    .Y(_578_)
);

AOI22X1 _10364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [27]),
    .B(_495__bF$buf2),
    .C(_494__bF$buf2),
    .D(_0_[27]),
    .Y(_579_)
);

AOI22X1 _10365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [27]),
    .B(_498__bF$buf2),
    .C(_497__bF$buf2),
    .D(\datapath.registers.regb_data [27]),
    .Y(_580_)
);

NAND3X1 _10366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_578_),
    .B(_579_),
    .C(_580_),
    .Y(_250_[27])
);

NAND2X1 _10367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [28]),
    .B(_490__bF$buf1),
    .Y(_581_)
);

AOI22X1 _10368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [28]),
    .B(_495__bF$buf1),
    .C(_494__bF$buf1),
    .D(_0_[28]),
    .Y(_582_)
);

AOI22X1 _10369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [28]),
    .B(_498__bF$buf1),
    .C(_497__bF$buf1),
    .D(\datapath.registers.regb_data [28]),
    .Y(_583_)
);

NAND3X1 _10370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_581_),
    .B(_582_),
    .C(_583_),
    .Y(_250_[28])
);

NAND2X1 _10371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [29]),
    .B(_490__bF$buf0),
    .Y(_584_)
);

AOI22X1 _10372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [29]),
    .B(_495__bF$buf0),
    .C(_494__bF$buf0),
    .D(_0_[29]),
    .Y(_585_)
);

AOI22X1 _10373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [29]),
    .B(_498__bF$buf0),
    .C(_497__bF$buf0),
    .D(\datapath.registers.regb_data [29]),
    .Y(_586_)
);

NAND3X1 _10374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_584_),
    .B(_585_),
    .C(_586_),
    .Y(_250_[29])
);

NAND2X1 _10375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [30]),
    .B(_490__bF$buf4),
    .Y(_587_)
);

AOI22X1 _10376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [30]),
    .B(_495__bF$buf4),
    .C(_494__bF$buf4),
    .D(_0_[30]),
    .Y(_588_)
);

AOI22X1 _10377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [30]),
    .B(_498__bF$buf4),
    .C(_497__bF$buf4),
    .D(\datapath.registers.regb_data [30]),
    .Y(_589_)
);

NAND3X1 _10378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_587_),
    .B(_588_),
    .C(_589_),
    .Y(_250_[30])
);

NAND2X1 _10379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [31]),
    .B(_490__bF$buf3),
    .Y(_590_)
);

AOI22X1 _10380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [31]),
    .B(_495__bF$buf3),
    .C(_494__bF$buf3),
    .D(_0_[31]),
    .Y(_591_)
);

AOI22X1 _10381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [31]),
    .B(_498__bF$buf3),
    .C(_497__bF$buf3),
    .D(\datapath.registers.regb_data [31]),
    .Y(_592_)
);

NAND3X1 _10382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_590_),
    .B(_591_),
    .C(_592_),
    .Y(_250_[31])
);

INVX1 _10383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [0]),
    .Y(_593_)
);

INVX1 _10384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bsel[0]),
    .Y(_594_)
);

AND2X2 _10385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_594_),
    .B(bsel[1]),
    .Y(_595_)
);

NOR2X1 _10386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bsel[1]),
    .B(_594_),
    .Y(_596_)
);

NOR2X1 _10387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_596__bF$buf4),
    .B(_595__bF$buf4),
    .Y(_597_)
);

NAND2X1 _10388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_593_),
    .B(_597__bF$buf4),
    .Y(_598_)
);

INVX1 _10389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.immediatedecoder._06_ ),
    .Y(_599_)
);

NAND2X1 _10390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_599_),
    .B(_596__bF$buf3),
    .Y(_600_)
);

INVX1 _10391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [0]),
    .Y(_601_)
);

INVX1 _10392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bbpsel[2]),
    .Y(_602_)
);

NOR2X1 _10393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bbpsel[0]),
    .B(bbpsel[1]),
    .Y(_603_)
);

NAND2X1 _10394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_602_),
    .B(_603_),
    .Y(_604_)
);

AOI21X1 _10395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_601_),
    .B(_595__bF$buf3),
    .C(_604__bF$buf4),
    .Y(_605_)
);

NAND3X1 _10396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_600_),
    .B(_605_),
    .C(_598_),
    .Y(_606_)
);

INVX1 _10397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bbpsel[1]),
    .Y(_607_)
);

NOR2X1 _10398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bbpsel[2]),
    .B(_607_),
    .Y(_608_)
);

AND2X2 _10399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_608_),
    .B(bbpsel[0]),
    .Y(_609_)
);

INVX1 _10400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_603_),
    .Y(_610_)
);

NOR2X1 _10401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_602_),
    .B(_610_),
    .Y(_611_)
);

AOI22X1 _10402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [0]),
    .B(_611__bF$buf4),
    .C(_609__bF$buf4),
    .D(_0__0_bF$buf3),
    .Y(_612_)
);

INVX1 _10403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [0]),
    .Y(_613_)
);

OAI21X1 _10404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bbpsel[2]),
    .B(_607_),
    .C(_610_),
    .Y(_614_)
);

NOR2X1 _10405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_613_),
    .B(_614__bF$buf4),
    .Y(_615_)
);

INVX1 _10406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_608_),
    .Y(_616_)
);

NOR2X1 _10407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bbpsel[0]),
    .B(_616_),
    .Y(_617_)
);

AOI21X1 _10408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.condtrue ),
    .B(_617__bF$buf4),
    .C(_615_),
    .Y(_618_)
);

NAND3X1 _10409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_612_),
    .B(_618_),
    .C(_606_),
    .Y(_249_[0])
);

INVX1 _10410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [1]),
    .Y(_619_)
);

NAND2X1 _10411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_619_),
    .B(_597__bF$buf3),
    .Y(_620_)
);

INVX1 _10412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [1]),
    .Y(_621_)
);

NAND2X1 _10413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_621_),
    .B(_596__bF$buf2),
    .Y(_622_)
);

INVX1 _10414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [1]),
    .Y(_623_)
);

AOI21X1 _10415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_623_),
    .B(_595__bF$buf2),
    .C(_604__bF$buf3),
    .Y(_624_)
);

NAND3X1 _10416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_622_),
    .B(_624_),
    .C(_620_),
    .Y(_625_)
);

AOI22X1 _10417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [1]),
    .B(_611__bF$buf3),
    .C(_617__bF$buf3),
    .D(\datapath.alu.c [1]),
    .Y(_626_)
);

INVX1 _10418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [1]),
    .Y(_627_)
);

NOR2X1 _10419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_627_),
    .B(_614__bF$buf3),
    .Y(_628_)
);

AOI21X1 _10420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf8),
    .B(_609__bF$buf3),
    .C(_628_),
    .Y(_629_)
);

NAND3X1 _10421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_626_),
    .B(_629_),
    .C(_625_),
    .Y(_249_[1])
);

INVX1 _10422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [2]),
    .Y(_630_)
);

NAND2X1 _10423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_630_),
    .B(_597__bF$buf2),
    .Y(_631_)
);

INVX1 _10424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [2]),
    .Y(_632_)
);

NAND2X1 _10425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_632_),
    .B(_596__bF$buf1),
    .Y(_633_)
);

INVX1 _10426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [2]),
    .Y(_634_)
);

AOI21X1 _10427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_634_),
    .B(_595__bF$buf1),
    .C(_604__bF$buf2),
    .Y(_635_)
);

NAND3X1 _10428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_633_),
    .B(_635_),
    .C(_631_),
    .Y(_636_)
);

AOI22X1 _10429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [2]),
    .B(_611__bF$buf2),
    .C(_609__bF$buf2),
    .D(_0_[2]),
    .Y(_637_)
);

INVX1 _10430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [2]),
    .Y(_638_)
);

NOR2X1 _10431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_638_),
    .B(_614__bF$buf2),
    .Y(_639_)
);

AOI21X1 _10432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [2]),
    .B(_617__bF$buf2),
    .C(_639_),
    .Y(_640_)
);

NAND3X1 _10433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_637_),
    .B(_640_),
    .C(_636_),
    .Y(_249_[2])
);

INVX1 _10434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [3]),
    .Y(_641_)
);

NAND2X1 _10435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_641_),
    .B(_597__bF$buf1),
    .Y(_642_)
);

INVX1 _10436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [3]),
    .Y(_643_)
);

NAND2X1 _10437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_643_),
    .B(_596__bF$buf0),
    .Y(_644_)
);

INVX1 _10438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [3]),
    .Y(_645_)
);

AOI21X1 _10439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_645_),
    .B(_595__bF$buf0),
    .C(_604__bF$buf1),
    .Y(_646_)
);

NAND3X1 _10440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_644_),
    .B(_646_),
    .C(_642_),
    .Y(_647_)
);

AOI22X1 _10441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [3]),
    .B(_611__bF$buf1),
    .C(_617__bF$buf1),
    .D(\datapath.alu.c [3]),
    .Y(_648_)
);

INVX1 _10442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [3]),
    .Y(_649_)
);

NOR2X1 _10443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_649_),
    .B(_614__bF$buf1),
    .Y(_650_)
);

AOI21X1 _10444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[3]),
    .B(_609__bF$buf1),
    .C(_650_),
    .Y(_651_)
);

NAND3X1 _10445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_648_),
    .B(_651_),
    .C(_647_),
    .Y(_249_[3])
);

INVX1 _10446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [4]),
    .Y(_652_)
);

NAND2X1 _10447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_652_),
    .B(_597__bF$buf0),
    .Y(_653_)
);

INVX1 _10448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [4]),
    .Y(_654_)
);

NAND2X1 _10449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_654_),
    .B(_596__bF$buf4),
    .Y(_655_)
);

INVX1 _10450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [4]),
    .Y(_656_)
);

AOI21X1 _10451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_656_),
    .B(_595__bF$buf4),
    .C(_604__bF$buf0),
    .Y(_657_)
);

NAND3X1 _10452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_655_),
    .B(_657_),
    .C(_653_),
    .Y(_658_)
);

AOI22X1 _10453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [4]),
    .B(_611__bF$buf0),
    .C(_617__bF$buf0),
    .D(\datapath.alu.c [4]),
    .Y(_659_)
);

INVX1 _10454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [4]),
    .Y(_660_)
);

NOR2X1 _10455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_660_),
    .B(_614__bF$buf0),
    .Y(_661_)
);

AOI21X1 _10456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[4]),
    .B(_609__bF$buf0),
    .C(_661_),
    .Y(_662_)
);

NAND3X1 _10457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_659_),
    .B(_662_),
    .C(_658_),
    .Y(_249_[4])
);

INVX1 _10458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [5]),
    .Y(_663_)
);

NAND2X1 _10459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_663_),
    .B(_597__bF$buf4),
    .Y(_664_)
);

INVX1 _10460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [5]),
    .Y(_665_)
);

NAND2X1 _10461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_665_),
    .B(_596__bF$buf3),
    .Y(_666_)
);

INVX1 _10462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [5]),
    .Y(_667_)
);

AOI21X1 _10463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_667_),
    .B(_595__bF$buf3),
    .C(_604__bF$buf4),
    .Y(_668_)
);

NAND3X1 _10464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_666_),
    .B(_668_),
    .C(_664_),
    .Y(_669_)
);

AOI22X1 _10465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [5]),
    .B(_611__bF$buf4),
    .C(_617__bF$buf4),
    .D(\datapath.alu.c [5]),
    .Y(_670_)
);

INVX1 _10466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [5]),
    .Y(_671_)
);

NOR2X1 _10467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_671_),
    .B(_614__bF$buf4),
    .Y(_672_)
);

AOI21X1 _10468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[5]),
    .B(_609__bF$buf4),
    .C(_672_),
    .Y(_673_)
);

NAND3X1 _10469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_670_),
    .B(_673_),
    .C(_669_),
    .Y(_249_[5])
);

INVX1 _10470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [6]),
    .Y(_674_)
);

NAND2X1 _10471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_674_),
    .B(_597__bF$buf3),
    .Y(_675_)
);

INVX1 _10472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [6]),
    .Y(_676_)
);

NAND2X1 _10473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_676_),
    .B(_596__bF$buf2),
    .Y(_677_)
);

INVX1 _10474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [6]),
    .Y(_678_)
);

AOI21X1 _10475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_678_),
    .B(_595__bF$buf2),
    .C(_604__bF$buf3),
    .Y(_679_)
);

NAND3X1 _10476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_677_),
    .B(_679_),
    .C(_675_),
    .Y(_680_)
);

AOI22X1 _10477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [6]),
    .B(_611__bF$buf3),
    .C(_609__bF$buf3),
    .D(_0_[6]),
    .Y(_681_)
);

INVX1 _10478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [6]),
    .Y(_682_)
);

NOR2X1 _10479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_682_),
    .B(_614__bF$buf3),
    .Y(_683_)
);

AOI21X1 _10480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [6]),
    .B(_617__bF$buf3),
    .C(_683_),
    .Y(_684_)
);

NAND3X1 _10481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_681_),
    .B(_684_),
    .C(_680_),
    .Y(_249_[6])
);

INVX1 _10482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [7]),
    .Y(_685_)
);

NAND2X1 _10483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_685_),
    .B(_597__bF$buf2),
    .Y(_686_)
);

INVX1 _10484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [7]),
    .Y(_687_)
);

NAND2X1 _10485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_687_),
    .B(_596__bF$buf1),
    .Y(_688_)
);

INVX1 _10486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [7]),
    .Y(_689_)
);

AOI21X1 _10487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_689_),
    .B(_595__bF$buf1),
    .C(_604__bF$buf2),
    .Y(_690_)
);

NAND3X1 _10488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_688_),
    .B(_690_),
    .C(_686_),
    .Y(_691_)
);

AOI22X1 _10489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [7]),
    .B(_611__bF$buf2),
    .C(_609__bF$buf2),
    .D(_0_[7]),
    .Y(_692_)
);

INVX1 _10490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [7]),
    .Y(_693_)
);

NOR2X1 _10491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_693_),
    .B(_614__bF$buf2),
    .Y(_694_)
);

AOI21X1 _10492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [7]),
    .B(_617__bF$buf2),
    .C(_694_),
    .Y(_695_)
);

NAND3X1 _10493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_692_),
    .B(_695_),
    .C(_691_),
    .Y(_249_[7])
);

INVX1 _10494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [8]),
    .Y(_696_)
);

NAND2X1 _10495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_696_),
    .B(_597__bF$buf1),
    .Y(_697_)
);

INVX1 _10496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [8]),
    .Y(_698_)
);

NAND2X1 _10497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_698_),
    .B(_596__bF$buf0),
    .Y(_699_)
);

INVX1 _10498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [8]),
    .Y(_700_)
);

AOI21X1 _10499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_700_),
    .B(_595__bF$buf0),
    .C(_604__bF$buf1),
    .Y(_701_)
);

NAND3X1 _10500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_699_),
    .B(_701_),
    .C(_697_),
    .Y(_702_)
);

AOI22X1 _10501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [8]),
    .B(_611__bF$buf1),
    .C(_617__bF$buf1),
    .D(\datapath.alu.c [8]),
    .Y(_703_)
);

INVX1 _10502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [8]),
    .Y(_704_)
);

NOR2X1 _10503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_704_),
    .B(_614__bF$buf1),
    .Y(_705_)
);

AOI21X1 _10504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[8]),
    .B(_609__bF$buf1),
    .C(_705_),
    .Y(_706_)
);

NAND3X1 _10505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_703_),
    .B(_706_),
    .C(_702_),
    .Y(_249_[8])
);

INVX1 _10506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [9]),
    .Y(_707_)
);

NAND2X1 _10507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_707_),
    .B(_597__bF$buf0),
    .Y(_708_)
);

INVX1 _10508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [9]),
    .Y(_709_)
);

NAND2X1 _10509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_709_),
    .B(_596__bF$buf4),
    .Y(_710_)
);

INVX1 _10510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [9]),
    .Y(_711_)
);

AOI21X1 _10511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_711_),
    .B(_595__bF$buf4),
    .C(_604__bF$buf0),
    .Y(_712_)
);

NAND3X1 _10512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_710_),
    .B(_712_),
    .C(_708_),
    .Y(_713_)
);

AOI22X1 _10513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [9]),
    .B(_611__bF$buf0),
    .C(_609__bF$buf0),
    .D(_0_[9]),
    .Y(_714_)
);

INVX1 _10514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [9]),
    .Y(_715_)
);

NOR2X1 _10515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_715_),
    .B(_614__bF$buf0),
    .Y(_716_)
);

AOI21X1 _10516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [9]),
    .B(_617__bF$buf0),
    .C(_716_),
    .Y(_717_)
);

NAND3X1 _10517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_714_),
    .B(_717_),
    .C(_713_),
    .Y(_249_[9])
);

INVX1 _10518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [10]),
    .Y(_718_)
);

NAND2X1 _10519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_718_),
    .B(_597__bF$buf4),
    .Y(_719_)
);

INVX1 _10520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [10]),
    .Y(_720_)
);

NAND2X1 _10521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_720_),
    .B(_596__bF$buf3),
    .Y(_721_)
);

INVX1 _10522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [10]),
    .Y(_722_)
);

AOI21X1 _10523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_722_),
    .B(_595__bF$buf3),
    .C(_604__bF$buf4),
    .Y(_723_)
);

NAND3X1 _10524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_721_),
    .B(_723_),
    .C(_719_),
    .Y(_724_)
);

AOI22X1 _10525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [10]),
    .B(_611__bF$buf4),
    .C(_609__bF$buf4),
    .D(_0_[10]),
    .Y(_725_)
);

INVX1 _10526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [10]),
    .Y(_726_)
);

NOR2X1 _10527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_726_),
    .B(_614__bF$buf4),
    .Y(_727_)
);

AOI21X1 _10528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [10]),
    .B(_617__bF$buf4),
    .C(_727_),
    .Y(_728_)
);

NAND3X1 _10529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_725_),
    .B(_728_),
    .C(_724_),
    .Y(_249_[10])
);

INVX1 _10530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [11]),
    .Y(_729_)
);

NAND2X1 _10531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_729_),
    .B(_597__bF$buf3),
    .Y(_730_)
);

INVX1 _10532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.immediatedecoder._09_ ),
    .Y(_731_)
);

NAND2X1 _10533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_731_),
    .B(_596__bF$buf2),
    .Y(_732_)
);

INVX1 _10534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [11]),
    .Y(_733_)
);

AOI21X1 _10535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_733_),
    .B(_595__bF$buf2),
    .C(_604__bF$buf3),
    .Y(_734_)
);

NAND3X1 _10536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_732_),
    .B(_734_),
    .C(_730_),
    .Y(_735_)
);

AOI22X1 _10537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [11]),
    .B(_611__bF$buf3),
    .C(_609__bF$buf3),
    .D(_0_[11]),
    .Y(_736_)
);

INVX1 _10538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [11]),
    .Y(_737_)
);

NOR2X1 _10539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_737_),
    .B(_614__bF$buf3),
    .Y(_738_)
);

AOI21X1 _10540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [11]),
    .B(_617__bF$buf3),
    .C(_738_),
    .Y(_739_)
);

NAND3X1 _10541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_736_),
    .B(_739_),
    .C(_735_),
    .Y(_249_[11])
);

INVX1 _10542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [12]),
    .Y(_740_)
);

NAND2X1 _10543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_740_),
    .B(_597__bF$buf2),
    .Y(_741_)
);

INVX1 _10544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [12]),
    .Y(_742_)
);

NAND2X1 _10545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_742_),
    .B(_596__bF$buf1),
    .Y(_743_)
);

INVX1 _10546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [12]),
    .Y(_744_)
);

AOI21X1 _10547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_744_),
    .B(_595__bF$buf1),
    .C(_604__bF$buf2),
    .Y(_745_)
);

NAND3X1 _10548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_743_),
    .B(_745_),
    .C(_741_),
    .Y(_746_)
);

AOI22X1 _10549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [12]),
    .B(_611__bF$buf2),
    .C(_609__bF$buf2),
    .D(_0_[12]),
    .Y(_747_)
);

INVX1 _10550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [12]),
    .Y(_748_)
);

NOR2X1 _10551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_748_),
    .B(_614__bF$buf2),
    .Y(_749_)
);

AOI21X1 _10552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [12]),
    .B(_617__bF$buf2),
    .C(_749_),
    .Y(_750_)
);

NAND3X1 _10553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_747_),
    .B(_750_),
    .C(_746_),
    .Y(_249_[12])
);

INVX1 _10554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [13]),
    .Y(_751_)
);

NAND2X1 _10555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_751_),
    .B(_597__bF$buf1),
    .Y(_752_)
);

INVX1 _10556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [13]),
    .Y(_753_)
);

NAND2X1 _10557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_753_),
    .B(_596__bF$buf0),
    .Y(_754_)
);

INVX1 _10558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [13]),
    .Y(_755_)
);

AOI21X1 _10559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_),
    .B(_595__bF$buf0),
    .C(_604__bF$buf1),
    .Y(_756_)
);

NAND3X1 _10560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_754_),
    .B(_756_),
    .C(_752_),
    .Y(_757_)
);

AOI22X1 _10561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [13]),
    .B(_611__bF$buf1),
    .C(_617__bF$buf1),
    .D(\datapath.alu.c [13]),
    .Y(_758_)
);

INVX1 _10562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [13]),
    .Y(_759_)
);

NOR2X1 _10563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_759_),
    .B(_614__bF$buf1),
    .Y(_760_)
);

AOI21X1 _10564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[13]),
    .B(_609__bF$buf1),
    .C(_760_),
    .Y(_761_)
);

NAND3X1 _10565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_758_),
    .B(_761_),
    .C(_757_),
    .Y(_249_[13])
);

INVX1 _10566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [14]),
    .Y(_762_)
);

NAND2X1 _10567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_762_),
    .B(_597__bF$buf0),
    .Y(_763_)
);

INVX1 _10568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [14]),
    .Y(_764_)
);

NAND2X1 _10569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_764_),
    .B(_596__bF$buf4),
    .Y(_765_)
);

INVX1 _10570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [14]),
    .Y(_766_)
);

AOI21X1 _10571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_766_),
    .B(_595__bF$buf4),
    .C(_604__bF$buf0),
    .Y(_767_)
);

NAND3X1 _10572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_765_),
    .B(_767_),
    .C(_763_),
    .Y(_768_)
);

AOI22X1 _10573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [14]),
    .B(_611__bF$buf0),
    .C(_609__bF$buf0),
    .D(_0_[14]),
    .Y(_769_)
);

INVX1 _10574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [14]),
    .Y(_770_)
);

NOR2X1 _10575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_770_),
    .B(_614__bF$buf0),
    .Y(_771_)
);

AOI21X1 _10576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [14]),
    .B(_617__bF$buf0),
    .C(_771_),
    .Y(_772_)
);

NAND3X1 _10577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_769_),
    .B(_772_),
    .C(_768_),
    .Y(_249_[14])
);

INVX1 _10578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [15]),
    .Y(_773_)
);

NAND2X1 _10579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_773_),
    .B(_597__bF$buf4),
    .Y(_774_)
);

INVX1 _10580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [15]),
    .Y(_775_)
);

NAND2X1 _10581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_775_),
    .B(_596__bF$buf3),
    .Y(_776_)
);

INVX1 _10582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [15]),
    .Y(_777_)
);

AOI21X1 _10583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_777_),
    .B(_595__bF$buf3),
    .C(_604__bF$buf4),
    .Y(_778_)
);

NAND3X1 _10584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_776_),
    .B(_778_),
    .C(_774_),
    .Y(_779_)
);

AOI22X1 _10585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [15]),
    .B(_611__bF$buf4),
    .C(_609__bF$buf4),
    .D(_0_[15]),
    .Y(_780_)
);

INVX1 _10586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [15]),
    .Y(_781_)
);

NOR2X1 _10587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_781_),
    .B(_614__bF$buf4),
    .Y(_782_)
);

AOI21X1 _10588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [15]),
    .B(_617__bF$buf4),
    .C(_782_),
    .Y(_783_)
);

NAND3X1 _10589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_780_),
    .B(_783_),
    .C(_779_),
    .Y(_249_[15])
);

INVX1 _10590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [16]),
    .Y(_784_)
);

NAND2X1 _10591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_784_),
    .B(_597__bF$buf3),
    .Y(_785_)
);

INVX1 _10592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [16]),
    .Y(_786_)
);

NAND2X1 _10593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_786_),
    .B(_596__bF$buf2),
    .Y(_787_)
);

INVX1 _10594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [16]),
    .Y(_788_)
);

AOI21X1 _10595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_788_),
    .B(_595__bF$buf2),
    .C(_604__bF$buf3),
    .Y(_789_)
);

NAND3X1 _10596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_787_),
    .B(_789_),
    .C(_785_),
    .Y(_790_)
);

AOI22X1 _10597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [16]),
    .B(_611__bF$buf3),
    .C(_609__bF$buf3),
    .D(_0_[16]),
    .Y(_791_)
);

INVX1 _10598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [16]),
    .Y(_792_)
);

NOR2X1 _10599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_792_),
    .B(_614__bF$buf3),
    .Y(_793_)
);

AOI21X1 _10600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [16]),
    .B(_617__bF$buf3),
    .C(_793_),
    .Y(_794_)
);

NAND3X1 _10601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_791_),
    .B(_794_),
    .C(_790_),
    .Y(_249_[16])
);

INVX1 _10602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [17]),
    .Y(_795_)
);

NAND2X1 _10603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_795_),
    .B(_597__bF$buf2),
    .Y(_796_)
);

INVX1 _10604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [17]),
    .Y(_797_)
);

NAND2X1 _10605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_797_),
    .B(_596__bF$buf1),
    .Y(_798_)
);

INVX1 _10606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [17]),
    .Y(_799_)
);

AOI21X1 _10607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_799_),
    .B(_595__bF$buf1),
    .C(_604__bF$buf2),
    .Y(_800_)
);

NAND3X1 _10608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_798_),
    .B(_800_),
    .C(_796_),
    .Y(_801_)
);

AOI22X1 _10609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [17]),
    .B(_611__bF$buf2),
    .C(_609__bF$buf2),
    .D(_0_[17]),
    .Y(_802_)
);

INVX1 _10610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [17]),
    .Y(_803_)
);

NOR2X1 _10611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_803_),
    .B(_614__bF$buf2),
    .Y(_804_)
);

AOI21X1 _10612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [17]),
    .B(_617__bF$buf2),
    .C(_804_),
    .Y(_805_)
);

NAND3X1 _10613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_802_),
    .B(_805_),
    .C(_801_),
    .Y(_249_[17])
);

INVX1 _10614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [18]),
    .Y(_806_)
);

NAND2X1 _10615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_806_),
    .B(_597__bF$buf1),
    .Y(_807_)
);

INVX1 _10616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [18]),
    .Y(_808_)
);

NAND2X1 _10617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_808_),
    .B(_596__bF$buf0),
    .Y(_809_)
);

INVX1 _10618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [18]),
    .Y(_810_)
);

AOI21X1 _10619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_810_),
    .B(_595__bF$buf0),
    .C(_604__bF$buf1),
    .Y(_811_)
);

NAND3X1 _10620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_809_),
    .B(_811_),
    .C(_807_),
    .Y(_812_)
);

AOI22X1 _10621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [18]),
    .B(_611__bF$buf1),
    .C(_609__bF$buf1),
    .D(_0_[18]),
    .Y(_813_)
);

INVX1 _10622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [18]),
    .Y(_814_)
);

NOR2X1 _10623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_814_),
    .B(_614__bF$buf1),
    .Y(_815_)
);

AOI21X1 _10624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [18]),
    .B(_617__bF$buf1),
    .C(_815_),
    .Y(_816_)
);

NAND3X1 _10625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_813_),
    .B(_816_),
    .C(_812_),
    .Y(_249_[18])
);

INVX1 _10626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [19]),
    .Y(_817_)
);

NAND2X1 _10627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_817_),
    .B(_597__bF$buf0),
    .Y(_818_)
);

INVX1 _10628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [19]),
    .Y(_819_)
);

NAND2X1 _10629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_819_),
    .B(_596__bF$buf4),
    .Y(_820_)
);

INVX1 _10630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [19]),
    .Y(_821_)
);

AOI21X1 _10631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_821_),
    .B(_595__bF$buf4),
    .C(_604__bF$buf0),
    .Y(_822_)
);

NAND3X1 _10632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_820_),
    .B(_822_),
    .C(_818_),
    .Y(_823_)
);

AOI22X1 _10633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [19]),
    .B(_611__bF$buf0),
    .C(_609__bF$buf0),
    .D(_0_[19]),
    .Y(_824_)
);

INVX1 _10634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [19]),
    .Y(_825_)
);

NOR2X1 _10635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_825_),
    .B(_614__bF$buf0),
    .Y(_826_)
);

AOI21X1 _10636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [19]),
    .B(_617__bF$buf0),
    .C(_826_),
    .Y(_827_)
);

NAND3X1 _10637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_824_),
    .B(_827_),
    .C(_823_),
    .Y(_249_[19])
);

INVX1 _10638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [20]),
    .Y(_828_)
);

NAND2X1 _10639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_828_),
    .B(_597__bF$buf4),
    .Y(_829_)
);

INVX1 _10640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [20]),
    .Y(_830_)
);

NAND2X1 _10641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_830_),
    .B(_596__bF$buf3),
    .Y(_831_)
);

INVX1 _10642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [20]),
    .Y(_832_)
);

AOI21X1 _10643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_832_),
    .B(_595__bF$buf3),
    .C(_604__bF$buf4),
    .Y(_833_)
);

NAND3X1 _10644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_831_),
    .B(_833_),
    .C(_829_),
    .Y(_834_)
);

AOI22X1 _10645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [20]),
    .B(_611__bF$buf4),
    .C(_617__bF$buf4),
    .D(\datapath.alu.c [20]),
    .Y(_835_)
);

INVX1 _10646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [20]),
    .Y(_836_)
);

NOR2X1 _10647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_836_),
    .B(_614__bF$buf4),
    .Y(_837_)
);

AOI21X1 _10648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[20]),
    .B(_609__bF$buf4),
    .C(_837_),
    .Y(_838_)
);

NAND3X1 _10649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_835_),
    .B(_838_),
    .C(_834_),
    .Y(_249_[20])
);

INVX1 _10650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [21]),
    .Y(_839_)
);

NAND2X1 _10651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_839_),
    .B(_597__bF$buf3),
    .Y(_840_)
);

INVX1 _10652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [21]),
    .Y(_841_)
);

NAND2X1 _10653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_841_),
    .B(_596__bF$buf2),
    .Y(_842_)
);

INVX1 _10654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [21]),
    .Y(_843_)
);

AOI21X1 _10655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_843_),
    .B(_595__bF$buf2),
    .C(_604__bF$buf3),
    .Y(_844_)
);

NAND3X1 _10656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_842_),
    .B(_844_),
    .C(_840_),
    .Y(_845_)
);

AOI22X1 _10657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [21]),
    .B(_611__bF$buf3),
    .C(_609__bF$buf3),
    .D(_0_[21]),
    .Y(_846_)
);

INVX1 _10658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [21]),
    .Y(_847_)
);

NOR2X1 _10659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_847_),
    .B(_614__bF$buf3),
    .Y(_848_)
);

AOI21X1 _10660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [21]),
    .B(_617__bF$buf3),
    .C(_848_),
    .Y(_849_)
);

NAND3X1 _10661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_846_),
    .B(_849_),
    .C(_845_),
    .Y(_249_[21])
);

INVX1 _10662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [22]),
    .Y(_850_)
);

NAND2X1 _10663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_850_),
    .B(_597__bF$buf2),
    .Y(_851_)
);

INVX1 _10664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [22]),
    .Y(_852_)
);

NAND2X1 _10665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_852_),
    .B(_596__bF$buf1),
    .Y(_853_)
);

INVX1 _10666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [22]),
    .Y(_854_)
);

AOI21X1 _10667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_854_),
    .B(_595__bF$buf1),
    .C(_604__bF$buf2),
    .Y(_855_)
);

NAND3X1 _10668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853_),
    .B(_855_),
    .C(_851_),
    .Y(_856_)
);

AOI22X1 _10669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [22]),
    .B(_611__bF$buf2),
    .C(_609__bF$buf2),
    .D(_0_[22]),
    .Y(_857_)
);

INVX1 _10670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [22]),
    .Y(_858_)
);

NOR2X1 _10671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_858_),
    .B(_614__bF$buf2),
    .Y(_859_)
);

AOI21X1 _10672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [22]),
    .B(_617__bF$buf2),
    .C(_859_),
    .Y(_860_)
);

NAND3X1 _10673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_857_),
    .B(_860_),
    .C(_856_),
    .Y(_249_[22])
);

INVX1 _10674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [23]),
    .Y(_861_)
);

NAND2X1 _10675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_861_),
    .B(_597__bF$buf1),
    .Y(_862_)
);

INVX1 _10676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [23]),
    .Y(_863_)
);

NAND2X1 _10677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_863_),
    .B(_596__bF$buf0),
    .Y(_864_)
);

INVX1 _10678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [23]),
    .Y(_865_)
);

AOI21X1 _10679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_865_),
    .B(_595__bF$buf0),
    .C(_604__bF$buf1),
    .Y(_866_)
);

NAND3X1 _10680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_864_),
    .B(_866_),
    .C(_862_),
    .Y(_867_)
);

AOI22X1 _10681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [23]),
    .B(_611__bF$buf1),
    .C(_617__bF$buf1),
    .D(\datapath.alu.c [23]),
    .Y(_868_)
);

INVX1 _10682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [23]),
    .Y(_869_)
);

NOR2X1 _10683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869_),
    .B(_614__bF$buf1),
    .Y(_870_)
);

AOI21X1 _10684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[23]),
    .B(_609__bF$buf1),
    .C(_870_),
    .Y(_871_)
);

NAND3X1 _10685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_868_),
    .B(_871_),
    .C(_867_),
    .Y(_249_[23])
);

INVX1 _10686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [24]),
    .Y(_872_)
);

NAND2X1 _10687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_872_),
    .B(_597__bF$buf0),
    .Y(_873_)
);

INVX1 _10688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [24]),
    .Y(_874_)
);

NAND2X1 _10689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_874_),
    .B(_596__bF$buf4),
    .Y(_875_)
);

INVX1 _10690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [24]),
    .Y(_876_)
);

AOI21X1 _10691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_876_),
    .B(_595__bF$buf4),
    .C(_604__bF$buf0),
    .Y(_877_)
);

NAND3X1 _10692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_875_),
    .B(_877_),
    .C(_873_),
    .Y(_878_)
);

AOI22X1 _10693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [24]),
    .B(_611__bF$buf0),
    .C(_609__bF$buf0),
    .D(_0_[24]),
    .Y(_879_)
);

INVX1 _10694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [24]),
    .Y(_880_)
);

NOR2X1 _10695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_880_),
    .B(_614__bF$buf0),
    .Y(_881_)
);

AOI21X1 _10696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [24]),
    .B(_617__bF$buf0),
    .C(_881_),
    .Y(_882_)
);

NAND3X1 _10697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_879_),
    .B(_882_),
    .C(_878_),
    .Y(_249_[24])
);

INVX1 _10698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [25]),
    .Y(_883_)
);

NAND2X1 _10699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_883_),
    .B(_597__bF$buf4),
    .Y(_884_)
);

INVX1 _10700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [25]),
    .Y(_885_)
);

NAND2X1 _10701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_885_),
    .B(_596__bF$buf3),
    .Y(_886_)
);

INVX1 _10702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [25]),
    .Y(_887_)
);

AOI21X1 _10703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887_),
    .B(_595__bF$buf3),
    .C(_604__bF$buf4),
    .Y(_888_)
);

NAND3X1 _10704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_),
    .B(_888_),
    .C(_884_),
    .Y(_889_)
);

AOI22X1 _10705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [25]),
    .B(_611__bF$buf4),
    .C(_617__bF$buf4),
    .D(\datapath.alu.c [25]),
    .Y(_890_)
);

INVX1 _10706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [25]),
    .Y(_891_)
);

NOR2X1 _10707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_891_),
    .B(_614__bF$buf4),
    .Y(_892_)
);

AOI21X1 _10708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[25]),
    .B(_609__bF$buf4),
    .C(_892_),
    .Y(_893_)
);

NAND3X1 _10709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_890_),
    .B(_893_),
    .C(_889_),
    .Y(_249_[25])
);

INVX1 _10710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [26]),
    .Y(_894_)
);

NAND2X1 _10711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_894_),
    .B(_597__bF$buf3),
    .Y(_895_)
);

INVX1 _10712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [26]),
    .Y(_896_)
);

NAND2X1 _10713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_896_),
    .B(_596__bF$buf2),
    .Y(_897_)
);

INVX1 _10714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [26]),
    .Y(_898_)
);

AOI21X1 _10715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_898_),
    .B(_595__bF$buf2),
    .C(_604__bF$buf3),
    .Y(_899_)
);

NAND3X1 _10716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_897_),
    .B(_899_),
    .C(_895_),
    .Y(_900_)
);

AOI22X1 _10717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [26]),
    .B(_611__bF$buf3),
    .C(_609__bF$buf3),
    .D(_0_[26]),
    .Y(_901_)
);

INVX1 _10718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [26]),
    .Y(_902_)
);

NOR2X1 _10719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_902_),
    .B(_614__bF$buf3),
    .Y(_903_)
);

AOI21X1 _10720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [26]),
    .B(_617__bF$buf3),
    .C(_903_),
    .Y(_904_)
);

NAND3X1 _10721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_901_),
    .B(_904_),
    .C(_900_),
    .Y(_249_[26])
);

INVX1 _10722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [27]),
    .Y(_905_)
);

NAND2X1 _10723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_905_),
    .B(_597__bF$buf2),
    .Y(_906_)
);

INVX1 _10724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [27]),
    .Y(_907_)
);

NAND2X1 _10725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_907_),
    .B(_596__bF$buf1),
    .Y(_908_)
);

INVX1 _10726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [27]),
    .Y(_909_)
);

AOI21X1 _10727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_909_),
    .B(_595__bF$buf1),
    .C(_604__bF$buf2),
    .Y(_910_)
);

NAND3X1 _10728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_908_),
    .B(_910_),
    .C(_906_),
    .Y(_911_)
);

AOI22X1 _10729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [27]),
    .B(_611__bF$buf2),
    .C(_617__bF$buf2),
    .D(\datapath.alu.c [27]),
    .Y(_912_)
);

INVX1 _10730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [27]),
    .Y(_913_)
);

NOR2X1 _10731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_913_),
    .B(_614__bF$buf2),
    .Y(_914_)
);

AOI21X1 _10732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[27]),
    .B(_609__bF$buf2),
    .C(_914_),
    .Y(_915_)
);

NAND3X1 _10733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_912_),
    .B(_915_),
    .C(_911_),
    .Y(_249_[27])
);

INVX1 _10734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [28]),
    .Y(_916_)
);

NAND2X1 _10735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_916_),
    .B(_597__bF$buf1),
    .Y(_917_)
);

INVX1 _10736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [28]),
    .Y(_918_)
);

NAND2X1 _10737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918_),
    .B(_596__bF$buf0),
    .Y(_919_)
);

INVX1 _10738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [28]),
    .Y(_920_)
);

AOI21X1 _10739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_920_),
    .B(_595__bF$buf0),
    .C(_604__bF$buf1),
    .Y(_921_)
);

NAND3X1 _10740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_919_),
    .B(_921_),
    .C(_917_),
    .Y(_922_)
);

AOI22X1 _10741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [28]),
    .B(_611__bF$buf1),
    .C(_609__bF$buf1),
    .D(_0_[28]),
    .Y(_923_)
);

INVX1 _10742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [28]),
    .Y(_924_)
);

NOR2X1 _10743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_924_),
    .B(_614__bF$buf1),
    .Y(_925_)
);

AOI21X1 _10744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [28]),
    .B(_617__bF$buf1),
    .C(_925_),
    .Y(_926_)
);

NAND3X1 _10745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_923_),
    .B(_926_),
    .C(_922_),
    .Y(_249_[28])
);

INVX1 _10746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [29]),
    .Y(_927_)
);

NAND2X1 _10747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_927_),
    .B(_597__bF$buf0),
    .Y(_928_)
);

INVX1 _10748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [29]),
    .Y(_929_)
);

NAND2X1 _10749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_929_),
    .B(_596__bF$buf4),
    .Y(_930_)
);

INVX1 _10750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [29]),
    .Y(_931_)
);

AOI21X1 _10751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_931_),
    .B(_595__bF$buf4),
    .C(_604__bF$buf0),
    .Y(_932_)
);

NAND3X1 _10752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_930_),
    .B(_932_),
    .C(_928_),
    .Y(_933_)
);

AOI22X1 _10753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [29]),
    .B(_611__bF$buf0),
    .C(_609__bF$buf0),
    .D(_0_[29]),
    .Y(_934_)
);

INVX1 _10754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [29]),
    .Y(_935_)
);

NOR2X1 _10755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_935_),
    .B(_614__bF$buf0),
    .Y(_936_)
);

AOI21X1 _10756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [29]),
    .B(_617__bF$buf0),
    .C(_936_),
    .Y(_937_)
);

NAND3X1 _10757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_934_),
    .B(_937_),
    .C(_933_),
    .Y(_249_[29])
);

INVX1 _10758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [30]),
    .Y(_938_)
);

NAND2X1 _10759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_938_),
    .B(_597__bF$buf4),
    .Y(_939_)
);

INVX1 _10760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.imm [30]),
    .Y(_940_)
);

NAND2X1 _10761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_940_),
    .B(_596__bF$buf3),
    .Y(_941_)
);

INVX1 _10762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [30]),
    .Y(_942_)
);

AOI21X1 _10763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_942_),
    .B(_595__bF$buf3),
    .C(_604__bF$buf4),
    .Y(_943_)
);

NAND3X1 _10764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_941_),
    .B(_943_),
    .C(_939_),
    .Y(_944_)
);

AOI22X1 _10765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [30]),
    .B(_611__bF$buf4),
    .C(_609__bF$buf4),
    .D(_0_[30]),
    .Y(_945_)
);

INVX1 _10766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [30]),
    .Y(_946_)
);

NOR2X1 _10767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_946_),
    .B(_614__bF$buf4),
    .Y(_947_)
);

AOI21X1 _10768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [30]),
    .B(_617__bF$buf4),
    .C(_947_),
    .Y(_948_)
);

NAND3X1 _10769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_945_),
    .B(_948_),
    .C(_944_),
    .Y(_249_[30])
);

INVX1 _10770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_data [31]),
    .Y(_949_)
);

NAND2X1 _10771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bsel[1]),
    .B(_594_),
    .Y(_950_)
);

NAND2X1 _10772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.immediatedecoder._12_ ),
    .B(_596__bF$buf2),
    .Y(_951_)
);

OAI21X1 _10773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_949_),
    .B(_950_),
    .C(_951_),
    .Y(_952_)
);

MUX2X1 _10774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.regb_data [31]),
    .B(_952_),
    .S(_597__bF$buf3),
    .Y(_953_)
);

NAND2X1 _10775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[31]),
    .B(_609__bF$buf3),
    .Y(_954_)
);

NAND2X1 _10776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [31]),
    .B(_611__bF$buf3),
    .Y(_955_)
);

NAND2X1 _10777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_955_),
    .B(_954_),
    .Y(_956_)
);

INVX1 _10778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [31]),
    .Y(_957_)
);

NAND2X1 _10779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [31]),
    .B(_617__bF$buf3),
    .Y(_958_)
);

OAI21X1 _10780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_957_),
    .B(_614__bF$buf3),
    .C(_958_),
    .Y(_959_)
);

NOR2X1 _10781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_956_),
    .B(_959_),
    .Y(_960_)
);

OAI21X1 _10782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_604__bF$buf3),
    .B(_953_),
    .C(_960_),
    .Y(_249_[31])
);

INVX1 _10783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [0]),
    .Y(_961_)
);

INVX1 _10784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(asel[0]),
    .Y(_962_)
);

AND2X2 _10785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_962_),
    .B(asel[1]),
    .Y(_963_)
);

NOR2X1 _10786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(asel[1]),
    .B(_962_),
    .Y(_964_)
);

NOR2X1 _10787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_964__bF$buf4),
    .B(_963__bF$buf4),
    .Y(_965_)
);

NAND2X1 _10788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_961_),
    .B(_965__bF$buf4),
    .Y(_966_)
);

NAND2X1 _10789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_601_),
    .B(_963__bF$buf3),
    .Y(_967_)
);

INVX1 _10790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(abpsel[2]),
    .Y(_968_)
);

NOR2X1 _10791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(abpsel[0]),
    .B(abpsel[1]),
    .Y(_969_)
);

NAND2X1 _10792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_968_),
    .B(_969_),
    .Y(_970_)
);

AOI21X1 _10793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_358_),
    .B(_964__bF$buf3),
    .C(_970__bF$buf4),
    .Y(_971_)
);

NAND3X1 _10794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_967_),
    .B(_971_),
    .C(_966_),
    .Y(_972_)
);

INVX1 _10795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_969_),
    .Y(_973_)
);

NOR2X1 _10796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_968_),
    .B(_973_),
    .Y(_974_)
);

INVX1 _10797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(abpsel[1]),
    .Y(_975_)
);

NOR2X1 _10798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(abpsel[2]),
    .B(_975_),
    .Y(_976_)
);

AND2X2 _10799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_976_),
    .B(abpsel[0]),
    .Y(_977_)
);

AOI22X1 _10800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [0]),
    .B(_974__bF$buf4),
    .C(_977__bF$buf4),
    .D(_0__0_bF$buf2),
    .Y(_978_)
);

OAI21X1 _10801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(abpsel[2]),
    .B(_975_),
    .C(_973_),
    .Y(_979_)
);

NOR2X1 _10802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_613_),
    .B(_979__bF$buf4),
    .Y(_980_)
);

INVX1 _10803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_976_),
    .Y(_981_)
);

NOR2X1 _10804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(abpsel[0]),
    .B(_981_),
    .Y(_982_)
);

AOI21X1 _10805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.condtrue ),
    .B(_982__bF$buf4),
    .C(_980_),
    .Y(_983_)
);

NAND3X1 _10806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_978_),
    .B(_983_),
    .C(_972_),
    .Y(_248_[0])
);

INVX1 _10807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [1]),
    .Y(_984_)
);

NAND2X1 _10808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_984_),
    .B(_965__bF$buf3),
    .Y(_985_)
);

NAND2X1 _10809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_623_),
    .B(_963__bF$buf2),
    .Y(_986_)
);

AOI21X1 _10810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_360_),
    .B(_964__bF$buf2),
    .C(_970__bF$buf3),
    .Y(_987_)
);

NAND3X1 _10811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_986_),
    .B(_987_),
    .C(_985_),
    .Y(_988_)
);

AOI22X1 _10812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [1]),
    .B(_974__bF$buf3),
    .C(_982__bF$buf3),
    .D(\datapath.alu.c [1]),
    .Y(_989_)
);

NOR2X1 _10813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_627_),
    .B(_979__bF$buf3),
    .Y(_990_)
);

AOI21X1 _10814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf7),
    .B(_977__bF$buf3),
    .C(_990_),
    .Y(_991_)
);

NAND3X1 _10815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_989_),
    .B(_991_),
    .C(_988_),
    .Y(_248_[1])
);

INVX1 _10816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [2]),
    .Y(_992_)
);

NAND2X1 _10817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_992_),
    .B(_965__bF$buf2),
    .Y(_993_)
);

NAND2X1 _10818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_634_),
    .B(_963__bF$buf1),
    .Y(_994_)
);

AOI21X1 _10819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_362_),
    .B(_964__bF$buf1),
    .C(_970__bF$buf2),
    .Y(_995_)
);

NAND3X1 _10820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_994_),
    .B(_995_),
    .C(_993_),
    .Y(_996_)
);

AOI22X1 _10821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [2]),
    .B(_974__bF$buf2),
    .C(_977__bF$buf2),
    .D(_0_[2]),
    .Y(_997_)
);

NOR2X1 _10822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_638_),
    .B(_979__bF$buf2),
    .Y(_998_)
);

AOI21X1 _10823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [2]),
    .B(_982__bF$buf2),
    .C(_998_),
    .Y(_999_)
);

NAND3X1 _10824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_997_),
    .B(_999_),
    .C(_996_),
    .Y(_248_[2])
);

INVX1 _10825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [3]),
    .Y(_1000_)
);

NAND2X1 _10826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1000_),
    .B(_965__bF$buf1),
    .Y(_1001_)
);

NAND2X1 _10827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_645_),
    .B(_963__bF$buf0),
    .Y(_1002_)
);

AOI21X1 _10828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_364_),
    .B(_964__bF$buf0),
    .C(_970__bF$buf1),
    .Y(_1003_)
);

NAND3X1 _10829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002_),
    .B(_1003_),
    .C(_1001_),
    .Y(_1004_)
);

AOI22X1 _10830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [3]),
    .B(_974__bF$buf1),
    .C(_982__bF$buf1),
    .D(\datapath.alu.c [3]),
    .Y(_1005_)
);

NOR2X1 _10831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_649_),
    .B(_979__bF$buf1),
    .Y(_1006_)
);

AOI21X1 _10832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[3]),
    .B(_977__bF$buf1),
    .C(_1006_),
    .Y(_1007_)
);

NAND3X1 _10833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1005_),
    .B(_1007_),
    .C(_1004_),
    .Y(_248_[3])
);

INVX1 _10834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [4]),
    .Y(_1008_)
);

NAND2X1 _10835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1008_),
    .B(_965__bF$buf0),
    .Y(_1009_)
);

NAND2X1 _10836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_656_),
    .B(_963__bF$buf4),
    .Y(_1010_)
);

AOI21X1 _10837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_366_),
    .B(_964__bF$buf4),
    .C(_970__bF$buf0),
    .Y(_1011_)
);

NAND3X1 _10838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010_),
    .B(_1011_),
    .C(_1009_),
    .Y(_1012_)
);

AOI22X1 _10839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [4]),
    .B(_974__bF$buf0),
    .C(_982__bF$buf0),
    .D(\datapath.alu.c [4]),
    .Y(_1013_)
);

NOR2X1 _10840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_660_),
    .B(_979__bF$buf0),
    .Y(_1014_)
);

AOI21X1 _10841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[4]),
    .B(_977__bF$buf0),
    .C(_1014_),
    .Y(_1015_)
);

NAND3X1 _10842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1013_),
    .B(_1015_),
    .C(_1012_),
    .Y(_248_[4])
);

INVX1 _10843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [5]),
    .Y(_1016_)
);

NAND2X1 _10844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1016_),
    .B(_965__bF$buf4),
    .Y(_1017_)
);

NAND2X1 _10845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_667_),
    .B(_963__bF$buf3),
    .Y(_1018_)
);

AOI21X1 _10846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_368_),
    .B(_964__bF$buf3),
    .C(_970__bF$buf4),
    .Y(_1019_)
);

NAND3X1 _10847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1018_),
    .B(_1019_),
    .C(_1017_),
    .Y(_1020_)
);

AOI22X1 _10848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [5]),
    .B(_974__bF$buf4),
    .C(_982__bF$buf4),
    .D(\datapath.alu.c [5]),
    .Y(_1021_)
);

NOR2X1 _10849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_671_),
    .B(_979__bF$buf4),
    .Y(_1022_)
);

AOI21X1 _10850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[5]),
    .B(_977__bF$buf4),
    .C(_1022_),
    .Y(_1023_)
);

NAND3X1 _10851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1021_),
    .B(_1023_),
    .C(_1020_),
    .Y(_248_[5])
);

INVX1 _10852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [6]),
    .Y(_1024_)
);

NAND2X1 _10853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1024_),
    .B(_965__bF$buf3),
    .Y(_1025_)
);

NAND2X1 _10854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_678_),
    .B(_963__bF$buf2),
    .Y(_1026_)
);

AOI21X1 _10855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_370_),
    .B(_964__bF$buf2),
    .C(_970__bF$buf3),
    .Y(_1027_)
);

NAND3X1 _10856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1026_),
    .B(_1027_),
    .C(_1025_),
    .Y(_1028_)
);

AOI22X1 _10857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [6]),
    .B(_974__bF$buf3),
    .C(_977__bF$buf3),
    .D(_0_[6]),
    .Y(_1029_)
);

NOR2X1 _10858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_682_),
    .B(_979__bF$buf3),
    .Y(_1030_)
);

AOI21X1 _10859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [6]),
    .B(_982__bF$buf3),
    .C(_1030_),
    .Y(_1031_)
);

NAND3X1 _10860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1029_),
    .B(_1031_),
    .C(_1028_),
    .Y(_248_[6])
);

INVX1 _10861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [7]),
    .Y(_1032_)
);

NAND2X1 _10862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1032_),
    .B(_965__bF$buf2),
    .Y(_1033_)
);

NAND2X1 _10863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_689_),
    .B(_963__bF$buf1),
    .Y(_1034_)
);

AOI21X1 _10864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_372_),
    .B(_964__bF$buf1),
    .C(_970__bF$buf2),
    .Y(_1035_)
);

NAND3X1 _10865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1034_),
    .B(_1035_),
    .C(_1033_),
    .Y(_1036_)
);

AOI22X1 _10866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [7]),
    .B(_974__bF$buf2),
    .C(_982__bF$buf2),
    .D(\datapath.alu.c [7]),
    .Y(_1037_)
);

NOR2X1 _10867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_693_),
    .B(_979__bF$buf2),
    .Y(_1038_)
);

AOI21X1 _10868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[7]),
    .B(_977__bF$buf2),
    .C(_1038_),
    .Y(_1039_)
);

NAND3X1 _10869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1037_),
    .B(_1039_),
    .C(_1036_),
    .Y(_248_[7])
);

INVX1 _10870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [8]),
    .Y(_1040_)
);

NAND2X1 _10871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1040_),
    .B(_965__bF$buf1),
    .Y(_1041_)
);

NAND2X1 _10872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_700_),
    .B(_963__bF$buf0),
    .Y(_1042_)
);

AOI21X1 _10873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_374_),
    .B(_964__bF$buf0),
    .C(_970__bF$buf1),
    .Y(_1043_)
);

NAND3X1 _10874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1042_),
    .B(_1043_),
    .C(_1041_),
    .Y(_1044_)
);

AOI22X1 _10875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [8]),
    .B(_974__bF$buf1),
    .C(_982__bF$buf1),
    .D(\datapath.alu.c [8]),
    .Y(_1045_)
);

NOR2X1 _10876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_704_),
    .B(_979__bF$buf1),
    .Y(_1046_)
);

AOI21X1 _10877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[8]),
    .B(_977__bF$buf1),
    .C(_1046_),
    .Y(_1047_)
);

NAND3X1 _10878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1045_),
    .B(_1047_),
    .C(_1044_),
    .Y(_248_[8])
);

INVX1 _10879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [9]),
    .Y(_1048_)
);

NAND2X1 _10880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1048_),
    .B(_965__bF$buf0),
    .Y(_1049_)
);

NAND2X1 _10881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_711_),
    .B(_963__bF$buf4),
    .Y(_1050_)
);

AOI21X1 _10882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_376_),
    .B(_964__bF$buf4),
    .C(_970__bF$buf0),
    .Y(_1051_)
);

NAND3X1 _10883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1050_),
    .B(_1051_),
    .C(_1049_),
    .Y(_1052_)
);

AOI22X1 _10884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [9]),
    .B(_974__bF$buf0),
    .C(_977__bF$buf0),
    .D(_0_[9]),
    .Y(_1053_)
);

NOR2X1 _10885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_715_),
    .B(_979__bF$buf0),
    .Y(_1054_)
);

AOI21X1 _10886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [9]),
    .B(_982__bF$buf0),
    .C(_1054_),
    .Y(_1055_)
);

NAND3X1 _10887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1053_),
    .B(_1055_),
    .C(_1052_),
    .Y(_248_[9])
);

INVX1 _10888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [10]),
    .Y(_1056_)
);

NAND2X1 _10889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1056_),
    .B(_965__bF$buf4),
    .Y(_1057_)
);

NAND2X1 _10890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_722_),
    .B(_963__bF$buf3),
    .Y(_1058_)
);

AOI21X1 _10891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_378_),
    .B(_964__bF$buf3),
    .C(_970__bF$buf4),
    .Y(_1059_)
);

NAND3X1 _10892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1058_),
    .B(_1059_),
    .C(_1057_),
    .Y(_1060_)
);

AOI22X1 _10893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [10]),
    .B(_974__bF$buf4),
    .C(_982__bF$buf4),
    .D(\datapath.alu.c [10]),
    .Y(_1061_)
);

NOR2X1 _10894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_726_),
    .B(_979__bF$buf4),
    .Y(_1062_)
);

AOI21X1 _10895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[10]),
    .B(_977__bF$buf4),
    .C(_1062_),
    .Y(_1063_)
);

NAND3X1 _10896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1061_),
    .B(_1063_),
    .C(_1060_),
    .Y(_248_[10])
);

INVX1 _10897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [11]),
    .Y(_1064_)
);

NAND2X1 _10898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1064_),
    .B(_965__bF$buf3),
    .Y(_1065_)
);

NAND2X1 _10899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_733_),
    .B(_963__bF$buf2),
    .Y(_1066_)
);

AOI21X1 _10900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_380_),
    .B(_964__bF$buf2),
    .C(_970__bF$buf3),
    .Y(_1067_)
);

NAND3X1 _10901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1066_),
    .B(_1067_),
    .C(_1065_),
    .Y(_1068_)
);

AOI22X1 _10902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [11]),
    .B(_974__bF$buf3),
    .C(_977__bF$buf3),
    .D(_0_[11]),
    .Y(_1069_)
);

NOR2X1 _10903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_737_),
    .B(_979__bF$buf3),
    .Y(_1070_)
);

AOI21X1 _10904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [11]),
    .B(_982__bF$buf3),
    .C(_1070_),
    .Y(_1071_)
);

NAND3X1 _10905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1069_),
    .B(_1071_),
    .C(_1068_),
    .Y(_248_[11])
);

INVX1 _10906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [12]),
    .Y(_1072_)
);

NAND2X1 _10907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1072_),
    .B(_965__bF$buf2),
    .Y(_1073_)
);

NAND2X1 _10908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_744_),
    .B(_963__bF$buf1),
    .Y(_1074_)
);

AOI21X1 _10909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_382_),
    .B(_964__bF$buf1),
    .C(_970__bF$buf2),
    .Y(_1075_)
);

NAND3X1 _10910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1074_),
    .B(_1075_),
    .C(_1073_),
    .Y(_1076_)
);

AOI22X1 _10911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [12]),
    .B(_974__bF$buf2),
    .C(_977__bF$buf2),
    .D(_0_[12]),
    .Y(_1077_)
);

NOR2X1 _10912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_748_),
    .B(_979__bF$buf2),
    .Y(_1078_)
);

AOI21X1 _10913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [12]),
    .B(_982__bF$buf2),
    .C(_1078_),
    .Y(_1079_)
);

NAND3X1 _10914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1077_),
    .B(_1079_),
    .C(_1076_),
    .Y(_248_[12])
);

INVX1 _10915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [13]),
    .Y(_1080_)
);

NAND2X1 _10916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1080_),
    .B(_965__bF$buf1),
    .Y(_1081_)
);

NAND2X1 _10917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_),
    .B(_963__bF$buf0),
    .Y(_1082_)
);

AOI21X1 _10918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_384_),
    .B(_964__bF$buf0),
    .C(_970__bF$buf1),
    .Y(_1083_)
);

NAND3X1 _10919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1082_),
    .B(_1083_),
    .C(_1081_),
    .Y(_1084_)
);

AOI22X1 _10920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [13]),
    .B(_974__bF$buf1),
    .C(_977__bF$buf1),
    .D(_0_[13]),
    .Y(_1085_)
);

NOR2X1 _10921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_759_),
    .B(_979__bF$buf1),
    .Y(_1086_)
);

AOI21X1 _10922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [13]),
    .B(_982__bF$buf1),
    .C(_1086_),
    .Y(_1087_)
);

NAND3X1 _10923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1085_),
    .B(_1087_),
    .C(_1084_),
    .Y(_248_[13])
);

INVX1 _10924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [14]),
    .Y(_1088_)
);

NAND2X1 _10925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1088_),
    .B(_965__bF$buf0),
    .Y(_1089_)
);

NAND2X1 _10926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_766_),
    .B(_963__bF$buf4),
    .Y(_1090_)
);

AOI21X1 _10927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_386_),
    .B(_964__bF$buf4),
    .C(_970__bF$buf0),
    .Y(_1091_)
);

NAND3X1 _10928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1090_),
    .B(_1091_),
    .C(_1089_),
    .Y(_1092_)
);

AOI22X1 _10929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [14]),
    .B(_974__bF$buf0),
    .C(_977__bF$buf0),
    .D(_0_[14]),
    .Y(_1093_)
);

NOR2X1 _10930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_770_),
    .B(_979__bF$buf0),
    .Y(_1094_)
);

AOI21X1 _10931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [14]),
    .B(_982__bF$buf0),
    .C(_1094_),
    .Y(_1095_)
);

NAND3X1 _10932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1093_),
    .B(_1095_),
    .C(_1092_),
    .Y(_248_[14])
);

INVX1 _10933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [15]),
    .Y(_1096_)
);

NAND2X1 _10934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1096_),
    .B(_965__bF$buf4),
    .Y(_1097_)
);

NAND2X1 _10935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_777_),
    .B(_963__bF$buf3),
    .Y(_1098_)
);

AOI21X1 _10936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_388_),
    .B(_964__bF$buf3),
    .C(_970__bF$buf4),
    .Y(_1099_)
);

NAND3X1 _10937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1098_),
    .B(_1099_),
    .C(_1097_),
    .Y(_1100_)
);

AOI22X1 _10938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [15]),
    .B(_974__bF$buf4),
    .C(_977__bF$buf4),
    .D(_0_[15]),
    .Y(_1101_)
);

NOR2X1 _10939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_781_),
    .B(_979__bF$buf4),
    .Y(_1102_)
);

AOI21X1 _10940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [15]),
    .B(_982__bF$buf4),
    .C(_1102_),
    .Y(_1103_)
);

NAND3X1 _10941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1101_),
    .B(_1103_),
    .C(_1100_),
    .Y(_248_[15])
);

INVX1 _10942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [16]),
    .Y(_1104_)
);

NAND2X1 _10943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1104_),
    .B(_965__bF$buf3),
    .Y(_1105_)
);

NAND2X1 _10944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_788_),
    .B(_963__bF$buf2),
    .Y(_1106_)
);

AOI21X1 _10945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_390_),
    .B(_964__bF$buf2),
    .C(_970__bF$buf3),
    .Y(_1107_)
);

NAND3X1 _10946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1106_),
    .B(_1107_),
    .C(_1105_),
    .Y(_1108_)
);

AOI22X1 _10947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [16]),
    .B(_974__bF$buf3),
    .C(_982__bF$buf3),
    .D(\datapath.alu.c [16]),
    .Y(_1109_)
);

NOR2X1 _10948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_792_),
    .B(_979__bF$buf3),
    .Y(_1110_)
);

AOI21X1 _10949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[16]),
    .B(_977__bF$buf3),
    .C(_1110_),
    .Y(_1111_)
);

NAND3X1 _10950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1109_),
    .B(_1111_),
    .C(_1108_),
    .Y(_248_[16])
);

INVX1 _10951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [17]),
    .Y(_1112_)
);

NAND2X1 _10952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1112_),
    .B(_965__bF$buf2),
    .Y(_1113_)
);

NAND2X1 _10953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_799_),
    .B(_963__bF$buf1),
    .Y(_1114_)
);

AOI21X1 _10954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_392_),
    .B(_964__bF$buf1),
    .C(_970__bF$buf2),
    .Y(_1115_)
);

NAND3X1 _10955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1114_),
    .B(_1115_),
    .C(_1113_),
    .Y(_1116_)
);

AOI22X1 _10956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [17]),
    .B(_974__bF$buf2),
    .C(_982__bF$buf2),
    .D(\datapath.alu.c [17]),
    .Y(_1117_)
);

NOR2X1 _10957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_803_),
    .B(_979__bF$buf2),
    .Y(_1118_)
);

AOI21X1 _10958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[17]),
    .B(_977__bF$buf2),
    .C(_1118_),
    .Y(_1119_)
);

NAND3X1 _10959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1117_),
    .B(_1119_),
    .C(_1116_),
    .Y(_248_[17])
);

INVX1 _10960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [18]),
    .Y(_1120_)
);

NAND2X1 _10961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1120_),
    .B(_965__bF$buf1),
    .Y(_1121_)
);

NAND2X1 _10962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_810_),
    .B(_963__bF$buf0),
    .Y(_1122_)
);

AOI21X1 _10963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_394_),
    .B(_964__bF$buf0),
    .C(_970__bF$buf1),
    .Y(_1123_)
);

NAND3X1 _10964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1122_),
    .B(_1123_),
    .C(_1121_),
    .Y(_1124_)
);

AOI22X1 _10965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [18]),
    .B(_974__bF$buf1),
    .C(_982__bF$buf1),
    .D(\datapath.alu.c [18]),
    .Y(_1125_)
);

NOR2X1 _10966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_814_),
    .B(_979__bF$buf1),
    .Y(_1126_)
);

AOI21X1 _10967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[18]),
    .B(_977__bF$buf1),
    .C(_1126_),
    .Y(_1127_)
);

NAND3X1 _10968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1125_),
    .B(_1127_),
    .C(_1124_),
    .Y(_248_[18])
);

INVX1 _10969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [19]),
    .Y(_1128_)
);

NAND2X1 _10970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1128_),
    .B(_965__bF$buf0),
    .Y(_1129_)
);

NAND2X1 _10971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_821_),
    .B(_963__bF$buf4),
    .Y(_1130_)
);

AOI21X1 _10972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_396_),
    .B(_964__bF$buf4),
    .C(_970__bF$buf0),
    .Y(_1131_)
);

NAND3X1 _10973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1130_),
    .B(_1131_),
    .C(_1129_),
    .Y(_1132_)
);

AOI22X1 _10974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [19]),
    .B(_974__bF$buf0),
    .C(_977__bF$buf0),
    .D(_0_[19]),
    .Y(_1133_)
);

NOR2X1 _10975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_825_),
    .B(_979__bF$buf0),
    .Y(_1134_)
);

AOI21X1 _10976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [19]),
    .B(_982__bF$buf0),
    .C(_1134_),
    .Y(_1135_)
);

NAND3X1 _10977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1133_),
    .B(_1135_),
    .C(_1132_),
    .Y(_248_[19])
);

INVX1 _10978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [20]),
    .Y(_1136_)
);

NAND2X1 _10979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1136_),
    .B(_965__bF$buf4),
    .Y(_1137_)
);

NAND2X1 _10980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_832_),
    .B(_963__bF$buf3),
    .Y(_1138_)
);

AOI21X1 _10981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_398_),
    .B(_964__bF$buf3),
    .C(_970__bF$buf4),
    .Y(_1139_)
);

NAND3X1 _10982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1138_),
    .B(_1139_),
    .C(_1137_),
    .Y(_1140_)
);

AOI22X1 _10983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [20]),
    .B(_974__bF$buf4),
    .C(_982__bF$buf4),
    .D(\datapath.alu.c [20]),
    .Y(_1141_)
);

NOR2X1 _10984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_836_),
    .B(_979__bF$buf4),
    .Y(_1142_)
);

AOI21X1 _10985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[20]),
    .B(_977__bF$buf4),
    .C(_1142_),
    .Y(_1143_)
);

NAND3X1 _10986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1141_),
    .B(_1143_),
    .C(_1140_),
    .Y(_248_[20])
);

INVX1 _10987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [21]),
    .Y(_1144_)
);

NAND2X1 _10988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1144_),
    .B(_965__bF$buf3),
    .Y(_1145_)
);

NAND2X1 _10989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_843_),
    .B(_963__bF$buf2),
    .Y(_1146_)
);

AOI21X1 _10990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_400_),
    .B(_964__bF$buf2),
    .C(_970__bF$buf3),
    .Y(_1147_)
);

NAND3X1 _10991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1146_),
    .B(_1147_),
    .C(_1145_),
    .Y(_1148_)
);

AOI22X1 _10992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [21]),
    .B(_974__bF$buf3),
    .C(_982__bF$buf3),
    .D(\datapath.alu.c [21]),
    .Y(_1149_)
);

NOR2X1 _10993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_847_),
    .B(_979__bF$buf3),
    .Y(_1150_)
);

AOI21X1 _10994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[21]),
    .B(_977__bF$buf3),
    .C(_1150_),
    .Y(_1151_)
);

NAND3X1 _10995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1149_),
    .B(_1151_),
    .C(_1148_),
    .Y(_248_[21])
);

INVX1 _10996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [22]),
    .Y(_1152_)
);

NAND2X1 _10997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1152_),
    .B(_965__bF$buf2),
    .Y(_1153_)
);

NAND2X1 _10998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_854_),
    .B(_963__bF$buf1),
    .Y(_1154_)
);

AOI21X1 _10999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_402_),
    .B(_964__bF$buf1),
    .C(_970__bF$buf2),
    .Y(_1155_)
);

NAND3X1 _11000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1154_),
    .B(_1155_),
    .C(_1153_),
    .Y(_1156_)
);

AOI22X1 _11001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [22]),
    .B(_974__bF$buf2),
    .C(_977__bF$buf2),
    .D(_0_[22]),
    .Y(_1157_)
);

NOR2X1 _11002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_858_),
    .B(_979__bF$buf2),
    .Y(_1158_)
);

AOI21X1 _11003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [22]),
    .B(_982__bF$buf2),
    .C(_1158_),
    .Y(_1159_)
);

NAND3X1 _11004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1157_),
    .B(_1159_),
    .C(_1156_),
    .Y(_248_[22])
);

INVX1 _11005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [23]),
    .Y(_1160_)
);

NAND2X1 _11006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1160_),
    .B(_965__bF$buf1),
    .Y(_1161_)
);

NAND2X1 _11007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_865_),
    .B(_963__bF$buf0),
    .Y(_1162_)
);

AOI21X1 _11008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_404_),
    .B(_964__bF$buf0),
    .C(_970__bF$buf1),
    .Y(_1163_)
);

NAND3X1 _11009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1162_),
    .B(_1163_),
    .C(_1161_),
    .Y(_1164_)
);

AOI22X1 _11010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [23]),
    .B(_974__bF$buf1),
    .C(_982__bF$buf1),
    .D(\datapath.alu.c [23]),
    .Y(_1165_)
);

NOR2X1 _11011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869_),
    .B(_979__bF$buf1),
    .Y(_1166_)
);

AOI21X1 _11012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[23]),
    .B(_977__bF$buf1),
    .C(_1166_),
    .Y(_1167_)
);

NAND3X1 _11013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1165_),
    .B(_1167_),
    .C(_1164_),
    .Y(_248_[23])
);

INVX1 _11014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [24]),
    .Y(_1168_)
);

NAND2X1 _11015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1168_),
    .B(_965__bF$buf0),
    .Y(_1169_)
);

NAND2X1 _11016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_876_),
    .B(_963__bF$buf4),
    .Y(_1170_)
);

AOI21X1 _11017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_406_),
    .B(_964__bF$buf4),
    .C(_970__bF$buf0),
    .Y(_1171_)
);

NAND3X1 _11018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1170_),
    .B(_1171_),
    .C(_1169_),
    .Y(_1172_)
);

AOI22X1 _11019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [24]),
    .B(_974__bF$buf0),
    .C(_982__bF$buf0),
    .D(\datapath.alu.c [24]),
    .Y(_1173_)
);

NOR2X1 _11020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_880_),
    .B(_979__bF$buf0),
    .Y(_1174_)
);

AOI21X1 _11021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[24]),
    .B(_977__bF$buf0),
    .C(_1174_),
    .Y(_1175_)
);

NAND3X1 _11022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1173_),
    .B(_1175_),
    .C(_1172_),
    .Y(_248_[24])
);

INVX1 _11023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [25]),
    .Y(_1176_)
);

NAND2X1 _11024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1176_),
    .B(_965__bF$buf4),
    .Y(_1177_)
);

NAND2X1 _11025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887_),
    .B(_963__bF$buf3),
    .Y(_1178_)
);

AOI21X1 _11026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_408_),
    .B(_964__bF$buf3),
    .C(_970__bF$buf4),
    .Y(_1179_)
);

NAND3X1 _11027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1178_),
    .B(_1179_),
    .C(_1177_),
    .Y(_1180_)
);

AOI22X1 _11028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [25]),
    .B(_974__bF$buf4),
    .C(_977__bF$buf4),
    .D(_0_[25]),
    .Y(_1181_)
);

NOR2X1 _11029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_891_),
    .B(_979__bF$buf4),
    .Y(_1182_)
);

AOI21X1 _11030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [25]),
    .B(_982__bF$buf4),
    .C(_1182_),
    .Y(_1183_)
);

NAND3X1 _11031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1181_),
    .B(_1183_),
    .C(_1180_),
    .Y(_248_[25])
);

INVX1 _11032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [26]),
    .Y(_1184_)
);

NAND2X1 _11033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1184_),
    .B(_965__bF$buf3),
    .Y(_1185_)
);

NAND2X1 _11034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_898_),
    .B(_963__bF$buf2),
    .Y(_1186_)
);

AOI21X1 _11035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_410_),
    .B(_964__bF$buf2),
    .C(_970__bF$buf3),
    .Y(_1187_)
);

NAND3X1 _11036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1186_),
    .B(_1187_),
    .C(_1185_),
    .Y(_1188_)
);

AOI22X1 _11037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [26]),
    .B(_974__bF$buf3),
    .C(_982__bF$buf3),
    .D(\datapath.alu.c [26]),
    .Y(_1189_)
);

NOR2X1 _11038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_902_),
    .B(_979__bF$buf3),
    .Y(_1190_)
);

AOI21X1 _11039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[26]),
    .B(_977__bF$buf3),
    .C(_1190_),
    .Y(_1191_)
);

NAND3X1 _11040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1189_),
    .B(_1191_),
    .C(_1188_),
    .Y(_248_[26])
);

INVX1 _11041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [27]),
    .Y(_1192_)
);

NAND2X1 _11042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1192_),
    .B(_965__bF$buf2),
    .Y(_1193_)
);

NAND2X1 _11043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_909_),
    .B(_963__bF$buf1),
    .Y(_1194_)
);

AOI21X1 _11044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_412_),
    .B(_964__bF$buf1),
    .C(_970__bF$buf2),
    .Y(_1195_)
);

NAND3X1 _11045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1194_),
    .B(_1195_),
    .C(_1193_),
    .Y(_1196_)
);

AOI22X1 _11046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [27]),
    .B(_974__bF$buf2),
    .C(_982__bF$buf2),
    .D(\datapath.alu.c [27]),
    .Y(_1197_)
);

NOR2X1 _11047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_913_),
    .B(_979__bF$buf2),
    .Y(_1198_)
);

AOI21X1 _11048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[27]),
    .B(_977__bF$buf2),
    .C(_1198_),
    .Y(_1199_)
);

NAND3X1 _11049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1197_),
    .B(_1199_),
    .C(_1196_),
    .Y(_248_[27])
);

INVX1 _11050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [28]),
    .Y(_1200_)
);

NAND2X1 _11051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1200_),
    .B(_965__bF$buf1),
    .Y(_1201_)
);

NAND2X1 _11052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_920_),
    .B(_963__bF$buf0),
    .Y(_1202_)
);

AOI21X1 _11053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_414_),
    .B(_964__bF$buf0),
    .C(_970__bF$buf1),
    .Y(_1203_)
);

NAND3X1 _11054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1202_),
    .B(_1203_),
    .C(_1201_),
    .Y(_1204_)
);

AOI22X1 _11055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [28]),
    .B(_974__bF$buf1),
    .C(_982__bF$buf1),
    .D(\datapath.alu.c [28]),
    .Y(_1205_)
);

NOR2X1 _11056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_924_),
    .B(_979__bF$buf1),
    .Y(_1206_)
);

AOI21X1 _11057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[28]),
    .B(_977__bF$buf1),
    .C(_1206_),
    .Y(_1207_)
);

NAND3X1 _11058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1205_),
    .B(_1207_),
    .C(_1204_),
    .Y(_248_[28])
);

INVX1 _11059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [29]),
    .Y(_1208_)
);

NAND2X1 _11060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1208_),
    .B(_965__bF$buf0),
    .Y(_1209_)
);

NAND2X1 _11061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_931_),
    .B(_963__bF$buf4),
    .Y(_1210_)
);

AOI21X1 _11062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_416_),
    .B(_964__bF$buf4),
    .C(_970__bF$buf0),
    .Y(_1211_)
);

NAND3X1 _11063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1210_),
    .B(_1211_),
    .C(_1209_),
    .Y(_1212_)
);

AOI22X1 _11064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [29]),
    .B(_974__bF$buf0),
    .C(_977__bF$buf0),
    .D(_0_[29]),
    .Y(_1213_)
);

NOR2X1 _11065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_935_),
    .B(_979__bF$buf0),
    .Y(_1214_)
);

AOI21X1 _11066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [29]),
    .B(_982__bF$buf0),
    .C(_1214_),
    .Y(_1215_)
);

NAND3X1 _11067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1213_),
    .B(_1215_),
    .C(_1212_),
    .Y(_248_[29])
);

NAND2X1 _11068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(asel[1]),
    .B(_962_),
    .Y(_1216_)
);

NAND2X1 _11069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [30]),
    .B(_964__bF$buf3),
    .Y(_1217_)
);

OAI21X1 _11070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_942_),
    .B(_1216_),
    .C(_1217_),
    .Y(_1218_)
);

MUX2X1 _11071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [30]),
    .B(_1218_),
    .S(_965__bF$buf4),
    .Y(_1219_)
);

NAND2X1 _11072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [30]),
    .B(_974__bF$buf4),
    .Y(_1220_)
);

NAND2X1 _11073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[30]),
    .B(_977__bF$buf4),
    .Y(_1221_)
);

NAND2X1 _11074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1220_),
    .B(_1221_),
    .Y(_1222_)
);

NAND2X1 _11075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [30]),
    .B(_982__bF$buf4),
    .Y(_1223_)
);

OAI21X1 _11076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_946_),
    .B(_979__bF$buf4),
    .C(_1223_),
    .Y(_1224_)
);

NOR2X1 _11077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1222_),
    .B(_1224_),
    .Y(_1225_)
);

OAI21X1 _11078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_970__bF$buf4),
    .B(_1219_),
    .C(_1225_),
    .Y(_248_[30])
);

NAND2X1 _11079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [31]),
    .B(_964__bF$buf2),
    .Y(_1226_)
);

OAI21X1 _11080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_949_),
    .B(_1216_),
    .C(_1226_),
    .Y(_1227_)
);

MUX2X1 _11081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.rega_data [31]),
    .B(_1227_),
    .S(_965__bF$buf3),
    .Y(_1228_)
);

NAND2X1 _11082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [31]),
    .B(_982__bF$buf3),
    .Y(_1229_)
);

NAND2X1 _11083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memdataload [31]),
    .B(_974__bF$buf3),
    .Y(_1230_)
);

NAND2X1 _11084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1230_),
    .B(_1229_),
    .Y(_1231_)
);

NAND2X1 _11085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[31]),
    .B(_977__bF$buf3),
    .Y(_1232_)
);

OAI21X1 _11086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_957_),
    .B(_979__bF$buf3),
    .C(_1232_),
    .Y(_1233_)
);

NOR2X1 _11087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1233_),
    .B(_1231_),
    .Y(_1234_)
);

OAI21X1 _11088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_970__bF$buf3),
    .B(_1228_),
    .C(_1234_),
    .Y(_248_[31])
);

INVX1 _11089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.wb_sel [1]),
    .Y(_1235_)
);

NOR2X1 _11090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.wb_sel [0]),
    .B(_1235_),
    .Y(_1236_)
);

INVX1 _11091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.wb_sel [0]),
    .Y(_1237_)
);

NOR2X1 _11092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1237_),
    .B(_1235_),
    .Y(_1238_)
);

AOI22X1 _11093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236__bF$buf4),
    .B(\datapath.wbpc_4 [0]),
    .C(\datapath.regcsrwb [0]),
    .D(_1238__bF$buf4),
    .Y(_1239_)
);

NOR2X1 _11094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.wb_sel [0]),
    .B(\controlunit.wb_sel [1]),
    .Y(_1240_)
);

NAND2X1 _11095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [0]),
    .B(_1240__bF$buf4),
    .Y(_1241_)
);

NOR2X1 _11096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.wb_sel [1]),
    .B(_1237_),
    .Y(_1242_)
);

NAND2X1 _11097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [0]),
    .B(_1242__bF$buf4),
    .Y(_1243_)
);

NAND3X1 _11098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1241_),
    .B(_1243_),
    .C(_1239_),
    .Y(\datapath.rd [0])
);

AOI22X1 _11099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [1]),
    .B(_1240__bF$buf3),
    .C(_1236__bF$buf3),
    .D(\datapath.wbpc_4 [1]),
    .Y(_1244_)
);

NAND2X1 _11100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [1]),
    .B(_1242__bF$buf3),
    .Y(_1245_)
);

NAND2X1 _11101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrwb [1]),
    .B(_1238__bF$buf3),
    .Y(_1246_)
);

NAND3X1 _11102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1245_),
    .B(_1246_),
    .C(_1244_),
    .Y(\datapath.rd [1])
);

NAND2X1 _11103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [2]),
    .B(_1242__bF$buf2),
    .Y(_1247_)
);

NAND2X1 _11104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrwb [2]),
    .B(_1238__bF$buf2),
    .Y(_1248_)
);

AOI22X1 _11105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [2]),
    .B(_1240__bF$buf2),
    .C(_1236__bF$buf2),
    .D(\datapath.wbpc_4 [2]),
    .Y(_1249_)
);

NAND3X1 _11106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1247_),
    .B(_1248_),
    .C(_1249_),
    .Y(\datapath.rd [2])
);

AOI22X1 _11107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236__bF$buf1),
    .B(\datapath.wbpc_4 [3]),
    .C(\datapath.regcsrwb [3]),
    .D(_1238__bF$buf1),
    .Y(_1250_)
);

NAND2X1 _11108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [3]),
    .B(_1240__bF$buf1),
    .Y(_1251_)
);

NAND2X1 _11109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [3]),
    .B(_1242__bF$buf1),
    .Y(_1252_)
);

NAND3X1 _11110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1251_),
    .B(_1252_),
    .C(_1250_),
    .Y(\datapath.rd [3])
);

AOI22X1 _11111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [4]),
    .B(_1240__bF$buf0),
    .C(_1236__bF$buf0),
    .D(\datapath.wbpc_4 [4]),
    .Y(_1253_)
);

NAND2X1 _11112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [4]),
    .B(_1242__bF$buf0),
    .Y(_1254_)
);

NAND2X1 _11113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrwb [4]),
    .B(_1238__bF$buf0),
    .Y(_1255_)
);

NAND3X1 _11114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1254_),
    .B(_1255_),
    .C(_1253_),
    .Y(\datapath.rd [4])
);

AOI22X1 _11115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236__bF$buf4),
    .B(\datapath.wbpc_4 [5]),
    .C(\datapath.regcsrwb [5]),
    .D(_1238__bF$buf4),
    .Y(_1256_)
);

NAND2X1 _11116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [5]),
    .B(_1240__bF$buf4),
    .Y(_1257_)
);

NAND2X1 _11117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [5]),
    .B(_1242__bF$buf4),
    .Y(_1258_)
);

NAND3X1 _11118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1257_),
    .B(_1258_),
    .C(_1256_),
    .Y(\datapath.rd [5])
);

NAND2X1 _11119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [6]),
    .B(_1242__bF$buf3),
    .Y(_1259_)
);

NAND2X1 _11120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrwb [6]),
    .B(_1238__bF$buf3),
    .Y(_1260_)
);

AOI22X1 _11121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [6]),
    .B(_1240__bF$buf3),
    .C(_1236__bF$buf3),
    .D(\datapath.wbpc_4 [6]),
    .Y(_1261_)
);

NAND3X1 _11122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1259_),
    .B(_1260_),
    .C(_1261_),
    .Y(\datapath.rd [6])
);

AOI22X1 _11123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236__bF$buf2),
    .B(\datapath.wbpc_4 [7]),
    .C(\datapath.regcsrwb [7]),
    .D(_1238__bF$buf2),
    .Y(_1262_)
);

NAND2X1 _11124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [7]),
    .B(_1240__bF$buf2),
    .Y(_1263_)
);

NAND2X1 _11125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [7]),
    .B(_1242__bF$buf2),
    .Y(_1264_)
);

NAND3X1 _11126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1263_),
    .B(_1264_),
    .C(_1262_),
    .Y(\datapath.rd [7])
);

AOI22X1 _11127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236__bF$buf1),
    .B(\datapath.wbpc_4 [8]),
    .C(\datapath.regcsrwb [8]),
    .D(_1238__bF$buf1),
    .Y(_1265_)
);

NAND2X1 _11128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [8]),
    .B(_1240__bF$buf1),
    .Y(_1266_)
);

NAND2X1 _11129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [8]),
    .B(_1242__bF$buf1),
    .Y(_1267_)
);

NAND3X1 _11130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1266_),
    .B(_1267_),
    .C(_1265_),
    .Y(\datapath.rd [8])
);

AOI22X1 _11131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [9]),
    .B(_1240__bF$buf0),
    .C(_1236__bF$buf0),
    .D(\datapath.wbpc_4 [9]),
    .Y(_1268_)
);

NAND2X1 _11132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [9]),
    .B(_1242__bF$buf0),
    .Y(_1269_)
);

NAND2X1 _11133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrwb [9]),
    .B(_1238__bF$buf0),
    .Y(_1270_)
);

NAND3X1 _11134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1269_),
    .B(_1270_),
    .C(_1268_),
    .Y(\datapath.rd [9])
);

NAND2X1 _11135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [10]),
    .B(_1242__bF$buf4),
    .Y(_1271_)
);

NAND2X1 _11136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrwb [10]),
    .B(_1238__bF$buf4),
    .Y(_1272_)
);

AOI22X1 _11137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [10]),
    .B(_1240__bF$buf4),
    .C(_1236__bF$buf4),
    .D(\datapath.wbpc_4 [10]),
    .Y(_1273_)
);

NAND3X1 _11138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1271_),
    .B(_1272_),
    .C(_1273_),
    .Y(\datapath.rd [10])
);

AOI22X1 _11139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236__bF$buf3),
    .B(\datapath.wbpc_4 [11]),
    .C(\datapath.regcsrwb [11]),
    .D(_1238__bF$buf3),
    .Y(_1274_)
);

NAND2X1 _11140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [11]),
    .B(_1240__bF$buf3),
    .Y(_1275_)
);

NAND2X1 _11141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [11]),
    .B(_1242__bF$buf3),
    .Y(_1276_)
);

NAND3X1 _11142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1275_),
    .B(_1276_),
    .C(_1274_),
    .Y(\datapath.rd [11])
);

AOI22X1 _11143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [12]),
    .B(_1240__bF$buf2),
    .C(_1236__bF$buf2),
    .D(\datapath.wbpc_4 [12]),
    .Y(_1277_)
);

NAND2X1 _11144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [12]),
    .B(_1242__bF$buf2),
    .Y(_1278_)
);

NAND2X1 _11145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrwb [12]),
    .B(_1238__bF$buf2),
    .Y(_1279_)
);

NAND3X1 _11146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1278_),
    .B(_1279_),
    .C(_1277_),
    .Y(\datapath.rd [12])
);

AOI22X1 _11147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236__bF$buf1),
    .B(\datapath.wbpc_4 [13]),
    .C(\datapath.regcsrwb [13]),
    .D(_1238__bF$buf1),
    .Y(_1280_)
);

NAND2X1 _11148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [13]),
    .B(_1240__bF$buf1),
    .Y(_1281_)
);

NAND2X1 _11149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [13]),
    .B(_1242__bF$buf1),
    .Y(_1282_)
);

NAND3X1 _11150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1281_),
    .B(_1282_),
    .C(_1280_),
    .Y(\datapath.rd [13])
);

NAND2X1 _11151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [14]),
    .B(_1242__bF$buf0),
    .Y(_1283_)
);

NAND2X1 _11152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrwb [14]),
    .B(_1238__bF$buf0),
    .Y(_1284_)
);

AOI22X1 _11153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [14]),
    .B(_1240__bF$buf0),
    .C(_1236__bF$buf0),
    .D(\datapath.wbpc_4 [14]),
    .Y(_1285_)
);

NAND3X1 _11154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1283_),
    .B(_1284_),
    .C(_1285_),
    .Y(\datapath.rd [14])
);

AOI22X1 _11155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236__bF$buf4),
    .B(\datapath.wbpc_4 [15]),
    .C(\datapath.regcsrwb [15]),
    .D(_1238__bF$buf4),
    .Y(_1286_)
);

NAND2X1 _11156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [15]),
    .B(_1240__bF$buf4),
    .Y(_1287_)
);

NAND2X1 _11157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [15]),
    .B(_1242__bF$buf4),
    .Y(_1288_)
);

NAND3X1 _11158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1287_),
    .B(_1288_),
    .C(_1286_),
    .Y(\datapath.rd [15])
);

AOI22X1 _11159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236__bF$buf3),
    .B(\datapath.wbpc_4 [16]),
    .C(\datapath.regcsrwb [16]),
    .D(_1238__bF$buf3),
    .Y(_1289_)
);

NAND2X1 _11160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [16]),
    .B(_1240__bF$buf3),
    .Y(_1290_)
);

NAND2X1 _11161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [16]),
    .B(_1242__bF$buf3),
    .Y(_1291_)
);

NAND3X1 _11162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1290_),
    .B(_1291_),
    .C(_1289_),
    .Y(\datapath.rd [16])
);

AOI22X1 _11163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [17]),
    .B(_1240__bF$buf2),
    .C(_1236__bF$buf2),
    .D(\datapath.wbpc_4 [17]),
    .Y(_1292_)
);

NAND2X1 _11164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [17]),
    .B(_1242__bF$buf2),
    .Y(_1293_)
);

NAND2X1 _11165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrwb [17]),
    .B(_1238__bF$buf2),
    .Y(_1294_)
);

NAND3X1 _11166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1293_),
    .B(_1294_),
    .C(_1292_),
    .Y(\datapath.rd [17])
);

NAND2X1 _11167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [18]),
    .B(_1242__bF$buf1),
    .Y(_1295_)
);

NAND2X1 _11168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrwb [18]),
    .B(_1238__bF$buf1),
    .Y(_1296_)
);

AOI22X1 _11169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [18]),
    .B(_1240__bF$buf1),
    .C(_1236__bF$buf1),
    .D(\datapath.wbpc_4 [18]),
    .Y(_1297_)
);

NAND3X1 _11170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1295_),
    .B(_1296_),
    .C(_1297_),
    .Y(\datapath.rd [18])
);

AOI22X1 _11171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236__bF$buf0),
    .B(\datapath.wbpc_4 [19]),
    .C(\datapath.regcsrwb [19]),
    .D(_1238__bF$buf0),
    .Y(_1298_)
);

NAND2X1 _11172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [19]),
    .B(_1240__bF$buf0),
    .Y(_1299_)
);

NAND2X1 _11173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [19]),
    .B(_1242__bF$buf0),
    .Y(_1300_)
);

NAND3X1 _11174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1299_),
    .B(_1300_),
    .C(_1298_),
    .Y(\datapath.rd [19])
);

AOI22X1 _11175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [20]),
    .B(_1240__bF$buf4),
    .C(_1236__bF$buf4),
    .D(\datapath.wbpc_4 [20]),
    .Y(_1301_)
);

NAND2X1 _11176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [20]),
    .B(_1242__bF$buf4),
    .Y(_1302_)
);

NAND2X1 _11177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrwb [20]),
    .B(_1238__bF$buf4),
    .Y(_1303_)
);

NAND3X1 _11178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1302_),
    .B(_1303_),
    .C(_1301_),
    .Y(\datapath.rd [20])
);

AOI22X1 _11179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236__bF$buf3),
    .B(\datapath.wbpc_4 [21]),
    .C(\datapath.regcsrwb [21]),
    .D(_1238__bF$buf3),
    .Y(_1304_)
);

NAND2X1 _11180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [21]),
    .B(_1240__bF$buf3),
    .Y(_1305_)
);

NAND2X1 _11181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [21]),
    .B(_1242__bF$buf3),
    .Y(_1306_)
);

NAND3X1 _11182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1305_),
    .B(_1306_),
    .C(_1304_),
    .Y(\datapath.rd [21])
);

NAND2X1 _11183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [22]),
    .B(_1242__bF$buf2),
    .Y(_1307_)
);

NAND2X1 _11184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrwb [22]),
    .B(_1238__bF$buf2),
    .Y(_1308_)
);

AOI22X1 _11185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [22]),
    .B(_1240__bF$buf2),
    .C(_1236__bF$buf2),
    .D(\datapath.wbpc_4 [22]),
    .Y(_1309_)
);

NAND3X1 _11186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1307_),
    .B(_1308_),
    .C(_1309_),
    .Y(\datapath.rd [22])
);

AOI22X1 _11187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236__bF$buf1),
    .B(\datapath.wbpc_4 [23]),
    .C(\datapath.regcsrwb [23]),
    .D(_1238__bF$buf1),
    .Y(_1310_)
);

NAND2X1 _11188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [23]),
    .B(_1240__bF$buf1),
    .Y(_1311_)
);

NAND2X1 _11189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [23]),
    .B(_1242__bF$buf1),
    .Y(_1312_)
);

NAND3X1 _11190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1311_),
    .B(_1312_),
    .C(_1310_),
    .Y(\datapath.rd [23])
);

AOI22X1 _11191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236__bF$buf0),
    .B(\datapath.wbpc_4 [24]),
    .C(\datapath.regcsrwb [24]),
    .D(_1238__bF$buf0),
    .Y(_1313_)
);

NAND2X1 _11192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [24]),
    .B(_1240__bF$buf0),
    .Y(_1314_)
);

NAND2X1 _11193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [24]),
    .B(_1242__bF$buf0),
    .Y(_1315_)
);

NAND3X1 _11194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1314_),
    .B(_1315_),
    .C(_1313_),
    .Y(\datapath.rd [24])
);

AOI22X1 _11195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [25]),
    .B(_1240__bF$buf4),
    .C(_1236__bF$buf4),
    .D(\datapath.wbpc_4 [25]),
    .Y(_1316_)
);

NAND2X1 _11196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [25]),
    .B(_1242__bF$buf4),
    .Y(_1317_)
);

NAND2X1 _11197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrwb [25]),
    .B(_1238__bF$buf4),
    .Y(_1318_)
);

NAND3X1 _11198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1317_),
    .B(_1318_),
    .C(_1316_),
    .Y(\datapath.rd [25])
);

NAND2X1 _11199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [26]),
    .B(_1242__bF$buf3),
    .Y(_1319_)
);

NAND2X1 _11200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrwb [26]),
    .B(_1238__bF$buf3),
    .Y(_1320_)
);

AOI22X1 _11201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [26]),
    .B(_1240__bF$buf3),
    .C(_1236__bF$buf3),
    .D(\datapath.wbpc_4 [26]),
    .Y(_1321_)
);

NAND3X1 _11202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1319_),
    .B(_1320_),
    .C(_1321_),
    .Y(\datapath.rd [26])
);

AOI22X1 _11203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236__bF$buf2),
    .B(\datapath.wbpc_4 [27]),
    .C(\datapath.regcsrwb [27]),
    .D(_1238__bF$buf2),
    .Y(_1322_)
);

NAND2X1 _11204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [27]),
    .B(_1240__bF$buf2),
    .Y(_1323_)
);

NAND2X1 _11205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [27]),
    .B(_1242__bF$buf2),
    .Y(_1324_)
);

NAND3X1 _11206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1323_),
    .B(_1324_),
    .C(_1322_),
    .Y(\datapath.rd [27])
);

AOI22X1 _11207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [28]),
    .B(_1240__bF$buf1),
    .C(_1236__bF$buf1),
    .D(\datapath.wbpc_4 [28]),
    .Y(_1325_)
);

NAND2X1 _11208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [28]),
    .B(_1242__bF$buf1),
    .Y(_1326_)
);

NAND2X1 _11209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrwb [28]),
    .B(_1238__bF$buf1),
    .Y(_1327_)
);

NAND3X1 _11210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1326_),
    .B(_1327_),
    .C(_1325_),
    .Y(\datapath.rd [28])
);

AOI22X1 _11211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236__bF$buf0),
    .B(\datapath.wbpc_4 [29]),
    .C(\datapath.regcsrwb [29]),
    .D(_1238__bF$buf0),
    .Y(_1328_)
);

NAND2X1 _11212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [29]),
    .B(_1240__bF$buf0),
    .Y(_1329_)
);

NAND2X1 _11213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [29]),
    .B(_1242__bF$buf0),
    .Y(_1330_)
);

NAND3X1 _11214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1329_),
    .B(_1330_),
    .C(_1328_),
    .Y(\datapath.rd [29])
);

NAND2X1 _11215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [30]),
    .B(_1242__bF$buf4),
    .Y(_1331_)
);

NAND2X1 _11216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrwb [30]),
    .B(_1238__bF$buf4),
    .Y(_1332_)
);

AOI22X1 _11217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [30]),
    .B(_1240__bF$buf4),
    .C(_1236__bF$buf4),
    .D(\datapath.wbpc_4 [30]),
    .Y(_1333_)
);

NAND3X1 _11218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1331_),
    .B(_1332_),
    .C(_1333_),
    .Y(\datapath.rd [30])
);

AOI22X1 _11219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236__bF$buf3),
    .B(\datapath.wbpc_4 [31]),
    .C(\datapath.regcsrwb [31]),
    .D(_1238__bF$buf3),
    .Y(_1334_)
);

NAND2X1 _11220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcwb [31]),
    .B(_1240__bF$buf3),
    .Y(_1335_)
);

NAND2X1 _11221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regloadwb [31]),
    .B(_1242__bF$buf3),
    .Y(_1336_)
);

NAND3X1 _11222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1335_),
    .B(_1336_),
    .C(_1334_),
    .Y(\datapath.rd [31])
);

MUX2X1 _11223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcondt ),
    .B(\datapath.regz ),
    .S(\datapath.meminstr [14]),
    .Y(_1337_)
);

XNOR2X1 _11224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1337_),
    .B(\datapath.meminstr [12]),
    .Y(\datapath.tkbranch )
);

NOR2X1 _11225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regwbtrap ),
    .B(\datapath.regmret_bF$buf4 ),
    .Y(_1338_)
);

NOR2X1 _11226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regpcsel [0]),
    .B(branch),
    .Y(_1339_)
);

NAND2X1 _11227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1338_),
    .B(_1339_),
    .Y(\datapath._60_ )
);

INVX1 _11228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regpcsel [1]),
    .Y(_1340_)
);

NAND2X1 _11229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1340_),
    .B(_1338_),
    .Y(\datapath._62_ )
);

OAI21X1 _11230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.rs2_bypass_sel [0]),
    .B(\bypassandflushunit.rs2_bypass_sel [1]),
    .C(\bypassandflushunit.rs2_bypass_sel [2]),
    .Y(_251_)
);

OAI21X1 _11231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bbpsel[0]),
    .B(bbpsel[1]),
    .C(bbpsel[2]),
    .Y(_252_)
);

OAI21X1 _11232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(abpsel[0]),
    .B(abpsel[1]),
    .C(abpsel[2]),
    .Y(_253_)
);

NOR2X1 _11233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf1),
    .B(\datapath._62_ ),
    .Y(_1341_)
);

AND2X2 _11234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1339_),
    .B(_1341_),
    .Y(\datapath.pcstall )
);

INVX1 _11235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.csrfile_wen ),
    .Y(_1342_)
);

NOR2X1 _11236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [18]),
    .B(_261_),
    .Y(_1343_)
);

NOR2X1 _11237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [19]),
    .B(\datapath.meminstr [17]),
    .Y(_1344_)
);

NOR2X1 _11238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [16]),
    .B(\datapath.meminstr [15]),
    .Y(_1345_)
);

AND2X2 _11239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1344_),
    .B(_1345_),
    .Y(_1346_)
);

AOI21X1 _11240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1343_),
    .B(_1346_),
    .C(_1342_),
    .Y(\datapath.allowcsrwrite )
);

AND2X2 _11241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [0]),
    .B(\datapath.regimmalu [0]),
    .Y(_1347_)
);

OR2X2 _11242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [1]),
    .B(\datapath.regimmalu [1]),
    .Y(_1348_)
);

NAND2X1 _11243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [1]),
    .B(\datapath.regimmalu [1]),
    .Y(_1349_)
);

NAND2X1 _11244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1349_),
    .B(_1348_),
    .Y(_1350_)
);

XNOR2X1 _11245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1350_),
    .B(_1347_),
    .Y(\datapath.jumptarget [1])
);

NAND2X1 _11246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [0]),
    .B(\datapath.regimmalu [0]),
    .Y(_1351_)
);

NOR2X1 _11247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [1]),
    .B(\datapath.regimmalu [1]),
    .Y(_1352_)
);

OAI21X1 _11248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1352_),
    .B(_1351_),
    .C(_1349_),
    .Y(_1353_)
);

XNOR2X1 _11249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [2]),
    .B(\datapath.regimmalu [2]),
    .Y(_1354_)
);

XNOR2X1 _11250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1353_),
    .B(_1354_),
    .Y(\datapath.jumptarget [2])
);

AND2X2 _11251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [1]),
    .B(\datapath.regimmalu [1]),
    .Y(_1355_)
);

AOI21X1 _11252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1347_),
    .B(_1348_),
    .C(_1355_),
    .Y(_1356_)
);

NAND2X1 _11253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [2]),
    .B(\datapath.regimmalu [2]),
    .Y(_1357_)
);

OAI21X1 _11254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1356_),
    .B(_1354_),
    .C(_1357_),
    .Y(_1358_)
);

XNOR2X1 _11255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [3]),
    .B(\datapath.regimmalu [3]),
    .Y(_1359_)
);

XNOR2X1 _11256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1358_),
    .B(_1359_),
    .Y(\datapath.jumptarget [3])
);

INVX1 _11257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1354_),
    .Y(_1360_)
);

INVX1 _11258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1359_),
    .Y(_1361_)
);

NAND3X1 _11259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1353_),
    .B(_1360_),
    .C(_1361_),
    .Y(_1362_)
);

INVX1 _11260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [3]),
    .Y(_1363_)
);

INVX1 _11261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regimmalu [3]),
    .Y(_1364_)
);

NOR2X1 _11262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1363_),
    .B(_1364_),
    .Y(_1365_)
);

AOI21X1 _11263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1363_),
    .B(_1364_),
    .C(_1357_),
    .Y(_1366_)
);

NOR2X1 _11264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1365_),
    .B(_1366_),
    .Y(_1367_)
);

NAND2X1 _11265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1367_),
    .B(_1362_),
    .Y(_1368_)
);

XNOR2X1 _11266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [4]),
    .B(\datapath.regimmalu [4]),
    .Y(_1369_)
);

XNOR2X1 _11267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1368_),
    .B(_1369_),
    .Y(\datapath.jumptarget [4])
);

INVX1 _11268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1368_),
    .Y(_1370_)
);

NAND2X1 _11269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [4]),
    .B(\datapath.regimmalu [4]),
    .Y(_1371_)
);

OAI21X1 _11270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1370_),
    .B(_1369_),
    .C(_1371_),
    .Y(_1372_)
);

XNOR2X1 _11271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [5]),
    .B(\datapath.regimmalu [5]),
    .Y(_1373_)
);

XNOR2X1 _11272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1372_),
    .B(_1373_),
    .Y(\datapath.jumptarget [5])
);

NAND2X1 _11273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [5]),
    .B(\datapath.regimmalu [5]),
    .Y(_1374_)
);

INVX1 _11274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1371_),
    .Y(_1375_)
);

OAI21X1 _11275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [5]),
    .B(\datapath.regimmalu [5]),
    .C(_1375_),
    .Y(_1376_)
);

AND2X2 _11276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1376_),
    .B(_1374_),
    .Y(_1377_)
);

XOR2X1 _11277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [4]),
    .B(\datapath.regimmalu [4]),
    .Y(_1378_)
);

XOR2X1 _11278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [5]),
    .B(\datapath.regimmalu [5]),
    .Y(_1379_)
);

NAND2X1 _11279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1378_),
    .B(_1379_),
    .Y(_1380_)
);

OAI21X1 _11280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1370_),
    .B(_1380_),
    .C(_1377_),
    .Y(_1381_)
);

XNOR2X1 _11281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [6]),
    .B(\datapath.regimmalu [6]),
    .Y(_1382_)
);

XNOR2X1 _11282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1381_),
    .B(_1382_),
    .Y(\datapath.jumptarget [6])
);

NAND2X1 _11283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [6]),
    .B(\datapath.regimmalu [6]),
    .Y(_1383_)
);

INVX1 _11284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1383_),
    .Y(_1384_)
);

XOR2X1 _11285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [6]),
    .B(\datapath.regimmalu [6]),
    .Y(_1385_)
);

AOI21X1 _11286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1385_),
    .B(_1381_),
    .C(_1384_),
    .Y(_1386_)
);

XOR2X1 _11287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [7]),
    .B(\datapath.regimmalu [7]),
    .Y(_1387_)
);

XNOR2X1 _11288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1386_),
    .B(_1387_),
    .Y(\datapath.jumptarget [7])
);

NOR2X1 _11289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1369_),
    .B(_1373_),
    .Y(_1388_)
);

XNOR2X1 _11290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [7]),
    .B(\datapath.regimmalu [7]),
    .Y(_1389_)
);

NOR2X1 _11291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1382_),
    .B(_1389_),
    .Y(_1390_)
);

NAND2X1 _11292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1388_),
    .B(_1390_),
    .Y(_1391_)
);

AOI21X1 _11293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1367_),
    .B(_1362_),
    .C(_1391_),
    .Y(_1392_)
);

NAND2X1 _11294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1385_),
    .B(_1387_),
    .Y(_1393_)
);

NAND2X1 _11295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [7]),
    .B(\datapath.regimmalu [7]),
    .Y(_1394_)
);

OAI21X1 _11296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1389_),
    .B(_1383_),
    .C(_1394_),
    .Y(_1395_)
);

INVX1 _11297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1395_),
    .Y(_1396_)
);

OAI21X1 _11298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1377_),
    .B(_1393_),
    .C(_1396_),
    .Y(_1397_)
);

NOR2X1 _11299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1397_),
    .B(_1392_),
    .Y(_1398_)
);

XOR2X1 _11300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [8]),
    .B(\datapath.regimmalu [8]),
    .Y(_1399_)
);

XNOR2X1 _11301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1398_),
    .B(_1399_),
    .Y(\datapath.jumptarget [8])
);

INVX1 _11302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [8]),
    .Y(_1400_)
);

INVX1 _11303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regimmalu [8]),
    .Y(_1401_)
);

NOR2X1 _11304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1400_),
    .B(_1401_),
    .Y(_1402_)
);

INVX1 _11305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1402_),
    .Y(_1403_)
);

INVX1 _11306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1399_),
    .Y(_1404_)
);

OAI21X1 _11307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1398_),
    .B(_1404_),
    .C(_1403_),
    .Y(_1405_)
);

XOR2X1 _11308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [9]),
    .B(\datapath.regimmalu [9]),
    .Y(_1406_)
);

INVX1 _11309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1406_),
    .Y(_1407_)
);

XNOR2X1 _11310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1405_),
    .B(_1407_),
    .Y(\datapath.jumptarget [9])
);

INVX1 _11311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [9]),
    .Y(_1408_)
);

INVX1 _11312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regimmalu [9]),
    .Y(_1409_)
);

NAND2X1 _11313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1408_),
    .B(_1409_),
    .Y(_1410_)
);

NOR2X1 _11314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1408_),
    .B(_1409_),
    .Y(_1411_)
);

AOI21X1 _11315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1410_),
    .B(_1402_),
    .C(_1411_),
    .Y(_1412_)
);

NAND2X1 _11316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1399_),
    .B(_1406_),
    .Y(_1413_)
);

OAI21X1 _11317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1398_),
    .B(_1413_),
    .C(_1412_),
    .Y(_1414_)
);

XOR2X1 _11318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [10]),
    .B(\datapath.regimmalu [10]),
    .Y(_1415_)
);

XOR2X1 _11319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1414_),
    .B(_1415_),
    .Y(\datapath.jumptarget [10])
);

AND2X2 _11320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [10]),
    .B(\datapath.regimmalu [10]),
    .Y(_1416_)
);

AOI21X1 _11321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1415_),
    .B(_1414_),
    .C(_1416_),
    .Y(_1417_)
);

XOR2X1 _11322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [11]),
    .B(\datapath.regimmalu [11]),
    .Y(_1418_)
);

XNOR2X1 _11323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1417_),
    .B(_1418_),
    .Y(\datapath.jumptarget [11])
);

NAND2X1 _11324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1415_),
    .B(_1418_),
    .Y(_1419_)
);

AND2X2 _11325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [11]),
    .B(\datapath.regimmalu [11]),
    .Y(_1420_)
);

AOI21X1 _11326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1416_),
    .B(_1418_),
    .C(_1420_),
    .Y(_1421_)
);

OAI21X1 _11327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1419_),
    .B(_1412_),
    .C(_1421_),
    .Y(_1422_)
);

NOR2X1 _11328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1413_),
    .B(_1419_),
    .Y(_1423_)
);

INVX1 _11329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1423_),
    .Y(_1424_)
);

NOR2X1 _11330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1424_),
    .B(_1398_),
    .Y(_1425_)
);

NOR2X1 _11331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1422_),
    .B(_1425_),
    .Y(_1426_)
);

NOR2X1 _11332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [12]),
    .B(\datapath.regimmalu [12]),
    .Y(_1427_)
);

AND2X2 _11333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [12]),
    .B(\datapath.regimmalu [12]),
    .Y(_1428_)
);

NOR2X1 _11334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1427_),
    .B(_1428_),
    .Y(_1429_)
);

XNOR2X1 _11335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1426_),
    .B(_1429_),
    .Y(\datapath.jumptarget [12])
);

NAND2X1 _11336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [12]),
    .B(\datapath.regimmalu [12]),
    .Y(_1430_)
);

OAI21X1 _11337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1426_),
    .B(_1427_),
    .C(_1430_),
    .Y(_1431_)
);

XOR2X1 _11338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [13]),
    .B(\datapath.regimmalu [13]),
    .Y(_1432_)
);

XOR2X1 _11339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1431_),
    .B(_1432_),
    .Y(\datapath.jumptarget [13])
);

NAND2X1 _11340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [13]),
    .B(\datapath.regimmalu [13]),
    .Y(_1433_)
);

NAND2X1 _11341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1430_),
    .B(_1433_),
    .Y(_1434_)
);

OAI21X1 _11342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [13]),
    .B(\datapath.regimmalu [13]),
    .C(_1434_),
    .Y(_1435_)
);

NAND2X1 _11343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1432_),
    .B(_1429_),
    .Y(_1436_)
);

OAI21X1 _11344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1426_),
    .B(_1436_),
    .C(_1435_),
    .Y(_1437_)
);

XOR2X1 _11345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [14]),
    .B(\datapath.regimmalu [14]),
    .Y(_1438_)
);

XOR2X1 _11346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1437_),
    .B(_1438_),
    .Y(\datapath.jumptarget [14])
);

NAND2X1 _11347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [14]),
    .B(\datapath.regimmalu [14]),
    .Y(_1439_)
);

INVX1 _11348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1439_),
    .Y(_1440_)
);

AOI21X1 _11349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1438_),
    .B(_1437_),
    .C(_1440_),
    .Y(_1441_)
);

NOR2X1 _11350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [15]),
    .B(\datapath.regimmalu [15]),
    .Y(_1442_)
);

AND2X2 _11351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [15]),
    .B(\datapath.regimmalu [15]),
    .Y(_1443_)
);

NOR2X1 _11352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1442_),
    .B(_1443_),
    .Y(_1444_)
);

XNOR2X1 _11353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1441_),
    .B(_1444_),
    .Y(\datapath.jumptarget [15])
);

NAND2X1 _11354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1438_),
    .B(_1444_),
    .Y(_1445_)
);

NOR2X1 _11355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1436_),
    .B(_1445_),
    .Y(_1446_)
);

NAND2X1 _11356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1423_),
    .B(_1446_),
    .Y(_1447_)
);

AOI21X1 _11357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1440_),
    .B(_1444_),
    .C(_1443_),
    .Y(_1448_)
);

OAI21X1 _11358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1435_),
    .B(_1445_),
    .C(_1448_),
    .Y(_1449_)
);

AOI21X1 _11359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1422_),
    .B(_1446_),
    .C(_1449_),
    .Y(_1450_)
);

OAI21X1 _11360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1398_),
    .B(_1447_),
    .C(_1450_),
    .Y(_1451_)
);

INVX1 _11361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [16]),
    .Y(_1452_)
);

INVX1 _11362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regimmalu [16]),
    .Y(_1453_)
);

NAND2X1 _11363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1452_),
    .B(_1453_),
    .Y(_1454_)
);

NAND2X1 _11364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [16]),
    .B(\datapath.regimmalu [16]),
    .Y(_1455_)
);

AND2X2 _11365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1454_),
    .B(_1455_),
    .Y(_1456_)
);

INVX1 _11366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1456_),
    .Y(_1457_)
);

XNOR2X1 _11367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1451_),
    .B(_1457_),
    .Y(\datapath.jumptarget [16])
);

INVX1 _11368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1455_),
    .Y(_1458_)
);

AOI21X1 _11369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1454_),
    .B(_1451_),
    .C(_1458_),
    .Y(_1459_)
);

INVX1 _11370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [17]),
    .Y(_1460_)
);

INVX1 _11371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regimmalu [17]),
    .Y(_1461_)
);

NOR2X1 _11372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1460_),
    .B(_1461_),
    .Y(_1462_)
);

NOR2X1 _11373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [17]),
    .B(\datapath.regimmalu [17]),
    .Y(_1463_)
);

NOR2X1 _11374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1463_),
    .B(_1462_),
    .Y(_1464_)
);

XNOR2X1 _11375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1459_),
    .B(_1464_),
    .Y(\datapath.jumptarget [17])
);

OAI21X1 _11376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [17]),
    .B(\datapath.regimmalu [17]),
    .C(_1458_),
    .Y(_1465_)
);

OAI21X1 _11377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1460_),
    .B(_1461_),
    .C(_1465_),
    .Y(_1466_)
);

NAND2X1 _11378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1456_),
    .B(_1464_),
    .Y(_1467_)
);

INVX1 _11379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1467_),
    .Y(_1468_)
);

AOI21X1 _11380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1468_),
    .B(_1451_),
    .C(_1466_),
    .Y(_1469_)
);

NAND2X1 _11381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [18]),
    .B(\datapath.regimmalu [18]),
    .Y(_1470_)
);

OR2X2 _11382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [18]),
    .B(\datapath.regimmalu [18]),
    .Y(_1471_)
);

NAND2X1 _11383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1470_),
    .B(_1471_),
    .Y(_1472_)
);

INVX2 _11384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1472_),
    .Y(_1473_)
);

XNOR2X1 _11385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1469_),
    .B(_1473_),
    .Y(\datapath.jumptarget [18])
);

OAI21X1 _11386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1469_),
    .B(_1472_),
    .C(_1470_),
    .Y(_1474_)
);

AND2X2 _11387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [19]),
    .B(\datapath.regimmalu [19]),
    .Y(_1475_)
);

NOR2X1 _11388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [19]),
    .B(\datapath.regimmalu [19]),
    .Y(_1476_)
);

NOR2X1 _11389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1476_),
    .B(_1475_),
    .Y(_1477_)
);

INVX1 _11390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1477_),
    .Y(_1478_)
);

XNOR2X1 _11391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1474_),
    .B(_1478_),
    .Y(\datapath.jumptarget [19])
);

NAND3X1 _11392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1473_),
    .B(_1477_),
    .C(_1466_),
    .Y(_1479_)
);

NOR2X1 _11393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1470_),
    .B(_1476_),
    .Y(_1480_)
);

NOR2X1 _11394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1475_),
    .B(_1480_),
    .Y(_1481_)
);

NAND2X1 _11395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1481_),
    .B(_1479_),
    .Y(_1482_)
);

NAND2X1 _11396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1477_),
    .B(_1473_),
    .Y(_1483_)
);

NOR2X1 _11397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1467_),
    .B(_1483_),
    .Y(_1484_)
);

AOI21X1 _11398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1484_),
    .B(_1451_),
    .C(_1482_),
    .Y(_1485_)
);

NAND2X1 _11399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [20]),
    .B(\datapath.regimmalu [20]),
    .Y(_1486_)
);

OR2X2 _11400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [20]),
    .B(\datapath.regimmalu [20]),
    .Y(_1487_)
);

AND2X2 _11401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1487_),
    .B(_1486_),
    .Y(_1488_)
);

XNOR2X1 _11402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1485_),
    .B(_1488_),
    .Y(\datapath.jumptarget [20])
);

INVX1 _11403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1488_),
    .Y(_1489_)
);

OAI21X1 _11404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1485_),
    .B(_1489_),
    .C(_1486_),
    .Y(_1490_)
);

AND2X2 _11405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [21]),
    .B(\datapath.regimmalu [21]),
    .Y(_1491_)
);

NOR2X1 _11406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [21]),
    .B(\datapath.regimmalu [21]),
    .Y(_1492_)
);

NOR2X1 _11407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1492_),
    .B(_1491_),
    .Y(_1493_)
);

XOR2X1 _11408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1490_),
    .B(_1493_),
    .Y(\datapath.jumptarget [21])
);

NOR2X1 _11409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1486_),
    .B(_1492_),
    .Y(_1494_)
);

NOR2X1 _11410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1491_),
    .B(_1494_),
    .Y(_1495_)
);

NAND2X1 _11411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1493_),
    .B(_1488_),
    .Y(_1496_)
);

OAI21X1 _11412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1485_),
    .B(_1496_),
    .C(_1495_),
    .Y(_1497_)
);

AND2X2 _11413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [22]),
    .B(\datapath.regimmalu [22]),
    .Y(_1498_)
);

NOR2X1 _11414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [22]),
    .B(\datapath.regimmalu [22]),
    .Y(_1499_)
);

NOR2X1 _11415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1499_),
    .B(_1498_),
    .Y(_1500_)
);

XOR2X1 _11416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1497_),
    .B(_1500_),
    .Y(\datapath.jumptarget [22])
);

AOI21X1 _11417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1500_),
    .B(_1497_),
    .C(_1498_),
    .Y(_1501_)
);

AND2X2 _11418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [23]),
    .B(\datapath.regimmalu [23]),
    .Y(_1502_)
);

NOR2X1 _11419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [23]),
    .B(\datapath.regimmalu [23]),
    .Y(_1503_)
);

NOR2X1 _11420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1503_),
    .B(_1502_),
    .Y(_1504_)
);

XNOR2X1 _11421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1501_),
    .B(_1504_),
    .Y(\datapath.jumptarget [23])
);

AND2X2 _11422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1446_),
    .B(_1423_),
    .Y(_1505_)
);

OAI21X1 _11423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1392_),
    .B(_1397_),
    .C(_1505_),
    .Y(_1506_)
);

NAND2X1 _11424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1500_),
    .B(_1504_),
    .Y(_1507_)
);

NOR2X1 _11425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1507_),
    .B(_1496_),
    .Y(_1508_)
);

NAND2X1 _11426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1508_),
    .B(_1484_),
    .Y(_1509_)
);

AOI21X1 _11427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1450_),
    .B(_1506_),
    .C(_1509_),
    .Y(_1510_)
);

OR2X2 _11428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1496_),
    .B(_1507_),
    .Y(_1511_)
);

AOI21X1 _11429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1481_),
    .B(_1479_),
    .C(_1511_),
    .Y(_1512_)
);

AOI21X1 _11430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1498_),
    .B(_1504_),
    .C(_1502_),
    .Y(_1513_)
);

OAI21X1 _11431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1507_),
    .B(_1495_),
    .C(_1513_),
    .Y(_1514_)
);

OR2X2 _11432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1512_),
    .B(_1514_),
    .Y(_1515_)
);

NOR2X1 _11433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1515_),
    .B(_1510_),
    .Y(_1516_)
);

INVX1 _11434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [24]),
    .Y(_1517_)
);

INVX1 _11435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regimmalu [24]),
    .Y(_1518_)
);

NOR2X1 _11436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1517_),
    .B(_1518_),
    .Y(_1519_)
);

INVX2 _11437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1519_),
    .Y(_1520_)
);

NAND2X1 _11438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1517_),
    .B(_1518_),
    .Y(_1521_)
);

AND2X2 _11439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1520_),
    .B(_1521_),
    .Y(_1522_)
);

XNOR2X1 _11440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1516_),
    .B(_1522_),
    .Y(\datapath.jumptarget [24])
);

INVX1 _11441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1522_),
    .Y(_1523_)
);

OAI21X1 _11442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1516_),
    .B(_1523_),
    .C(_1520_),
    .Y(_1524_)
);

NAND2X1 _11443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [25]),
    .B(\datapath.regimmalu [25]),
    .Y(_1525_)
);

INVX1 _11444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1525_),
    .Y(_1526_)
);

NOR2X1 _11445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [25]),
    .B(\datapath.regimmalu [25]),
    .Y(_1527_)
);

NOR2X1 _11446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1527_),
    .B(_1526_),
    .Y(_1528_)
);

XOR2X1 _11447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1524_),
    .B(_1528_),
    .Y(\datapath.jumptarget [25])
);

OAI21X1 _11448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1520_),
    .B(_1527_),
    .C(_1525_),
    .Y(_1529_)
);

INVX1 _11449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1529_),
    .Y(_1530_)
);

NAND2X1 _11450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1528_),
    .B(_1522_),
    .Y(_1531_)
);

OAI21X1 _11451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1516_),
    .B(_1531_),
    .C(_1530_),
    .Y(_1532_)
);

NAND2X1 _11452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [26]),
    .B(\datapath.regimmalu [26]),
    .Y(_1533_)
);

INVX1 _11453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1533_),
    .Y(_1534_)
);

NOR2X1 _11454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [26]),
    .B(\datapath.regimmalu [26]),
    .Y(_1535_)
);

NOR2X1 _11455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1535_),
    .B(_1534_),
    .Y(_1536_)
);

XOR2X1 _11456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1532_),
    .B(_1536_),
    .Y(\datapath.jumptarget [26])
);

AOI21X1 _11457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1536_),
    .B(_1532_),
    .C(_1534_),
    .Y(_1537_)
);

NOR2X1 _11458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [27]),
    .B(\datapath.regimmalu [27]),
    .Y(_1538_)
);

NAND2X1 _11459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [27]),
    .B(\datapath.regimmalu [27]),
    .Y(_1539_)
);

INVX1 _11460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1539_),
    .Y(_1540_)
);

NOR2X1 _11461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1538_),
    .B(_1540_),
    .Y(_1541_)
);

XNOR2X1 _11462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1537_),
    .B(_1541_),
    .Y(\datapath.jumptarget [27])
);

NAND2X1 _11463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1536_),
    .B(_1541_),
    .Y(_1542_)
);

NOR2X1 _11464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1542_),
    .B(_1531_),
    .Y(_1543_)
);

INVX1 _11465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1543_),
    .Y(_1544_)
);

OAI21X1 _11466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1538_),
    .B(_1533_),
    .C(_1539_),
    .Y(_1545_)
);

INVX1 _11467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1545_),
    .Y(_1546_)
);

OAI21X1 _11468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1530_),
    .B(_1542_),
    .C(_1546_),
    .Y(_1547_)
);

INVX1 _11469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1547_),
    .Y(_1548_)
);

OAI21X1 _11470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1516_),
    .B(_1544_),
    .C(_1548_),
    .Y(_1549_)
);

NOR2X1 _11471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [28]),
    .B(\datapath.regimmalu [28]),
    .Y(_1550_)
);

NAND2X1 _11472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [28]),
    .B(\datapath.regimmalu [28]),
    .Y(_1551_)
);

INVX1 _11473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1551_),
    .Y(_1552_)
);

NOR2X1 _11474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1550_),
    .B(_1552_),
    .Y(_1553_)
);

XOR2X1 _11475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1549_),
    .B(_1553_),
    .Y(\datapath.jumptarget [28])
);

AOI21X1 _11476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1553_),
    .B(_1549_),
    .C(_1552_),
    .Y(_1554_)
);

NOR2X1 _11477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [29]),
    .B(\datapath.regimmalu [29]),
    .Y(_1555_)
);

NAND2X1 _11478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [29]),
    .B(\datapath.regimmalu [29]),
    .Y(_1556_)
);

INVX1 _11479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1556_),
    .Y(_1557_)
);

NOR2X1 _11480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1555_),
    .B(_1557_),
    .Y(_1558_)
);

XNOR2X1 _11481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1554_),
    .B(_1558_),
    .Y(\datapath.jumptarget [29])
);

OAI21X1 _11482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1510_),
    .B(_1515_),
    .C(_1543_),
    .Y(_1559_)
);

NAND2X1 _11483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1553_),
    .B(_1558_),
    .Y(_1560_)
);

AOI21X1 _11484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1548_),
    .B(_1559_),
    .C(_1560_),
    .Y(_1561_)
);

OAI21X1 _11485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1555_),
    .B(_1551_),
    .C(_1556_),
    .Y(_1562_)
);

NOR2X1 _11486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [30]),
    .B(\datapath.regimmalu [30]),
    .Y(_1563_)
);

NAND2X1 _11487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [30]),
    .B(\datapath.regimmalu [30]),
    .Y(_1564_)
);

INVX1 _11488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1564_),
    .Y(_1565_)
);

NOR2X1 _11489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1563_),
    .B(_1565_),
    .Y(_1566_)
);

OAI21X1 _11490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1561_),
    .B(_1562_),
    .C(_1566_),
    .Y(_1567_)
);

NOR3X1 _11491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1354_),
    .B(_1359_),
    .C(_1356_),
    .Y(_1568_)
);

INVX1 _11492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1367_),
    .Y(_1569_)
);

NOR2X1 _11493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1380_),
    .B(_1393_),
    .Y(_1570_)
);

OAI21X1 _11494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1568_),
    .B(_1569_),
    .C(_1570_),
    .Y(_1571_)
);

OAI21X1 _11495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1373_),
    .B(_1371_),
    .C(_1374_),
    .Y(_1572_)
);

AOI21X1 _11496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1390_),
    .B(_1572_),
    .C(_1395_),
    .Y(_1573_)
);

AOI21X1 _11497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1573_),
    .B(_1571_),
    .C(_1447_),
    .Y(_1574_)
);

INVX1 _11498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1450_),
    .Y(_1575_)
);

AND2X2 _11499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1484_),
    .B(_1508_),
    .Y(_1576_)
);

OAI21X1 _11500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1574_),
    .B(_1575_),
    .C(_1576_),
    .Y(_1577_)
);

NOR2X1 _11501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1514_),
    .B(_1512_),
    .Y(_1578_)
);

AOI21X1 _11502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1578_),
    .B(_1577_),
    .C(_1544_),
    .Y(_1579_)
);

INVX1 _11503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1560_),
    .Y(_1580_)
);

OAI21X1 _11504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1579_),
    .B(_1547_),
    .C(_1580_),
    .Y(_1581_)
);

INVX1 _11505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1562_),
    .Y(_1582_)
);

INVX1 _11506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1566_),
    .Y(_1583_)
);

NAND3X1 _11507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1582_),
    .B(_1583_),
    .C(_1581_),
    .Y(_1584_)
);

AND2X2 _11508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1567_),
    .B(_1584_),
    .Y(\datapath.jumptarget [30])
);

XNOR2X1 _11509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [31]),
    .B(\datapath.regimmalu [31]),
    .Y(_1585_)
);

INVX1 _11510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1585_),
    .Y(_1586_)
);

NAND3X1 _11511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1564_),
    .B(_1586_),
    .C(_1567_),
    .Y(_1587_)
);

AOI21X1 _11512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1582_),
    .B(_1581_),
    .C(_1583_),
    .Y(_1588_)
);

OAI21X1 _11513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1588_),
    .B(_1565_),
    .C(_1585_),
    .Y(_1589_)
);

NAND2X1 _11514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1589_),
    .B(_1587_),
    .Y(\datapath.jumptarget [31])
);

NOR2X1 _11515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alupc [0]),
    .B(\datapath.regimmalu [0]),
    .Y(_1590_)
);

NOR2X1 _11516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1590_),
    .B(_1347_),
    .Y(\datapath.jumptarget [0])
);

DFFPOSX1 _11517_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf153),
    .D(\datapath.regcsralu [0]),
    .Q(\datapath.regcsrmem [0])
);

DFFPOSX1 _11518_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf152),
    .D(\datapath.regcsralu [1]),
    .Q(\datapath.regcsrmem [1])
);

DFFPOSX1 _11519_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf151),
    .D(\datapath.regcsralu [2]),
    .Q(\datapath.regcsrmem [2])
);

DFFPOSX1 _11520_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf150),
    .D(\datapath.regcsralu [3]),
    .Q(\datapath.regcsrmem [3])
);

DFFPOSX1 _11521_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf149),
    .D(\datapath.regcsralu [4]),
    .Q(\datapath.regcsrmem [4])
);

DFFPOSX1 _11522_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf148),
    .D(\datapath.regcsralu [5]),
    .Q(\datapath.regcsrmem [5])
);

DFFPOSX1 _11523_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf147),
    .D(\datapath.regcsralu [6]),
    .Q(\datapath.regcsrmem [6])
);

DFFPOSX1 _11524_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf146),
    .D(\datapath.regcsralu [7]),
    .Q(\datapath.regcsrmem [7])
);

DFFPOSX1 _11525_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf145),
    .D(\datapath.regcsralu [8]),
    .Q(\datapath.regcsrmem [8])
);

DFFPOSX1 _11526_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf144),
    .D(\datapath.regcsralu [9]),
    .Q(\datapath.regcsrmem [9])
);

DFFPOSX1 _11527_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf143),
    .D(\datapath.regcsralu [10]),
    .Q(\datapath.regcsrmem [10])
);

DFFPOSX1 _11528_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf142),
    .D(\datapath.regcsralu [11]),
    .Q(\datapath.regcsrmem [11])
);

DFFPOSX1 _11529_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf141),
    .D(\datapath.regcsralu [12]),
    .Q(\datapath.regcsrmem [12])
);

DFFPOSX1 _11530_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf140),
    .D(\datapath.regcsralu [13]),
    .Q(\datapath.regcsrmem [13])
);

DFFPOSX1 _11531_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf139),
    .D(\datapath.regcsralu [14]),
    .Q(\datapath.regcsrmem [14])
);

DFFPOSX1 _11532_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf138),
    .D(\datapath.regcsralu [15]),
    .Q(\datapath.regcsrmem [15])
);

DFFPOSX1 _11533_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf137),
    .D(\datapath.regcsralu [16]),
    .Q(\datapath.regcsrmem [16])
);

DFFPOSX1 _11534_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf136),
    .D(\datapath.regcsralu [17]),
    .Q(\datapath.regcsrmem [17])
);

DFFPOSX1 _11535_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf135),
    .D(\datapath.regcsralu [18]),
    .Q(\datapath.regcsrmem [18])
);

DFFPOSX1 _11536_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf134),
    .D(\datapath.regcsralu [19]),
    .Q(\datapath.regcsrmem [19])
);

DFFPOSX1 _11537_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf133),
    .D(\datapath.regcsralu [20]),
    .Q(\datapath.regcsrmem [20])
);

DFFPOSX1 _11538_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf132),
    .D(\datapath.regcsralu [21]),
    .Q(\datapath.regcsrmem [21])
);

DFFPOSX1 _11539_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf131),
    .D(\datapath.regcsralu [22]),
    .Q(\datapath.regcsrmem [22])
);

DFFPOSX1 _11540_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf130),
    .D(\datapath.regcsralu [23]),
    .Q(\datapath.regcsrmem [23])
);

DFFPOSX1 _11541_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf129),
    .D(\datapath.regcsralu [24]),
    .Q(\datapath.regcsrmem [24])
);

DFFPOSX1 _11542_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf128),
    .D(\datapath.regcsralu [25]),
    .Q(\datapath.regcsrmem [25])
);

DFFPOSX1 _11543_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf127),
    .D(\datapath.regcsralu [26]),
    .Q(\datapath.regcsrmem [26])
);

DFFPOSX1 _11544_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf126),
    .D(\datapath.regcsralu [27]),
    .Q(\datapath.regcsrmem [27])
);

DFFPOSX1 _11545_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf125),
    .D(\datapath.regcsralu [28]),
    .Q(\datapath.regcsrmem [28])
);

DFFPOSX1 _11546_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf124),
    .D(\datapath.regcsralu [29]),
    .Q(\datapath.regcsrmem [29])
);

DFFPOSX1 _11547_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf123),
    .D(\datapath.regcsralu [30]),
    .Q(\datapath.regcsrmem [30])
);

DFFPOSX1 _11548_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf122),
    .D(\datapath.regcsralu [31]),
    .Q(\datapath.regcsrmem [31])
);

DFFPOSX1 _11549_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf121),
    .D(\datapath.regrs2alu [0]),
    .Q(\datapath.memoryinterface.data_store [0])
);

DFFPOSX1 _11550_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf120),
    .D(\datapath.regrs2alu [1]),
    .Q(\datapath.memoryinterface.data_store [1])
);

DFFPOSX1 _11551_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf119),
    .D(\datapath.regrs2alu [2]),
    .Q(\datapath.memoryinterface.data_store [2])
);

DFFPOSX1 _11552_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf118),
    .D(\datapath.regrs2alu [3]),
    .Q(\datapath.memoryinterface.data_store [3])
);

DFFPOSX1 _11553_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf117),
    .D(\datapath.regrs2alu [4]),
    .Q(\datapath.memoryinterface.data_store [4])
);

DFFPOSX1 _11554_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf116),
    .D(\datapath.regrs2alu [5]),
    .Q(\datapath.memoryinterface.data_store [5])
);

DFFPOSX1 _11555_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf115),
    .D(\datapath.regrs2alu [6]),
    .Q(\datapath.memoryinterface.data_store [6])
);

DFFPOSX1 _11556_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf114),
    .D(\datapath.regrs2alu [7]),
    .Q(\datapath.memoryinterface.data_store [7])
);

DFFPOSX1 _11557_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf113),
    .D(\datapath.regrs2alu [8]),
    .Q(\datapath.memoryinterface.data_store [8])
);

DFFPOSX1 _11558_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf112),
    .D(\datapath.regrs2alu [9]),
    .Q(\datapath.memoryinterface.data_store [9])
);

DFFPOSX1 _11559_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf111),
    .D(\datapath.regrs2alu [10]),
    .Q(\datapath.memoryinterface.data_store [10])
);

DFFPOSX1 _11560_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf110),
    .D(\datapath.regrs2alu [11]),
    .Q(\datapath.memoryinterface.data_store [11])
);

DFFPOSX1 _11561_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf109),
    .D(\datapath.regrs2alu [12]),
    .Q(\datapath.memoryinterface.data_store [12])
);

DFFPOSX1 _11562_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf108),
    .D(\datapath.regrs2alu [13]),
    .Q(\datapath.memoryinterface.data_store [13])
);

DFFPOSX1 _11563_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf107),
    .D(\datapath.regrs2alu [14]),
    .Q(\datapath.memoryinterface.data_store [14])
);

DFFPOSX1 _11564_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf106),
    .D(\datapath.regrs2alu [15]),
    .Q(\datapath.memoryinterface.data_store [15])
);

DFFPOSX1 _11565_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf105),
    .D(\datapath.regrs2alu [16]),
    .Q(\datapath.memoryinterface.data_store [16])
);

DFFPOSX1 _11566_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf104),
    .D(\datapath.regrs2alu [17]),
    .Q(\datapath.memoryinterface.data_store [17])
);

DFFPOSX1 _11567_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf103),
    .D(\datapath.regrs2alu [18]),
    .Q(\datapath.memoryinterface.data_store [18])
);

DFFPOSX1 _11568_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf102),
    .D(\datapath.regrs2alu [19]),
    .Q(\datapath.memoryinterface.data_store [19])
);

DFFPOSX1 _11569_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf101),
    .D(\datapath.regrs2alu [20]),
    .Q(\datapath.memoryinterface.data_store [20])
);

DFFPOSX1 _11570_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf100),
    .D(\datapath.regrs2alu [21]),
    .Q(\datapath.memoryinterface.data_store [21])
);

DFFPOSX1 _11571_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf99),
    .D(\datapath.regrs2alu [22]),
    .Q(\datapath.memoryinterface.data_store [22])
);

DFFPOSX1 _11572_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf98),
    .D(\datapath.regrs2alu [23]),
    .Q(\datapath.memoryinterface.data_store [23])
);

DFFPOSX1 _11573_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf97),
    .D(\datapath.regrs2alu [24]),
    .Q(\datapath.memoryinterface.data_store [24])
);

DFFPOSX1 _11574_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf96),
    .D(\datapath.regrs2alu [25]),
    .Q(\datapath.memoryinterface.data_store [25])
);

DFFPOSX1 _11575_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf95),
    .D(\datapath.regrs2alu [26]),
    .Q(\datapath.memoryinterface.data_store [26])
);

DFFPOSX1 _11576_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf94),
    .D(\datapath.regrs2alu [27]),
    .Q(\datapath.memoryinterface.data_store [27])
);

DFFPOSX1 _11577_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf93),
    .D(\datapath.regrs2alu [28]),
    .Q(\datapath.memoryinterface.data_store [28])
);

DFFPOSX1 _11578_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf92),
    .D(\datapath.regrs2alu [29]),
    .Q(\datapath.memoryinterface.data_store [29])
);

DFFPOSX1 _11579_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf91),
    .D(\datapath.regrs2alu [30]),
    .Q(\datapath.memoryinterface.data_store [30])
);

DFFPOSX1 _11580_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf90),
    .D(\datapath.regrs2alu [31]),
    .Q(\datapath.memoryinterface.data_store [31])
);

DFFPOSX1 _11581_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf89),
    .D(\datapath.alu.condtrue ),
    .Q(_0_[0])
);

DFFPOSX1 _11582_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf88),
    .D(\datapath.alu.c [1]),
    .Q(_0_[1])
);

DFFPOSX1 _11583_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf87),
    .D(\datapath.alu.c [2]),
    .Q(_0_[2])
);

DFFPOSX1 _11584_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf86),
    .D(\datapath.alu.c [3]),
    .Q(_0_[3])
);

DFFPOSX1 _11585_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf85),
    .D(\datapath.alu.c [4]),
    .Q(_0_[4])
);

DFFPOSX1 _11586_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf84),
    .D(\datapath.alu.c [5]),
    .Q(_0_[5])
);

DFFPOSX1 _11587_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf83),
    .D(\datapath.alu.c [6]),
    .Q(_0_[6])
);

DFFPOSX1 _11588_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf82),
    .D(\datapath.alu.c [7]),
    .Q(_0_[7])
);

DFFPOSX1 _11589_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf81),
    .D(\datapath.alu.c [8]),
    .Q(_0_[8])
);

DFFPOSX1 _11590_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf80),
    .D(\datapath.alu.c [9]),
    .Q(_0_[9])
);

DFFPOSX1 _11591_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf79),
    .D(\datapath.alu.c [10]),
    .Q(_0_[10])
);

DFFPOSX1 _11592_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf78),
    .D(\datapath.alu.c [11]),
    .Q(_0_[11])
);

DFFPOSX1 _11593_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf77),
    .D(\datapath.alu.c [12]),
    .Q(_0_[12])
);

DFFPOSX1 _11594_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf76),
    .D(\datapath.alu.c [13]),
    .Q(_0_[13])
);

DFFPOSX1 _11595_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf75),
    .D(\datapath.alu.c [14]),
    .Q(_0_[14])
);

DFFPOSX1 _11596_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf74),
    .D(\datapath.alu.c [15]),
    .Q(_0_[15])
);

DFFPOSX1 _11597_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf73),
    .D(\datapath.alu.c [16]),
    .Q(_0_[16])
);

DFFPOSX1 _11598_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf72),
    .D(\datapath.alu.c [17]),
    .Q(_0_[17])
);

DFFPOSX1 _11599_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf71),
    .D(\datapath.alu.c [18]),
    .Q(_0_[18])
);

DFFPOSX1 _11600_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf70),
    .D(\datapath.alu.c [19]),
    .Q(_0_[19])
);

DFFPOSX1 _11601_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf69),
    .D(\datapath.alu.c [20]),
    .Q(_0_[20])
);

DFFPOSX1 _11602_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf68),
    .D(\datapath.alu.c [21]),
    .Q(_0_[21])
);

DFFPOSX1 _11603_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf67),
    .D(\datapath.alu.c [22]),
    .Q(_0_[22])
);

DFFPOSX1 _11604_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf66),
    .D(\datapath.alu.c [23]),
    .Q(_0_[23])
);

DFFPOSX1 _11605_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf65),
    .D(\datapath.alu.c [24]),
    .Q(_0_[24])
);

DFFPOSX1 _11606_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf64),
    .D(\datapath.alu.c [25]),
    .Q(_0_[25])
);

DFFPOSX1 _11607_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf63),
    .D(\datapath.alu.c [26]),
    .Q(_0_[26])
);

DFFPOSX1 _11608_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf62),
    .D(\datapath.alu.c [27]),
    .Q(_0_[27])
);

DFFPOSX1 _11609_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf61),
    .D(\datapath.alu.c [28]),
    .Q(_0_[28])
);

DFFPOSX1 _11610_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf60),
    .D(\datapath.alu.c [29]),
    .Q(_0_[29])
);

DFFPOSX1 _11611_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf59),
    .D(\datapath.alu.c [30]),
    .Q(_0_[30])
);

DFFPOSX1 _11612_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf58),
    .D(\datapath.alu.c [31]),
    .Q(_0_[31])
);

DFFPOSX1 _11613_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf57),
    .D(\datapath.jumptarget [0]),
    .Q(\datapath.programcounter.jumps [0])
);

DFFPOSX1 _11614_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf56),
    .D(\datapath.jumptarget [1]),
    .Q(\datapath.programcounter.jumps [1])
);

DFFPOSX1 _11615_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf55),
    .D(\datapath.jumptarget [2]),
    .Q(\datapath.programcounter.jumps [2])
);

DFFPOSX1 _11616_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf54),
    .D(\datapath.jumptarget [3]),
    .Q(\datapath.programcounter.jumps [3])
);

DFFPOSX1 _11617_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf53),
    .D(\datapath.jumptarget [4]),
    .Q(\datapath.programcounter.jumps [4])
);

DFFPOSX1 _11618_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf52),
    .D(\datapath.jumptarget [5]),
    .Q(\datapath.programcounter.jumps [5])
);

DFFPOSX1 _11619_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf51),
    .D(\datapath.jumptarget [6]),
    .Q(\datapath.programcounter.jumps [6])
);

DFFPOSX1 _11620_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf50),
    .D(\datapath.jumptarget [7]),
    .Q(\datapath.programcounter.jumps [7])
);

DFFPOSX1 _11621_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf49),
    .D(\datapath.jumptarget [8]),
    .Q(\datapath.programcounter.jumps [8])
);

DFFPOSX1 _11622_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf48),
    .D(\datapath.jumptarget [9]),
    .Q(\datapath.programcounter.jumps [9])
);

DFFPOSX1 _11623_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf47),
    .D(\datapath.jumptarget [10]),
    .Q(\datapath.programcounter.jumps [10])
);

DFFPOSX1 _11624_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf46),
    .D(\datapath.jumptarget [11]),
    .Q(\datapath.programcounter.jumps [11])
);

DFFPOSX1 _11625_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf45),
    .D(\datapath.jumptarget [12]),
    .Q(\datapath.programcounter.jumps [12])
);

DFFPOSX1 _11626_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf44),
    .D(\datapath.jumptarget [13]),
    .Q(\datapath.programcounter.jumps [13])
);

DFFPOSX1 _11627_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf43),
    .D(\datapath.jumptarget [14]),
    .Q(\datapath.programcounter.jumps [14])
);

DFFPOSX1 _11628_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf42),
    .D(\datapath.jumptarget [15]),
    .Q(\datapath.programcounter.jumps [15])
);

DFFPOSX1 _11629_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf41),
    .D(\datapath.jumptarget [16]),
    .Q(\datapath.programcounter.jumps [16])
);

DFFPOSX1 _11630_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf40),
    .D(\datapath.jumptarget [17]),
    .Q(\datapath.programcounter.jumps [17])
);

DFFPOSX1 _11631_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf39),
    .D(\datapath.jumptarget [18]),
    .Q(\datapath.programcounter.jumps [18])
);

DFFPOSX1 _11632_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf38),
    .D(\datapath.jumptarget [19]),
    .Q(\datapath.programcounter.jumps [19])
);

DFFPOSX1 _11633_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf37),
    .D(\datapath.jumptarget [20]),
    .Q(\datapath.programcounter.jumps [20])
);

DFFPOSX1 _11634_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf36),
    .D(\datapath.jumptarget [21]),
    .Q(\datapath.programcounter.jumps [21])
);

DFFPOSX1 _11635_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf35),
    .D(\datapath.jumptarget [22]),
    .Q(\datapath.programcounter.jumps [22])
);

DFFPOSX1 _11636_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf34),
    .D(\datapath.jumptarget [23]),
    .Q(\datapath.programcounter.jumps [23])
);

DFFPOSX1 _11637_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf33),
    .D(\datapath.jumptarget [24]),
    .Q(\datapath.programcounter.jumps [24])
);

DFFPOSX1 _11638_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf32),
    .D(\datapath.jumptarget [25]),
    .Q(\datapath.programcounter.jumps [25])
);

DFFPOSX1 _11639_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf31),
    .D(\datapath.jumptarget [26]),
    .Q(\datapath.programcounter.jumps [26])
);

DFFPOSX1 _11640_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf30),
    .D(\datapath.jumptarget [27]),
    .Q(\datapath.programcounter.jumps [27])
);

DFFPOSX1 _11641_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf29),
    .D(\datapath.jumptarget [28]),
    .Q(\datapath.programcounter.jumps [28])
);

DFFPOSX1 _11642_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf28),
    .D(\datapath.jumptarget [29]),
    .Q(\datapath.programcounter.jumps [29])
);

DFFPOSX1 _11643_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf27),
    .D(\datapath.jumptarget [30]),
    .Q(\datapath.programcounter.jumps [30])
);

DFFPOSX1 _11644_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf26),
    .D(\datapath.jumptarget [31]),
    .Q(\datapath.programcounter.jumps [31])
);

DFFPOSX1 _11645_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf25),
    .D(\datapath._32_ [0]),
    .Q(\datapath.regpcsel [0])
);

DFFPOSX1 _11646_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf24),
    .D(\datapath._32_ [1]),
    .Q(\datapath.regpcsel [1])
);

DFFPOSX1 _11647_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf23),
    .D(\datapath.alu.condtrue ),
    .Q(\datapath.regcondt )
);

DFFPOSX1 _11648_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf22),
    .D(\datapath.alu.z ),
    .Q(\datapath.regz )
);

DFFPOSX1 _11649_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf21),
    .D(\datapath._31_ [0]),
    .Q(\datapath.memexecptions [0])
);

DFFPOSX1 _11650_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf20),
    .D(\datapath._31_ [1]),
    .Q(\datapath.memexecptions [1])
);

DFFPOSX1 _11651_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf19),
    .D(\datapath._31_ [2]),
    .Q(\datapath.memexecptions [2])
);

DFFPOSX1 _11652_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf18),
    .D(\datapath._30_ [0]),
    .Q(\datapath.meminstr [0])
);

DFFPOSX1 _11653_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf17),
    .D(\datapath._30_ [1]),
    .Q(\datapath.meminstr [1])
);

DFFPOSX1 _11654_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf16),
    .D(\datapath._30_ [2]),
    .Q(\datapath.meminstr [2])
);

DFFPOSX1 _11655_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf15),
    .D(\datapath._30_ [3]),
    .Q(\datapath.meminstr [3])
);

DFFPOSX1 _11656_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf14),
    .D(\datapath._30_ [4]),
    .Q(\datapath.meminstr [4])
);

DFFPOSX1 _11657_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf13),
    .D(\datapath._30_ [5]),
    .Q(\datapath.meminstr [5])
);

DFFPOSX1 _11658_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf12),
    .D(\datapath._30_ [6]),
    .Q(\datapath.meminstr [6])
);

DFFPOSX1 _11659_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf11),
    .D(\datapath._30_ [7]),
    .Q(\datapath.meminstr [7])
);

DFFPOSX1 _11660_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf10),
    .D(\datapath._30_ [8]),
    .Q(\datapath.meminstr [8])
);

DFFPOSX1 _11661_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf9),
    .D(\datapath._30_ [9]),
    .Q(\datapath.meminstr [9])
);

DFFPOSX1 _11662_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf8),
    .D(\datapath._30_ [10]),
    .Q(\datapath.meminstr [10])
);

DFFPOSX1 _11663_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf7),
    .D(\datapath._30_ [11]),
    .Q(\datapath.meminstr [11])
);

DFFPOSX1 _11664_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf6),
    .D(\datapath._30_ [12]),
    .Q(\datapath.meminstr [12])
);

DFFPOSX1 _11665_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf5),
    .D(\datapath._30_ [13]),
    .Q(\datapath.meminstr [13])
);

DFFPOSX1 _11666_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf4),
    .D(\datapath._30_ [14]),
    .Q(\datapath.meminstr [14])
);

DFFPOSX1 _11667_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf3),
    .D(\datapath._30_ [15]),
    .Q(\datapath.meminstr [15])
);

DFFPOSX1 _11668_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf2),
    .D(\datapath._30_ [16]),
    .Q(\datapath.meminstr [16])
);

DFFPOSX1 _11669_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf1),
    .D(\datapath._30_ [17]),
    .Q(\datapath.meminstr [17])
);

DFFPOSX1 _11670_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf0),
    .D(\datapath._30_ [18]),
    .Q(\datapath.meminstr [18])
);

DFFPOSX1 _11671_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf153),
    .D(\datapath._30_ [19]),
    .Q(\datapath.meminstr [19])
);

DFFPOSX1 _11672_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf152),
    .D(\datapath._30_ [20]),
    .Q(\datapath.meminstr [20])
);

DFFPOSX1 _11673_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf151),
    .D(\datapath._30_ [21]),
    .Q(\datapath.meminstr [21])
);

DFFPOSX1 _11674_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf150),
    .D(\datapath._30_ [22]),
    .Q(\datapath.meminstr [22])
);

DFFPOSX1 _11675_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf149),
    .D(\datapath._30_ [23]),
    .Q(\datapath.meminstr [23])
);

DFFPOSX1 _11676_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf148),
    .D(\datapath._30_ [24]),
    .Q(\datapath.meminstr [24])
);

DFFPOSX1 _11677_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf147),
    .D(\datapath._30_ [25]),
    .Q(\datapath.meminstr [25])
);

DFFPOSX1 _11678_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf146),
    .D(\datapath._30_ [26]),
    .Q(\datapath.meminstr [26])
);

DFFPOSX1 _11679_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf145),
    .D(\datapath._30_ [27]),
    .Q(\datapath.meminstr [27])
);

DFFPOSX1 _11680_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf144),
    .D(\datapath._30_ [28]),
    .Q(\datapath.meminstr [28])
);

DFFPOSX1 _11681_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf143),
    .D(\datapath._30_ [29]),
    .Q(\datapath.meminstr [29])
);

DFFPOSX1 _11682_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf142),
    .D(\datapath._30_ [30]),
    .Q(\datapath.meminstr [30])
);

DFFPOSX1 _11683_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf141),
    .D(\datapath._30_ [31]),
    .Q(\datapath.meminstr [31])
);

DFFPOSX1 _11684_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf140),
    .D(\datapath.alupc_4 [0]),
    .Q(\datapath.mempc_4 [0])
);

DFFPOSX1 _11685_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf139),
    .D(\datapath.alupc_4 [1]),
    .Q(\datapath.mempc_4 [1])
);

DFFPOSX1 _11686_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf138),
    .D(\datapath.alupc_4 [2]),
    .Q(\datapath.mempc_4 [2])
);

DFFPOSX1 _11687_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf137),
    .D(\datapath.alupc_4 [3]),
    .Q(\datapath.mempc_4 [3])
);

DFFPOSX1 _11688_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf136),
    .D(\datapath.alupc_4 [4]),
    .Q(\datapath.mempc_4 [4])
);

DFFPOSX1 _11689_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf135),
    .D(\datapath.alupc_4 [5]),
    .Q(\datapath.mempc_4 [5])
);

DFFPOSX1 _11690_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf134),
    .D(\datapath.alupc_4 [6]),
    .Q(\datapath.mempc_4 [6])
);

DFFPOSX1 _11691_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf133),
    .D(\datapath.alupc_4 [7]),
    .Q(\datapath.mempc_4 [7])
);

DFFPOSX1 _11692_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf132),
    .D(\datapath.alupc_4 [8]),
    .Q(\datapath.mempc_4 [8])
);

DFFPOSX1 _11693_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf131),
    .D(\datapath.alupc_4 [9]),
    .Q(\datapath.mempc_4 [9])
);

DFFPOSX1 _11694_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf130),
    .D(\datapath.alupc_4 [10]),
    .Q(\datapath.mempc_4 [10])
);

DFFPOSX1 _11695_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf129),
    .D(\datapath.alupc_4 [11]),
    .Q(\datapath.mempc_4 [11])
);

DFFPOSX1 _11696_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf128),
    .D(\datapath.alupc_4 [12]),
    .Q(\datapath.mempc_4 [12])
);

DFFPOSX1 _11697_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf127),
    .D(\datapath.alupc_4 [13]),
    .Q(\datapath.mempc_4 [13])
);

DFFPOSX1 _11698_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf126),
    .D(\datapath.alupc_4 [14]),
    .Q(\datapath.mempc_4 [14])
);

DFFPOSX1 _11699_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf125),
    .D(\datapath.alupc_4 [15]),
    .Q(\datapath.mempc_4 [15])
);

DFFPOSX1 _11700_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf124),
    .D(\datapath.alupc_4 [16]),
    .Q(\datapath.mempc_4 [16])
);

DFFPOSX1 _11701_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf123),
    .D(\datapath.alupc_4 [17]),
    .Q(\datapath.mempc_4 [17])
);

DFFPOSX1 _11702_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf122),
    .D(\datapath.alupc_4 [18]),
    .Q(\datapath.mempc_4 [18])
);

DFFPOSX1 _11703_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf121),
    .D(\datapath.alupc_4 [19]),
    .Q(\datapath.mempc_4 [19])
);

DFFPOSX1 _11704_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf120),
    .D(\datapath.alupc_4 [20]),
    .Q(\datapath.mempc_4 [20])
);

DFFPOSX1 _11705_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf119),
    .D(\datapath.alupc_4 [21]),
    .Q(\datapath.mempc_4 [21])
);

DFFPOSX1 _11706_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf118),
    .D(\datapath.alupc_4 [22]),
    .Q(\datapath.mempc_4 [22])
);

DFFPOSX1 _11707_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf117),
    .D(\datapath.alupc_4 [23]),
    .Q(\datapath.mempc_4 [23])
);

DFFPOSX1 _11708_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf116),
    .D(\datapath.alupc_4 [24]),
    .Q(\datapath.mempc_4 [24])
);

DFFPOSX1 _11709_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf115),
    .D(\datapath.alupc_4 [25]),
    .Q(\datapath.mempc_4 [25])
);

DFFPOSX1 _11710_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf114),
    .D(\datapath.alupc_4 [26]),
    .Q(\datapath.mempc_4 [26])
);

DFFPOSX1 _11711_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf113),
    .D(\datapath.alupc_4 [27]),
    .Q(\datapath.mempc_4 [27])
);

DFFPOSX1 _11712_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf112),
    .D(\datapath.alupc_4 [28]),
    .Q(\datapath.mempc_4 [28])
);

DFFPOSX1 _11713_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf111),
    .D(\datapath.alupc_4 [29]),
    .Q(\datapath.mempc_4 [29])
);

DFFPOSX1 _11714_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf110),
    .D(\datapath.alupc_4 [30]),
    .Q(\datapath.mempc_4 [30])
);

DFFPOSX1 _11715_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf109),
    .D(\datapath.alupc_4 [31]),
    .Q(\datapath.mempc_4 [31])
);

DFFPOSX1 _11716_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf108),
    .D(\datapath.alupc [2]),
    .Q(\datapath.mempc [2])
);

DFFPOSX1 _11717_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf107),
    .D(\datapath.alupc [3]),
    .Q(\datapath.mempc [3])
);

DFFPOSX1 _11718_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf106),
    .D(\datapath.alupc [4]),
    .Q(\datapath.mempc [4])
);

DFFPOSX1 _11719_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf105),
    .D(\datapath.alupc [5]),
    .Q(\datapath.mempc [5])
);

DFFPOSX1 _11720_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf104),
    .D(\datapath.alupc [6]),
    .Q(\datapath.mempc [6])
);

DFFPOSX1 _11721_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf103),
    .D(\datapath.alupc [7]),
    .Q(\datapath.mempc [7])
);

DFFPOSX1 _11722_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf102),
    .D(\datapath.alupc [8]),
    .Q(\datapath.mempc [8])
);

DFFPOSX1 _11723_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf101),
    .D(\datapath.alupc [9]),
    .Q(\datapath.mempc [9])
);

DFFPOSX1 _11724_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf100),
    .D(\datapath.alupc [10]),
    .Q(\datapath.mempc [10])
);

DFFPOSX1 _11725_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf99),
    .D(\datapath.alupc [11]),
    .Q(\datapath.mempc [11])
);

DFFPOSX1 _11726_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf98),
    .D(\datapath.alupc [12]),
    .Q(\datapath.mempc [12])
);

DFFPOSX1 _11727_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf97),
    .D(\datapath.alupc [13]),
    .Q(\datapath.mempc [13])
);

DFFPOSX1 _11728_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf96),
    .D(\datapath.alupc [14]),
    .Q(\datapath.mempc [14])
);

DFFPOSX1 _11729_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf95),
    .D(\datapath.alupc [15]),
    .Q(\datapath.mempc [15])
);

DFFPOSX1 _11730_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf94),
    .D(\datapath.alupc [16]),
    .Q(\datapath.mempc [16])
);

DFFPOSX1 _11731_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf93),
    .D(\datapath.alupc [17]),
    .Q(\datapath.mempc [17])
);

DFFPOSX1 _11732_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf92),
    .D(\datapath.alupc [18]),
    .Q(\datapath.mempc [18])
);

DFFPOSX1 _11733_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf91),
    .D(\datapath.alupc [19]),
    .Q(\datapath.mempc [19])
);

DFFPOSX1 _11734_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf90),
    .D(\datapath.alupc [20]),
    .Q(\datapath.mempc [20])
);

DFFPOSX1 _11735_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf89),
    .D(\datapath.alupc [21]),
    .Q(\datapath.mempc [21])
);

DFFPOSX1 _11736_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf88),
    .D(\datapath.alupc [22]),
    .Q(\datapath.mempc [22])
);

DFFPOSX1 _11737_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf87),
    .D(\datapath.alupc [23]),
    .Q(\datapath.mempc [23])
);

DFFPOSX1 _11738_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf86),
    .D(\datapath.alupc [24]),
    .Q(\datapath.mempc [24])
);

DFFPOSX1 _11739_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf85),
    .D(\datapath.alupc [25]),
    .Q(\datapath.mempc [25])
);

DFFPOSX1 _11740_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf84),
    .D(\datapath.alupc [26]),
    .Q(\datapath.mempc [26])
);

DFFPOSX1 _11741_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf83),
    .D(\datapath.alupc [27]),
    .Q(\datapath.mempc [27])
);

DFFPOSX1 _11742_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf82),
    .D(\datapath.alupc [28]),
    .Q(\datapath.mempc [28])
);

DFFPOSX1 _11743_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf81),
    .D(\datapath.alupc [29]),
    .Q(\datapath.mempc [29])
);

DFFPOSX1 _11744_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf80),
    .D(\datapath.alupc [30]),
    .Q(\datapath.mempc [30])
);

DFFPOSX1 _11745_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf79),
    .D(\datapath.alupc [31]),
    .Q(\datapath.mempc [31])
);

DFFPOSX1 _11746_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf78),
    .D(\datapath.immediatedecoder._06_ ),
    .Q(\datapath.regimmalu [0])
);

DFFPOSX1 _11747_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf77),
    .D(\datapath.imm [1]),
    .Q(\datapath.regimmalu [1])
);

DFFPOSX1 _11748_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf76),
    .D(\datapath.imm [2]),
    .Q(\datapath.regimmalu [2])
);

DFFPOSX1 _11749_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf75),
    .D(\datapath.imm [3]),
    .Q(\datapath.regimmalu [3])
);

DFFPOSX1 _11750_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf74),
    .D(\datapath.imm [4]),
    .Q(\datapath.regimmalu [4])
);

DFFPOSX1 _11751_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf73),
    .D(\datapath.imm [5]),
    .Q(\datapath.regimmalu [5])
);

DFFPOSX1 _11752_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf72),
    .D(\datapath.imm [6]),
    .Q(\datapath.regimmalu [6])
);

DFFPOSX1 _11753_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf71),
    .D(\datapath.imm [7]),
    .Q(\datapath.regimmalu [7])
);

DFFPOSX1 _11754_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf70),
    .D(\datapath.imm [8]),
    .Q(\datapath.regimmalu [8])
);

DFFPOSX1 _11755_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf69),
    .D(\datapath.imm [9]),
    .Q(\datapath.regimmalu [9])
);

DFFPOSX1 _11756_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf68),
    .D(\datapath.imm [10]),
    .Q(\datapath.regimmalu [10])
);

DFFPOSX1 _11757_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf67),
    .D(\datapath.immediatedecoder._09_ ),
    .Q(\datapath.regimmalu [11])
);

DFFPOSX1 _11758_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf66),
    .D(\datapath.imm [12]),
    .Q(\datapath.regimmalu [12])
);

DFFPOSX1 _11759_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf65),
    .D(\datapath.imm [13]),
    .Q(\datapath.regimmalu [13])
);

DFFPOSX1 _11760_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf64),
    .D(\datapath.imm [14]),
    .Q(\datapath.regimmalu [14])
);

DFFPOSX1 _11761_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf63),
    .D(\datapath.imm [15]),
    .Q(\datapath.regimmalu [15])
);

DFFPOSX1 _11762_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf62),
    .D(\datapath.imm [16]),
    .Q(\datapath.regimmalu [16])
);

DFFPOSX1 _11763_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf61),
    .D(\datapath.imm [17]),
    .Q(\datapath.regimmalu [17])
);

DFFPOSX1 _11764_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf60),
    .D(\datapath.imm [18]),
    .Q(\datapath.regimmalu [18])
);

DFFPOSX1 _11765_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf59),
    .D(\datapath.imm [19]),
    .Q(\datapath.regimmalu [19])
);

DFFPOSX1 _11766_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf58),
    .D(\datapath.imm [20]),
    .Q(\datapath.regimmalu [20])
);

DFFPOSX1 _11767_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf57),
    .D(\datapath.imm [21]),
    .Q(\datapath.regimmalu [21])
);

DFFPOSX1 _11768_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf56),
    .D(\datapath.imm [22]),
    .Q(\datapath.regimmalu [22])
);

DFFPOSX1 _11769_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf55),
    .D(\datapath.imm [23]),
    .Q(\datapath.regimmalu [23])
);

DFFPOSX1 _11770_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf54),
    .D(\datapath.imm [24]),
    .Q(\datapath.regimmalu [24])
);

DFFPOSX1 _11771_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf53),
    .D(\datapath.imm [25]),
    .Q(\datapath.regimmalu [25])
);

DFFPOSX1 _11772_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf52),
    .D(\datapath.imm [26]),
    .Q(\datapath.regimmalu [26])
);

DFFPOSX1 _11773_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf51),
    .D(\datapath.imm [27]),
    .Q(\datapath.regimmalu [27])
);

DFFPOSX1 _11774_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf50),
    .D(\datapath.imm [28]),
    .Q(\datapath.regimmalu [28])
);

DFFPOSX1 _11775_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf49),
    .D(\datapath.imm [29]),
    .Q(\datapath.regimmalu [29])
);

DFFPOSX1 _11776_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf48),
    .D(\datapath.imm [30]),
    .Q(\datapath.regimmalu [30])
);

DFFPOSX1 _11777_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf47),
    .D(\datapath.immediatedecoder._12_ ),
    .Q(\datapath.regimmalu [31])
);

DFFPOSX1 _11778_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf46),
    .D(\datapath.csr.csr_data [0]),
    .Q(\datapath.regcsralu [0])
);

DFFPOSX1 _11779_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf45),
    .D(\datapath.csr.csr_data [1]),
    .Q(\datapath.regcsralu [1])
);

DFFPOSX1 _11780_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf44),
    .D(\datapath.csr.csr_data [2]),
    .Q(\datapath.regcsralu [2])
);

DFFPOSX1 _11781_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf43),
    .D(\datapath.csr.csr_data [3]),
    .Q(\datapath.regcsralu [3])
);

DFFPOSX1 _11782_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf42),
    .D(\datapath.csr.csr_data [4]),
    .Q(\datapath.regcsralu [4])
);

DFFPOSX1 _11783_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf41),
    .D(\datapath.csr.csr_data [5]),
    .Q(\datapath.regcsralu [5])
);

DFFPOSX1 _11784_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf40),
    .D(\datapath.csr.csr_data [6]),
    .Q(\datapath.regcsralu [6])
);

DFFPOSX1 _11785_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf39),
    .D(\datapath.csr.csr_data [7]),
    .Q(\datapath.regcsralu [7])
);

DFFPOSX1 _11786_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf38),
    .D(\datapath.csr.csr_data [8]),
    .Q(\datapath.regcsralu [8])
);

DFFPOSX1 _11787_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf37),
    .D(\datapath.csr.csr_data [9]),
    .Q(\datapath.regcsralu [9])
);

DFFPOSX1 _11788_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf36),
    .D(\datapath.csr.csr_data [10]),
    .Q(\datapath.regcsralu [10])
);

DFFPOSX1 _11789_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf35),
    .D(\datapath.csr.csr_data [11]),
    .Q(\datapath.regcsralu [11])
);

DFFPOSX1 _11790_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf34),
    .D(\datapath.csr.csr_data [12]),
    .Q(\datapath.regcsralu [12])
);

DFFPOSX1 _11791_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf33),
    .D(\datapath.csr.csr_data [13]),
    .Q(\datapath.regcsralu [13])
);

DFFPOSX1 _11792_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf32),
    .D(\datapath.csr.csr_data [14]),
    .Q(\datapath.regcsralu [14])
);

DFFPOSX1 _11793_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf31),
    .D(\datapath.csr.csr_data [15]),
    .Q(\datapath.regcsralu [15])
);

DFFPOSX1 _11794_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf30),
    .D(\datapath.csr.csr_data [16]),
    .Q(\datapath.regcsralu [16])
);

DFFPOSX1 _11795_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf29),
    .D(\datapath.csr.csr_data [17]),
    .Q(\datapath.regcsralu [17])
);

DFFPOSX1 _11796_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf28),
    .D(\datapath.csr.csr_data [18]),
    .Q(\datapath.regcsralu [18])
);

DFFPOSX1 _11797_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf27),
    .D(\datapath.csr.csr_data [19]),
    .Q(\datapath.regcsralu [19])
);

DFFPOSX1 _11798_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf26),
    .D(\datapath.csr.csr_data [20]),
    .Q(\datapath.regcsralu [20])
);

DFFPOSX1 _11799_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf25),
    .D(\datapath.csr.csr_data [21]),
    .Q(\datapath.regcsralu [21])
);

DFFPOSX1 _11800_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf24),
    .D(\datapath.csr.csr_data [22]),
    .Q(\datapath.regcsralu [22])
);

DFFPOSX1 _11801_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf23),
    .D(\datapath.csr.csr_data [23]),
    .Q(\datapath.regcsralu [23])
);

DFFPOSX1 _11802_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf22),
    .D(\datapath.csr.csr_data [24]),
    .Q(\datapath.regcsralu [24])
);

DFFPOSX1 _11803_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf21),
    .D(\datapath.csr.csr_data [25]),
    .Q(\datapath.regcsralu [25])
);

DFFPOSX1 _11804_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf20),
    .D(\datapath.csr.csr_data [26]),
    .Q(\datapath.regcsralu [26])
);

DFFPOSX1 _11805_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf19),
    .D(\datapath.csr.csr_data [27]),
    .Q(\datapath.regcsralu [27])
);

DFFPOSX1 _11806_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf18),
    .D(\datapath.csr.csr_data [28]),
    .Q(\datapath.regcsralu [28])
);

DFFPOSX1 _11807_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf17),
    .D(\datapath.csr.csr_data [29]),
    .Q(\datapath.regcsralu [29])
);

DFFPOSX1 _11808_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf16),
    .D(\datapath.csr.csr_data [30]),
    .Q(\datapath.regcsralu [30])
);

DFFPOSX1 _11809_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf15),
    .D(\datapath.csr.csr_data [31]),
    .Q(\datapath.regcsralu [31])
);

DFFPOSX1 _11810_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf14),
    .D(\datapath.rs2bypass [0]),
    .Q(\datapath.regrs2alu [0])
);

DFFPOSX1 _11811_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf13),
    .D(\datapath.rs2bypass [1]),
    .Q(\datapath.regrs2alu [1])
);

DFFPOSX1 _11812_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf12),
    .D(\datapath.rs2bypass [2]),
    .Q(\datapath.regrs2alu [2])
);

DFFPOSX1 _11813_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf11),
    .D(\datapath.rs2bypass [3]),
    .Q(\datapath.regrs2alu [3])
);

DFFPOSX1 _11814_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf10),
    .D(\datapath.rs2bypass [4]),
    .Q(\datapath.regrs2alu [4])
);

DFFPOSX1 _11815_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf9),
    .D(\datapath.rs2bypass [5]),
    .Q(\datapath.regrs2alu [5])
);

DFFPOSX1 _11816_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf8),
    .D(\datapath.rs2bypass [6]),
    .Q(\datapath.regrs2alu [6])
);

DFFPOSX1 _11817_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf7),
    .D(\datapath.rs2bypass [7]),
    .Q(\datapath.regrs2alu [7])
);

DFFPOSX1 _11818_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf6),
    .D(\datapath.rs2bypass [8]),
    .Q(\datapath.regrs2alu [8])
);

DFFPOSX1 _11819_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf5),
    .D(\datapath.rs2bypass [9]),
    .Q(\datapath.regrs2alu [9])
);

DFFPOSX1 _11820_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf4),
    .D(\datapath.rs2bypass [10]),
    .Q(\datapath.regrs2alu [10])
);

DFFPOSX1 _11821_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf3),
    .D(\datapath.rs2bypass [11]),
    .Q(\datapath.regrs2alu [11])
);

DFFPOSX1 _11822_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf2),
    .D(\datapath.rs2bypass [12]),
    .Q(\datapath.regrs2alu [12])
);

DFFPOSX1 _11823_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf1),
    .D(\datapath.rs2bypass [13]),
    .Q(\datapath.regrs2alu [13])
);

DFFPOSX1 _11824_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf0),
    .D(\datapath.rs2bypass [14]),
    .Q(\datapath.regrs2alu [14])
);

DFFPOSX1 _11825_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf153),
    .D(\datapath.rs2bypass [15]),
    .Q(\datapath.regrs2alu [15])
);

DFFPOSX1 _11826_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf152),
    .D(\datapath.rs2bypass [16]),
    .Q(\datapath.regrs2alu [16])
);

DFFPOSX1 _11827_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf151),
    .D(\datapath.rs2bypass [17]),
    .Q(\datapath.regrs2alu [17])
);

DFFPOSX1 _11828_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf150),
    .D(\datapath.rs2bypass [18]),
    .Q(\datapath.regrs2alu [18])
);

DFFPOSX1 _11829_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf149),
    .D(\datapath.rs2bypass [19]),
    .Q(\datapath.regrs2alu [19])
);

DFFPOSX1 _11830_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf148),
    .D(\datapath.rs2bypass [20]),
    .Q(\datapath.regrs2alu [20])
);

DFFPOSX1 _11831_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf147),
    .D(\datapath.rs2bypass [21]),
    .Q(\datapath.regrs2alu [21])
);

DFFPOSX1 _11832_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf146),
    .D(\datapath.rs2bypass [22]),
    .Q(\datapath.regrs2alu [22])
);

DFFPOSX1 _11833_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf145),
    .D(\datapath.rs2bypass [23]),
    .Q(\datapath.regrs2alu [23])
);

DFFPOSX1 _11834_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf144),
    .D(\datapath.rs2bypass [24]),
    .Q(\datapath.regrs2alu [24])
);

DFFPOSX1 _11835_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf143),
    .D(\datapath.rs2bypass [25]),
    .Q(\datapath.regrs2alu [25])
);

DFFPOSX1 _11836_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf142),
    .D(\datapath.rs2bypass [26]),
    .Q(\datapath.regrs2alu [26])
);

DFFPOSX1 _11837_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf141),
    .D(\datapath.rs2bypass [27]),
    .Q(\datapath.regrs2alu [27])
);

DFFPOSX1 _11838_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf140),
    .D(\datapath.rs2bypass [28]),
    .Q(\datapath.regrs2alu [28])
);

DFFPOSX1 _11839_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf139),
    .D(\datapath.rs2bypass [29]),
    .Q(\datapath.regrs2alu [29])
);

DFFPOSX1 _11840_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf138),
    .D(\datapath.rs2bypass [30]),
    .Q(\datapath.regrs2alu [30])
);

DFFPOSX1 _11841_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf137),
    .D(\datapath.rs2bypass [31]),
    .Q(\datapath.regrs2alu [31])
);

DFFPOSX1 _11842_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf136),
    .D(\datapath.bbypass [0]),
    .Q(\datapath.alu.b [0])
);

DFFPOSX1 _11843_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf135),
    .D(\datapath.bbypass [1]),
    .Q(\datapath.alu.b [1])
);

DFFPOSX1 _11844_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf134),
    .D(\datapath.bbypass [2]),
    .Q(\datapath.alu.b [2])
);

DFFPOSX1 _11845_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf133),
    .D(\datapath.bbypass [3]),
    .Q(\datapath.alu.b [3])
);

DFFPOSX1 _11846_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf132),
    .D(\datapath.bbypass [4]),
    .Q(\datapath.alu.b [4])
);

DFFPOSX1 _11847_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf131),
    .D(\datapath.bbypass [5]),
    .Q(\datapath.alu.b [5])
);

DFFPOSX1 _11848_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf130),
    .D(\datapath.bbypass [6]),
    .Q(\datapath.alu.b [6])
);

DFFPOSX1 _11849_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf129),
    .D(\datapath.bbypass [7]),
    .Q(\datapath.alu.b [7])
);

DFFPOSX1 _11850_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf128),
    .D(\datapath.bbypass [8]),
    .Q(\datapath.alu.b [8])
);

DFFPOSX1 _11851_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf127),
    .D(\datapath.bbypass [9]),
    .Q(\datapath.alu.b [9])
);

DFFPOSX1 _11852_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf126),
    .D(\datapath.bbypass [10]),
    .Q(\datapath.alu.b [10])
);

DFFPOSX1 _11853_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf125),
    .D(\datapath.bbypass [11]),
    .Q(\datapath.alu.b [11])
);

DFFPOSX1 _11854_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf124),
    .D(\datapath.bbypass [12]),
    .Q(\datapath.alu.b [12])
);

DFFPOSX1 _11855_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf123),
    .D(\datapath.bbypass [13]),
    .Q(\datapath.alu.b [13])
);

DFFPOSX1 _11856_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf122),
    .D(\datapath.bbypass [14]),
    .Q(\datapath.alu.b [14])
);

DFFPOSX1 _11857_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf121),
    .D(\datapath.bbypass [15]),
    .Q(\datapath.alu.b [15])
);

DFFPOSX1 _11858_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf120),
    .D(\datapath.bbypass [16]),
    .Q(\datapath.alu.b [16])
);

DFFPOSX1 _11859_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf119),
    .D(\datapath.bbypass [17]),
    .Q(\datapath.alu.b [17])
);

DFFPOSX1 _11860_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf118),
    .D(\datapath.bbypass [18]),
    .Q(\datapath.alu.b [18])
);

DFFPOSX1 _11861_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf117),
    .D(\datapath.bbypass [19]),
    .Q(\datapath.alu.b [19])
);

DFFPOSX1 _11862_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf116),
    .D(\datapath.bbypass [20]),
    .Q(\datapath.alu.b [20])
);

DFFPOSX1 _11863_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf115),
    .D(\datapath.bbypass [21]),
    .Q(\datapath.alu.b [21])
);

DFFPOSX1 _11864_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf114),
    .D(\datapath.bbypass [22]),
    .Q(\datapath.alu.b [22])
);

DFFPOSX1 _11865_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf113),
    .D(\datapath.bbypass [23]),
    .Q(\datapath.alu.b [23])
);

DFFPOSX1 _11866_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf112),
    .D(\datapath.bbypass [24]),
    .Q(\datapath.alu.b [24])
);

DFFPOSX1 _11867_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf111),
    .D(\datapath.bbypass [25]),
    .Q(\datapath.alu.b [25])
);

DFFPOSX1 _11868_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf110),
    .D(\datapath.bbypass [26]),
    .Q(\datapath.alu.b [26])
);

DFFPOSX1 _11869_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf109),
    .D(\datapath.bbypass [27]),
    .Q(\datapath.alu.b [27])
);

DFFPOSX1 _11870_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf108),
    .D(\datapath.bbypass [28]),
    .Q(\datapath.alu.b [28])
);

DFFPOSX1 _11871_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf107),
    .D(\datapath.bbypass [29]),
    .Q(\datapath.alu.b [29])
);

DFFPOSX1 _11872_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf106),
    .D(\datapath.bbypass [30]),
    .Q(\datapath.alu.b [30])
);

DFFPOSX1 _11873_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf105),
    .D(\datapath.bbypass [31]),
    .Q(\datapath.alu.b [31])
);

DFFPOSX1 _11874_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf104),
    .D(\datapath.abypass [0]),
    .Q(\datapath.alu.a [0])
);

DFFPOSX1 _11875_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf103),
    .D(\datapath.abypass [1]),
    .Q(\datapath.alu.a [1])
);

DFFPOSX1 _11876_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf102),
    .D(\datapath.abypass [2]),
    .Q(\datapath.alu.a [2])
);

DFFPOSX1 _11877_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf101),
    .D(\datapath.abypass [3]),
    .Q(\datapath.alu.a [3])
);

DFFPOSX1 _11878_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf100),
    .D(\datapath.abypass [4]),
    .Q(\datapath.alu.a [4])
);

DFFPOSX1 _11879_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf99),
    .D(\datapath.abypass [5]),
    .Q(\datapath.alu.a [5])
);

DFFPOSX1 _11880_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf98),
    .D(\datapath.abypass [6]),
    .Q(\datapath.alu.a [6])
);

DFFPOSX1 _11881_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf97),
    .D(\datapath.abypass [7]),
    .Q(\datapath.alu.a [7])
);

DFFPOSX1 _11882_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf96),
    .D(\datapath.abypass [8]),
    .Q(\datapath.alu.a [8])
);

DFFPOSX1 _11883_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf95),
    .D(\datapath.abypass [9]),
    .Q(\datapath.alu.a [9])
);

DFFPOSX1 _11884_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf94),
    .D(\datapath.abypass [10]),
    .Q(\datapath.alu.a [10])
);

DFFPOSX1 _11885_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf93),
    .D(\datapath.abypass [11]),
    .Q(\datapath.alu.a [11])
);

DFFPOSX1 _11886_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf92),
    .D(\datapath.abypass [12]),
    .Q(\datapath.alu.a [12])
);

DFFPOSX1 _11887_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf91),
    .D(\datapath.abypass [13]),
    .Q(\datapath.alu.a [13])
);

DFFPOSX1 _11888_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf90),
    .D(\datapath.abypass [14]),
    .Q(\datapath.alu.a [14])
);

DFFPOSX1 _11889_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf89),
    .D(\datapath.abypass [15]),
    .Q(\datapath.alu.a [15])
);

DFFPOSX1 _11890_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf88),
    .D(\datapath.abypass [16]),
    .Q(\datapath.alu.a [16])
);

DFFPOSX1 _11891_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf87),
    .D(\datapath.abypass [17]),
    .Q(\datapath.alu.a [17])
);

DFFPOSX1 _11892_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf86),
    .D(\datapath.abypass [18]),
    .Q(\datapath.alu.a [18])
);

DFFPOSX1 _11893_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf85),
    .D(\datapath.abypass [19]),
    .Q(\datapath.alu.a [19])
);

DFFPOSX1 _11894_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf84),
    .D(\datapath.abypass [20]),
    .Q(\datapath.alu.a [20])
);

DFFPOSX1 _11895_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf83),
    .D(\datapath.abypass [21]),
    .Q(\datapath.alu.a [21])
);

DFFPOSX1 _11896_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf82),
    .D(\datapath.abypass [22]),
    .Q(\datapath.alu.a [22])
);

DFFPOSX1 _11897_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf81),
    .D(\datapath.abypass [23]),
    .Q(\datapath.alu.a [23])
);

DFFPOSX1 _11898_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf80),
    .D(\datapath.abypass [24]),
    .Q(\datapath.alu.a [24])
);

DFFPOSX1 _11899_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf79),
    .D(\datapath.abypass [25]),
    .Q(\datapath.alu.a [25])
);

DFFPOSX1 _11900_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf78),
    .D(\datapath.abypass [26]),
    .Q(\datapath.alu.a [26])
);

DFFPOSX1 _11901_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf77),
    .D(\datapath.abypass [27]),
    .Q(\datapath.alu.a [27])
);

DFFPOSX1 _11902_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf76),
    .D(\datapath.abypass [28]),
    .Q(\datapath.alu.a [28])
);

DFFPOSX1 _11903_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf75),
    .D(\datapath.abypass [29]),
    .Q(\datapath.alu.a [29])
);

DFFPOSX1 _11904_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf74),
    .D(\datapath.abypass [30]),
    .Q(\datapath.alu.a [30])
);

DFFPOSX1 _11905_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf73),
    .D(\datapath.abypass [31]),
    .Q(\datapath.alu.a [31])
);

DFFPOSX1 _11906_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf72),
    .D(alusel[0]),
    .Q(\datapath.alu.funsel [0])
);

DFFPOSX1 _11907_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf71),
    .D(alusel[1]),
    .Q(\datapath.alu.funsel [1])
);

DFFPOSX1 _11908_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf70),
    .D(alusel[2]),
    .Q(\datapath.alu.funsel [2])
);

DFFPOSX1 _11909_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf69),
    .D(alusel[3]),
    .Q(\datapath.alu.funsel [3])
);

DFFPOSX1 _11910_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf68),
    .D(\datapath._29_ [0]),
    .Q(\datapath.aluexecptions [0])
);

DFFPOSX1 _11911_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf67),
    .D(\datapath._29_ [1]),
    .Q(\datapath.aluexecptions [1])
);

DFFPOSX1 _11912_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf66),
    .D(\datapath._29_ [2]),
    .Q(\datapath.aluexecptions [2])
);

DFFPOSX1 _11913_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf65),
    .D(\datapath._28_ [0]),
    .Q(\datapath.aluinstr [0])
);

DFFPOSX1 _11914_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf64),
    .D(\datapath._28_ [1]),
    .Q(\datapath.aluinstr [1])
);

DFFPOSX1 _11915_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf63),
    .D(\datapath._28_ [2]),
    .Q(\datapath.aluinstr [2])
);

DFFPOSX1 _11916_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf62),
    .D(\datapath._28_ [3]),
    .Q(\datapath.aluinstr [3])
);

DFFPOSX1 _11917_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf61),
    .D(\datapath._28_ [4]),
    .Q(\datapath.aluinstr [4])
);

DFFPOSX1 _11918_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf60),
    .D(\datapath._28_ [5]),
    .Q(\datapath.aluinstr [5])
);

DFFPOSX1 _11919_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf59),
    .D(\datapath._28_ [6]),
    .Q(\datapath.aluinstr [6])
);

DFFPOSX1 _11920_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf58),
    .D(\datapath._28_ [7]),
    .Q(\datapath.aluinstr [7])
);

DFFPOSX1 _11921_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf57),
    .D(\datapath._28_ [8]),
    .Q(\datapath.aluinstr [8])
);

DFFPOSX1 _11922_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf56),
    .D(\datapath._28_ [9]),
    .Q(\datapath.aluinstr [9])
);

DFFPOSX1 _11923_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf55),
    .D(\datapath._28_ [10]),
    .Q(\datapath.aluinstr [10])
);

DFFPOSX1 _11924_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf54),
    .D(\datapath._28_ [11]),
    .Q(\datapath.aluinstr [11])
);

DFFPOSX1 _11925_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf53),
    .D(\datapath._28_ [12]),
    .Q(\datapath.aluinstr [12])
);

DFFPOSX1 _11926_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf52),
    .D(\datapath._28_ [13]),
    .Q(\datapath.aluinstr [13])
);

DFFPOSX1 _11927_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf51),
    .D(\datapath._28_ [14]),
    .Q(\datapath.aluinstr [14])
);

DFFPOSX1 _11928_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf50),
    .D(\datapath._28_ [15]),
    .Q(\datapath.aluinstr [15])
);

DFFPOSX1 _11929_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf49),
    .D(\datapath._28_ [16]),
    .Q(\datapath.aluinstr [16])
);

DFFPOSX1 _11930_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf48),
    .D(\datapath._28_ [17]),
    .Q(\datapath.aluinstr [17])
);

DFFPOSX1 _11931_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf47),
    .D(\datapath._28_ [18]),
    .Q(\datapath.aluinstr [18])
);

DFFPOSX1 _11932_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf46),
    .D(\datapath._28_ [19]),
    .Q(\datapath.aluinstr [19])
);

DFFPOSX1 _11933_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf45),
    .D(\datapath._28_ [20]),
    .Q(\datapath.aluinstr [20])
);

DFFPOSX1 _11934_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf44),
    .D(\datapath._28_ [21]),
    .Q(\datapath.aluinstr [21])
);

DFFPOSX1 _11935_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf43),
    .D(\datapath._28_ [22]),
    .Q(\datapath.aluinstr [22])
);

DFFPOSX1 _11936_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf42),
    .D(\datapath._28_ [23]),
    .Q(\datapath.aluinstr [23])
);

DFFPOSX1 _11937_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf41),
    .D(\datapath._28_ [24]),
    .Q(\datapath.aluinstr [24])
);

DFFPOSX1 _11938_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf40),
    .D(\datapath._28_ [25]),
    .Q(\datapath.aluinstr [25])
);

DFFPOSX1 _11939_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf39),
    .D(\datapath._28_ [26]),
    .Q(\datapath.aluinstr [26])
);

DFFPOSX1 _11940_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf38),
    .D(\datapath._28_ [27]),
    .Q(\datapath.aluinstr [27])
);

DFFPOSX1 _11941_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf37),
    .D(\datapath._28_ [28]),
    .Q(\datapath.aluinstr [28])
);

DFFPOSX1 _11942_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf36),
    .D(\datapath._28_ [29]),
    .Q(\datapath.aluinstr [29])
);

DFFPOSX1 _11943_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf35),
    .D(\datapath._28_ [30]),
    .Q(\datapath.aluinstr [30])
);

DFFPOSX1 _11944_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf34),
    .D(\datapath._28_ [31]),
    .Q(\datapath.aluinstr [31])
);

DFFPOSX1 _11945_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf33),
    .D(\datapath.idpc_4 [0]),
    .Q(\datapath.alupc_4 [0])
);

DFFPOSX1 _11946_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf32),
    .D(\datapath.idpc_4 [1]),
    .Q(\datapath.alupc_4 [1])
);

DFFPOSX1 _11947_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf31),
    .D(\datapath.idpc_4 [2]),
    .Q(\datapath.alupc_4 [2])
);

DFFPOSX1 _11948_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf30),
    .D(\datapath.idpc_4 [3]),
    .Q(\datapath.alupc_4 [3])
);

DFFPOSX1 _11949_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf29),
    .D(\datapath.idpc_4 [4]),
    .Q(\datapath.alupc_4 [4])
);

DFFPOSX1 _11950_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf28),
    .D(\datapath.idpc_4 [5]),
    .Q(\datapath.alupc_4 [5])
);

DFFPOSX1 _11951_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf27),
    .D(\datapath.idpc_4 [6]),
    .Q(\datapath.alupc_4 [6])
);

DFFPOSX1 _11952_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf26),
    .D(\datapath.idpc_4 [7]),
    .Q(\datapath.alupc_4 [7])
);

DFFPOSX1 _11953_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf25),
    .D(\datapath.idpc_4 [8]),
    .Q(\datapath.alupc_4 [8])
);

DFFPOSX1 _11954_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf24),
    .D(\datapath.idpc_4 [9]),
    .Q(\datapath.alupc_4 [9])
);

DFFPOSX1 _11955_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf23),
    .D(\datapath.idpc_4 [10]),
    .Q(\datapath.alupc_4 [10])
);

DFFPOSX1 _11956_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf22),
    .D(\datapath.idpc_4 [11]),
    .Q(\datapath.alupc_4 [11])
);

DFFPOSX1 _11957_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf21),
    .D(\datapath.idpc_4 [12]),
    .Q(\datapath.alupc_4 [12])
);

DFFPOSX1 _11958_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf20),
    .D(\datapath.idpc_4 [13]),
    .Q(\datapath.alupc_4 [13])
);

DFFPOSX1 _11959_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf19),
    .D(\datapath.idpc_4 [14]),
    .Q(\datapath.alupc_4 [14])
);

DFFPOSX1 _11960_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf18),
    .D(\datapath.idpc_4 [15]),
    .Q(\datapath.alupc_4 [15])
);

DFFPOSX1 _11961_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf17),
    .D(\datapath.idpc_4 [16]),
    .Q(\datapath.alupc_4 [16])
);

DFFPOSX1 _11962_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf16),
    .D(\datapath.idpc_4 [17]),
    .Q(\datapath.alupc_4 [17])
);

DFFPOSX1 _11963_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf15),
    .D(\datapath.idpc_4 [18]),
    .Q(\datapath.alupc_4 [18])
);

DFFPOSX1 _11964_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf14),
    .D(\datapath.idpc_4 [19]),
    .Q(\datapath.alupc_4 [19])
);

DFFPOSX1 _11965_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf13),
    .D(\datapath.idpc_4 [20]),
    .Q(\datapath.alupc_4 [20])
);

DFFPOSX1 _11966_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf12),
    .D(\datapath.idpc_4 [21]),
    .Q(\datapath.alupc_4 [21])
);

DFFPOSX1 _11967_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf11),
    .D(\datapath.idpc_4 [22]),
    .Q(\datapath.alupc_4 [22])
);

DFFPOSX1 _11968_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf10),
    .D(\datapath.idpc_4 [23]),
    .Q(\datapath.alupc_4 [23])
);

DFFPOSX1 _11969_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf9),
    .D(\datapath.idpc_4 [24]),
    .Q(\datapath.alupc_4 [24])
);

DFFPOSX1 _11970_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf8),
    .D(\datapath.idpc_4 [25]),
    .Q(\datapath.alupc_4 [25])
);

DFFPOSX1 _11971_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf7),
    .D(\datapath.idpc_4 [26]),
    .Q(\datapath.alupc_4 [26])
);

DFFPOSX1 _11972_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf6),
    .D(\datapath.idpc_4 [27]),
    .Q(\datapath.alupc_4 [27])
);

DFFPOSX1 _11973_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf5),
    .D(\datapath.idpc_4 [28]),
    .Q(\datapath.alupc_4 [28])
);

DFFPOSX1 _11974_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf4),
    .D(\datapath.idpc_4 [29]),
    .Q(\datapath.alupc_4 [29])
);

DFFPOSX1 _11975_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf3),
    .D(\datapath.idpc_4 [30]),
    .Q(\datapath.alupc_4 [30])
);

DFFPOSX1 _11976_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf2),
    .D(\datapath.idpc_4 [31]),
    .Q(\datapath.alupc_4 [31])
);

DFFPOSX1 _11977_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf1),
    .D(\datapath.idpc [0]),
    .Q(\datapath.alupc [0])
);

DFFPOSX1 _11978_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf0),
    .D(\datapath.idpc [1]),
    .Q(\datapath.alupc [1])
);

DFFPOSX1 _11979_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf153),
    .D(\datapath.idpc [2]),
    .Q(\datapath.alupc [2])
);

DFFPOSX1 _11980_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf152),
    .D(\datapath.idpc [3]),
    .Q(\datapath.alupc [3])
);

DFFPOSX1 _11981_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf151),
    .D(\datapath.idpc [4]),
    .Q(\datapath.alupc [4])
);

DFFPOSX1 _11982_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf150),
    .D(\datapath.idpc [5]),
    .Q(\datapath.alupc [5])
);

DFFPOSX1 _11983_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf149),
    .D(\datapath.idpc [6]),
    .Q(\datapath.alupc [6])
);

DFFPOSX1 _11984_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf148),
    .D(\datapath.idpc [7]),
    .Q(\datapath.alupc [7])
);

DFFPOSX1 _11985_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf147),
    .D(\datapath.idpc [8]),
    .Q(\datapath.alupc [8])
);

DFFPOSX1 _11986_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf146),
    .D(\datapath.idpc [9]),
    .Q(\datapath.alupc [9])
);

DFFPOSX1 _11987_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf145),
    .D(\datapath.idpc [10]),
    .Q(\datapath.alupc [10])
);

DFFPOSX1 _11988_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf144),
    .D(\datapath.idpc [11]),
    .Q(\datapath.alupc [11])
);

DFFPOSX1 _11989_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf143),
    .D(\datapath.idpc [12]),
    .Q(\datapath.alupc [12])
);

DFFPOSX1 _11990_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf142),
    .D(\datapath.idpc [13]),
    .Q(\datapath.alupc [13])
);

DFFPOSX1 _11991_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf141),
    .D(\datapath.idpc [14]),
    .Q(\datapath.alupc [14])
);

DFFPOSX1 _11992_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf140),
    .D(\datapath.idpc [15]),
    .Q(\datapath.alupc [15])
);

DFFPOSX1 _11993_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf139),
    .D(\datapath.idpc [16]),
    .Q(\datapath.alupc [16])
);

DFFPOSX1 _11994_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf138),
    .D(\datapath.idpc [17]),
    .Q(\datapath.alupc [17])
);

DFFPOSX1 _11995_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf137),
    .D(\datapath.idpc [18]),
    .Q(\datapath.alupc [18])
);

DFFPOSX1 _11996_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf136),
    .D(\datapath.idpc [19]),
    .Q(\datapath.alupc [19])
);

DFFPOSX1 _11997_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf135),
    .D(\datapath.idpc [20]),
    .Q(\datapath.alupc [20])
);

DFFPOSX1 _11998_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf134),
    .D(\datapath.idpc [21]),
    .Q(\datapath.alupc [21])
);

DFFPOSX1 _11999_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf133),
    .D(\datapath.idpc [22]),
    .Q(\datapath.alupc [22])
);

DFFPOSX1 _12000_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf132),
    .D(\datapath.idpc [23]),
    .Q(\datapath.alupc [23])
);

DFFPOSX1 _12001_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf131),
    .D(\datapath.idpc [24]),
    .Q(\datapath.alupc [24])
);

DFFPOSX1 _12002_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf130),
    .D(\datapath.idpc [25]),
    .Q(\datapath.alupc [25])
);

DFFPOSX1 _12003_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf129),
    .D(\datapath.idpc [26]),
    .Q(\datapath.alupc [26])
);

DFFPOSX1 _12004_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf128),
    .D(\datapath.idpc [27]),
    .Q(\datapath.alupc [27])
);

DFFPOSX1 _12005_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf127),
    .D(\datapath.idpc [28]),
    .Q(\datapath.alupc [28])
);

DFFPOSX1 _12006_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf126),
    .D(\datapath.idpc [29]),
    .Q(\datapath.alupc [29])
);

DFFPOSX1 _12007_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf125),
    .D(\datapath.idpc [30]),
    .Q(\datapath.alupc [30])
);

DFFPOSX1 _12008_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf124),
    .D(\datapath.idpc [31]),
    .Q(\datapath.alupc [31])
);

DFFPOSX1 _12009_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf123),
    .D(\datapath._03_ [0]),
    .Q(\datapath.idinstr [0])
);

DFFPOSX1 _12010_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf122),
    .D(\datapath._03_ [1]),
    .Q(\datapath.idinstr [1])
);

DFFPOSX1 _12011_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf121),
    .D(\datapath._03_ [2]),
    .Q(\datapath.idinstr [2])
);

DFFPOSX1 _12012_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf120),
    .D(\datapath._03_ [3]),
    .Q(\datapath.idinstr [3])
);

DFFPOSX1 _12013_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf119),
    .D(\datapath._03_ [4]),
    .Q(\datapath.idinstr [4])
);

DFFPOSX1 _12014_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf118),
    .D(\datapath._03_ [5]),
    .Q(\datapath.idinstr [5])
);

DFFPOSX1 _12015_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf117),
    .D(\datapath._03_ [6]),
    .Q(\datapath.idinstr [6])
);

DFFPOSX1 _12016_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf116),
    .D(\datapath._03_ [7]),
    .Q(\datapath.idinstr [7])
);

DFFPOSX1 _12017_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf115),
    .D(\datapath._03_ [8]),
    .Q(\datapath.idinstr [8])
);

DFFPOSX1 _12018_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf114),
    .D(\datapath._03_ [9]),
    .Q(\datapath.idinstr [9])
);

DFFPOSX1 _12019_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf113),
    .D(\datapath._03_ [10]),
    .Q(\datapath.idinstr [10])
);

DFFPOSX1 _12020_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf112),
    .D(\datapath._03_ [11]),
    .Q(\datapath.idinstr [11])
);

DFFPOSX1 _12021_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf111),
    .D(\datapath._03_ [12]),
    .Q(\datapath.idinstr [12])
);

DFFPOSX1 _12022_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf110),
    .D(\datapath._03_ [13]),
    .Q(\datapath.idinstr [13])
);

DFFPOSX1 _12023_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf109),
    .D(\datapath._03_ [14]),
    .Q(\datapath.idinstr [14])
);

DFFPOSX1 _12024_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf108),
    .D(\datapath._03_ [15]),
    .Q(\datapath.idinstr [15])
);

DFFPOSX1 _12025_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf107),
    .D(\datapath._03_ [16]),
    .Q(\datapath.idinstr [16])
);

DFFPOSX1 _12026_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf106),
    .D(\datapath._03_ [17]),
    .Q(\datapath.idinstr [17])
);

DFFPOSX1 _12027_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf105),
    .D(\datapath._03_ [18]),
    .Q(\datapath.idinstr [18])
);

DFFPOSX1 _12028_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf104),
    .D(\datapath._03_ [19]),
    .Q(\datapath.idinstr [19])
);

DFFPOSX1 _12029_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf103),
    .D(\datapath._03_ [20]),
    .Q(\datapath.idinstr [20])
);

DFFPOSX1 _12030_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf102),
    .D(\datapath._03_ [21]),
    .Q(\datapath.idinstr [21])
);

DFFPOSX1 _12031_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf101),
    .D(\datapath._03_ [22]),
    .Q(\datapath.idinstr [22])
);

DFFPOSX1 _12032_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf100),
    .D(\datapath._03_ [23]),
    .Q(\datapath.idinstr [23])
);

DFFPOSX1 _12033_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf99),
    .D(\datapath._03_ [24]),
    .Q(\datapath.idinstr [24])
);

DFFPOSX1 _12034_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf98),
    .D(\datapath._03_ [25]),
    .Q(\datapath.idinstr [25])
);

DFFPOSX1 _12035_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf97),
    .D(\datapath._03_ [26]),
    .Q(\datapath.idinstr [26])
);

DFFPOSX1 _12036_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf96),
    .D(\datapath._03_ [27]),
    .Q(\datapath.idinstr [27])
);

DFFPOSX1 _12037_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf95),
    .D(\datapath._03_ [28]),
    .Q(\datapath.idinstr [28])
);

DFFPOSX1 _12038_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf94),
    .D(\datapath._03_ [29]),
    .Q(\datapath.idinstr [29])
);

DFFPOSX1 _12039_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf93),
    .D(\datapath._03_ [30]),
    .Q(\datapath.idinstr [30])
);

DFFPOSX1 _12040_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf92),
    .D(\datapath._03_ [31]),
    .Q(\datapath.idinstr [31])
);

DFFPOSX1 _12041_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf91),
    .D(\datapath._06_ [0]),
    .Q(\datapath.idpc_4 [0])
);

DFFPOSX1 _12042_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf90),
    .D(\datapath._06_ [1]),
    .Q(\datapath.idpc_4 [1])
);

DFFPOSX1 _12043_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf89),
    .D(\datapath._06_ [2]),
    .Q(\datapath.idpc_4 [2])
);

DFFPOSX1 _12044_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf88),
    .D(\datapath._06_ [3]),
    .Q(\datapath.idpc_4 [3])
);

DFFPOSX1 _12045_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf87),
    .D(\datapath._06_ [4]),
    .Q(\datapath.idpc_4 [4])
);

DFFPOSX1 _12046_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf86),
    .D(\datapath._06_ [5]),
    .Q(\datapath.idpc_4 [5])
);

DFFPOSX1 _12047_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf85),
    .D(\datapath._06_ [6]),
    .Q(\datapath.idpc_4 [6])
);

DFFPOSX1 _12048_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf84),
    .D(\datapath._06_ [7]),
    .Q(\datapath.idpc_4 [7])
);

DFFPOSX1 _12049_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf83),
    .D(\datapath._06_ [8]),
    .Q(\datapath.idpc_4 [8])
);

DFFPOSX1 _12050_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf82),
    .D(\datapath._06_ [9]),
    .Q(\datapath.idpc_4 [9])
);

DFFPOSX1 _12051_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf81),
    .D(\datapath._06_ [10]),
    .Q(\datapath.idpc_4 [10])
);

DFFPOSX1 _12052_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf80),
    .D(\datapath._06_ [11]),
    .Q(\datapath.idpc_4 [11])
);

DFFPOSX1 _12053_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf79),
    .D(\datapath._06_ [12]),
    .Q(\datapath.idpc_4 [12])
);

DFFPOSX1 _12054_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf78),
    .D(\datapath._06_ [13]),
    .Q(\datapath.idpc_4 [13])
);

DFFPOSX1 _12055_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf77),
    .D(\datapath._06_ [14]),
    .Q(\datapath.idpc_4 [14])
);

DFFPOSX1 _12056_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf76),
    .D(\datapath._06_ [15]),
    .Q(\datapath.idpc_4 [15])
);

DFFPOSX1 _12057_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf75),
    .D(\datapath._06_ [16]),
    .Q(\datapath.idpc_4 [16])
);

DFFPOSX1 _12058_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf74),
    .D(\datapath._06_ [17]),
    .Q(\datapath.idpc_4 [17])
);

DFFPOSX1 _12059_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf73),
    .D(\datapath._06_ [18]),
    .Q(\datapath.idpc_4 [18])
);

DFFPOSX1 _12060_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf72),
    .D(\datapath._06_ [19]),
    .Q(\datapath.idpc_4 [19])
);

DFFPOSX1 _12061_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf71),
    .D(\datapath._06_ [20]),
    .Q(\datapath.idpc_4 [20])
);

DFFPOSX1 _12062_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf70),
    .D(\datapath._06_ [21]),
    .Q(\datapath.idpc_4 [21])
);

DFFPOSX1 _12063_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf69),
    .D(\datapath._06_ [22]),
    .Q(\datapath.idpc_4 [22])
);

DFFPOSX1 _12064_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf68),
    .D(\datapath._06_ [23]),
    .Q(\datapath.idpc_4 [23])
);

DFFPOSX1 _12065_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf67),
    .D(\datapath._06_ [24]),
    .Q(\datapath.idpc_4 [24])
);

DFFPOSX1 _12066_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf66),
    .D(\datapath._06_ [25]),
    .Q(\datapath.idpc_4 [25])
);

DFFPOSX1 _12067_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf65),
    .D(\datapath._06_ [26]),
    .Q(\datapath.idpc_4 [26])
);

DFFPOSX1 _12068_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf64),
    .D(\datapath._06_ [27]),
    .Q(\datapath.idpc_4 [27])
);

DFFPOSX1 _12069_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf63),
    .D(\datapath._06_ [28]),
    .Q(\datapath.idpc_4 [28])
);

DFFPOSX1 _12070_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf62),
    .D(\datapath._06_ [29]),
    .Q(\datapath.idpc_4 [29])
);

DFFPOSX1 _12071_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf61),
    .D(\datapath._06_ [30]),
    .Q(\datapath.idpc_4 [30])
);

DFFPOSX1 _12072_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf60),
    .D(\datapath._06_ [31]),
    .Q(\datapath.idpc_4 [31])
);

DFFPOSX1 _12073_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf59),
    .D(\datapath._05_ [0]),
    .Q(\datapath.idpc [0])
);

DFFPOSX1 _12074_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf58),
    .D(\datapath._05_ [1]),
    .Q(\datapath.idpc [1])
);

DFFPOSX1 _12075_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf57),
    .D(\datapath._05_ [2]),
    .Q(\datapath.idpc [2])
);

DFFPOSX1 _12076_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf56),
    .D(\datapath._05_ [3]),
    .Q(\datapath.idpc [3])
);

DFFPOSX1 _12077_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf55),
    .D(\datapath._05_ [4]),
    .Q(\datapath.idpc [4])
);

DFFPOSX1 _12078_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf54),
    .D(\datapath._05_ [5]),
    .Q(\datapath.idpc [5])
);

DFFPOSX1 _12079_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf53),
    .D(\datapath._05_ [6]),
    .Q(\datapath.idpc [6])
);

DFFPOSX1 _12080_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf52),
    .D(\datapath._05_ [7]),
    .Q(\datapath.idpc [7])
);

DFFPOSX1 _12081_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf51),
    .D(\datapath._05_ [8]),
    .Q(\datapath.idpc [8])
);

DFFPOSX1 _12082_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf50),
    .D(\datapath._05_ [9]),
    .Q(\datapath.idpc [9])
);

DFFPOSX1 _12083_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf49),
    .D(\datapath._05_ [10]),
    .Q(\datapath.idpc [10])
);

DFFPOSX1 _12084_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf48),
    .D(\datapath._05_ [11]),
    .Q(\datapath.idpc [11])
);

DFFPOSX1 _12085_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf47),
    .D(\datapath._05_ [12]),
    .Q(\datapath.idpc [12])
);

DFFPOSX1 _12086_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf46),
    .D(\datapath._05_ [13]),
    .Q(\datapath.idpc [13])
);

DFFPOSX1 _12087_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf45),
    .D(\datapath._05_ [14]),
    .Q(\datapath.idpc [14])
);

DFFPOSX1 _12088_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf44),
    .D(\datapath._05_ [15]),
    .Q(\datapath.idpc [15])
);

DFFPOSX1 _12089_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf43),
    .D(\datapath._05_ [16]),
    .Q(\datapath.idpc [16])
);

DFFPOSX1 _12090_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf42),
    .D(\datapath._05_ [17]),
    .Q(\datapath.idpc [17])
);

DFFPOSX1 _12091_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf41),
    .D(\datapath._05_ [18]),
    .Q(\datapath.idpc [18])
);

DFFPOSX1 _12092_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf40),
    .D(\datapath._05_ [19]),
    .Q(\datapath.idpc [19])
);

DFFPOSX1 _12093_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf39),
    .D(\datapath._05_ [20]),
    .Q(\datapath.idpc [20])
);

DFFPOSX1 _12094_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf38),
    .D(\datapath._05_ [21]),
    .Q(\datapath.idpc [21])
);

DFFPOSX1 _12095_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf37),
    .D(\datapath._05_ [22]),
    .Q(\datapath.idpc [22])
);

DFFPOSX1 _12096_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf36),
    .D(\datapath._05_ [23]),
    .Q(\datapath.idpc [23])
);

DFFPOSX1 _12097_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf35),
    .D(\datapath._05_ [24]),
    .Q(\datapath.idpc [24])
);

DFFPOSX1 _12098_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf34),
    .D(\datapath._05_ [25]),
    .Q(\datapath.idpc [25])
);

DFFPOSX1 _12099_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf33),
    .D(\datapath._05_ [26]),
    .Q(\datapath.idpc [26])
);

DFFPOSX1 _12100_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf32),
    .D(\datapath._05_ [27]),
    .Q(\datapath.idpc [27])
);

DFFPOSX1 _12101_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf31),
    .D(\datapath._05_ [28]),
    .Q(\datapath.idpc [28])
);

DFFPOSX1 _12102_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf30),
    .D(\datapath._05_ [29]),
    .Q(\datapath.idpc [29])
);

DFFPOSX1 _12103_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf29),
    .D(\datapath._05_ [30]),
    .Q(\datapath.idpc [30])
);

DFFPOSX1 _12104_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf28),
    .D(\datapath._05_ [31]),
    .Q(\datapath.idpc [31])
);

DFFPOSX1 _12105_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf27),
    .D(\datapath.regcsrmem [0]),
    .Q(\datapath.regcsrwb [0])
);

DFFPOSX1 _12106_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf26),
    .D(\datapath.regcsrmem [1]),
    .Q(\datapath.regcsrwb [1])
);

DFFPOSX1 _12107_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf25),
    .D(\datapath.regcsrmem [2]),
    .Q(\datapath.regcsrwb [2])
);

DFFPOSX1 _12108_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf24),
    .D(\datapath.regcsrmem [3]),
    .Q(\datapath.regcsrwb [3])
);

DFFPOSX1 _12109_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf23),
    .D(\datapath.regcsrmem [4]),
    .Q(\datapath.regcsrwb [4])
);

DFFPOSX1 _12110_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf22),
    .D(\datapath.regcsrmem [5]),
    .Q(\datapath.regcsrwb [5])
);

DFFPOSX1 _12111_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf21),
    .D(\datapath.regcsrmem [6]),
    .Q(\datapath.regcsrwb [6])
);

DFFPOSX1 _12112_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf20),
    .D(\datapath.regcsrmem [7]),
    .Q(\datapath.regcsrwb [7])
);

DFFPOSX1 _12113_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf19),
    .D(\datapath.regcsrmem [8]),
    .Q(\datapath.regcsrwb [8])
);

DFFPOSX1 _12114_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf18),
    .D(\datapath.regcsrmem [9]),
    .Q(\datapath.regcsrwb [9])
);

DFFPOSX1 _12115_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf17),
    .D(\datapath.regcsrmem [10]),
    .Q(\datapath.regcsrwb [10])
);

DFFPOSX1 _12116_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf16),
    .D(\datapath.regcsrmem [11]),
    .Q(\datapath.regcsrwb [11])
);

DFFPOSX1 _12117_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf15),
    .D(\datapath.regcsrmem [12]),
    .Q(\datapath.regcsrwb [12])
);

DFFPOSX1 _12118_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf14),
    .D(\datapath.regcsrmem [13]),
    .Q(\datapath.regcsrwb [13])
);

DFFPOSX1 _12119_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf13),
    .D(\datapath.regcsrmem [14]),
    .Q(\datapath.regcsrwb [14])
);

DFFPOSX1 _12120_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf12),
    .D(\datapath.regcsrmem [15]),
    .Q(\datapath.regcsrwb [15])
);

DFFPOSX1 _12121_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf11),
    .D(\datapath.regcsrmem [16]),
    .Q(\datapath.regcsrwb [16])
);

DFFPOSX1 _12122_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf10),
    .D(\datapath.regcsrmem [17]),
    .Q(\datapath.regcsrwb [17])
);

DFFPOSX1 _12123_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf9),
    .D(\datapath.regcsrmem [18]),
    .Q(\datapath.regcsrwb [18])
);

DFFPOSX1 _12124_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf8),
    .D(\datapath.regcsrmem [19]),
    .Q(\datapath.regcsrwb [19])
);

DFFPOSX1 _12125_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf7),
    .D(\datapath.regcsrmem [20]),
    .Q(\datapath.regcsrwb [20])
);

DFFPOSX1 _12126_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf6),
    .D(\datapath.regcsrmem [21]),
    .Q(\datapath.regcsrwb [21])
);

DFFPOSX1 _12127_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf5),
    .D(\datapath.regcsrmem [22]),
    .Q(\datapath.regcsrwb [22])
);

DFFPOSX1 _12128_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf4),
    .D(\datapath.regcsrmem [23]),
    .Q(\datapath.regcsrwb [23])
);

DFFPOSX1 _12129_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf3),
    .D(\datapath.regcsrmem [24]),
    .Q(\datapath.regcsrwb [24])
);

DFFPOSX1 _12130_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf2),
    .D(\datapath.regcsrmem [25]),
    .Q(\datapath.regcsrwb [25])
);

DFFPOSX1 _12131_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf1),
    .D(\datapath.regcsrmem [26]),
    .Q(\datapath.regcsrwb [26])
);

DFFPOSX1 _12132_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf0),
    .D(\datapath.regcsrmem [27]),
    .Q(\datapath.regcsrwb [27])
);

DFFPOSX1 _12133_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf153),
    .D(\datapath.regcsrmem [28]),
    .Q(\datapath.regcsrwb [28])
);

DFFPOSX1 _12134_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf152),
    .D(\datapath.regcsrmem [29]),
    .Q(\datapath.regcsrwb [29])
);

DFFPOSX1 _12135_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf151),
    .D(\datapath.regcsrmem [30]),
    .Q(\datapath.regcsrwb [30])
);

DFFPOSX1 _12136_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf150),
    .D(\datapath.regcsrmem [31]),
    .Q(\datapath.regcsrwb [31])
);

DFFPOSX1 _12137_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf149),
    .D(\datapath.memdataload [0]),
    .Q(\datapath.regloadwb [0])
);

DFFPOSX1 _12138_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf148),
    .D(\datapath.memdataload [1]),
    .Q(\datapath.regloadwb [1])
);

DFFPOSX1 _12139_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf147),
    .D(\datapath.memdataload [2]),
    .Q(\datapath.regloadwb [2])
);

DFFPOSX1 _12140_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf146),
    .D(\datapath.memdataload [3]),
    .Q(\datapath.regloadwb [3])
);

DFFPOSX1 _12141_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf145),
    .D(\datapath.memdataload [4]),
    .Q(\datapath.regloadwb [4])
);

DFFPOSX1 _12142_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf144),
    .D(\datapath.memdataload [5]),
    .Q(\datapath.regloadwb [5])
);

DFFPOSX1 _12143_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf143),
    .D(\datapath.memdataload [6]),
    .Q(\datapath.regloadwb [6])
);

DFFPOSX1 _12144_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf142),
    .D(\datapath.memdataload [7]),
    .Q(\datapath.regloadwb [7])
);

DFFPOSX1 _12145_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf141),
    .D(\datapath.memdataload [8]),
    .Q(\datapath.regloadwb [8])
);

DFFPOSX1 _12146_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf140),
    .D(\datapath.memdataload [9]),
    .Q(\datapath.regloadwb [9])
);

DFFPOSX1 _12147_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf139),
    .D(\datapath.memdataload [10]),
    .Q(\datapath.regloadwb [10])
);

DFFPOSX1 _12148_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf138),
    .D(\datapath.memdataload [11]),
    .Q(\datapath.regloadwb [11])
);

DFFPOSX1 _12149_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf137),
    .D(\datapath.memdataload [12]),
    .Q(\datapath.regloadwb [12])
);

DFFPOSX1 _12150_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf136),
    .D(\datapath.memdataload [13]),
    .Q(\datapath.regloadwb [13])
);

DFFPOSX1 _12151_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf135),
    .D(\datapath.memdataload [14]),
    .Q(\datapath.regloadwb [14])
);

DFFPOSX1 _12152_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf134),
    .D(\datapath.memdataload [15]),
    .Q(\datapath.regloadwb [15])
);

DFFPOSX1 _12153_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf133),
    .D(\datapath.memdataload [16]),
    .Q(\datapath.regloadwb [16])
);

DFFPOSX1 _12154_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf132),
    .D(\datapath.memdataload [17]),
    .Q(\datapath.regloadwb [17])
);

DFFPOSX1 _12155_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf131),
    .D(\datapath.memdataload [18]),
    .Q(\datapath.regloadwb [18])
);

DFFPOSX1 _12156_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf130),
    .D(\datapath.memdataload [19]),
    .Q(\datapath.regloadwb [19])
);

DFFPOSX1 _12157_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf129),
    .D(\datapath.memdataload [20]),
    .Q(\datapath.regloadwb [20])
);

DFFPOSX1 _12158_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf128),
    .D(\datapath.memdataload [21]),
    .Q(\datapath.regloadwb [21])
);

DFFPOSX1 _12159_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf127),
    .D(\datapath.memdataload [22]),
    .Q(\datapath.regloadwb [22])
);

DFFPOSX1 _12160_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf126),
    .D(\datapath.memdataload [23]),
    .Q(\datapath.regloadwb [23])
);

DFFPOSX1 _12161_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf125),
    .D(\datapath.memdataload [24]),
    .Q(\datapath.regloadwb [24])
);

DFFPOSX1 _12162_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf124),
    .D(\datapath.memdataload [25]),
    .Q(\datapath.regloadwb [25])
);

DFFPOSX1 _12163_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf123),
    .D(\datapath.memdataload [26]),
    .Q(\datapath.regloadwb [26])
);

DFFPOSX1 _12164_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf122),
    .D(\datapath.memdataload [27]),
    .Q(\datapath.regloadwb [27])
);

DFFPOSX1 _12165_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf121),
    .D(\datapath.memdataload [28]),
    .Q(\datapath.regloadwb [28])
);

DFFPOSX1 _12166_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf120),
    .D(\datapath.memdataload [29]),
    .Q(\datapath.regloadwb [29])
);

DFFPOSX1 _12167_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf119),
    .D(\datapath.memdataload [30]),
    .Q(\datapath.regloadwb [30])
);

DFFPOSX1 _12168_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf118),
    .D(\datapath.memdataload [31]),
    .Q(\datapath.regloadwb [31])
);

DFFPOSX1 _12169_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf117),
    .D(_0__0_bF$buf1),
    .Q(\datapath.regcwb [0])
);

DFFPOSX1 _12170_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf116),
    .D(_0__1_bF$buf6),
    .Q(\datapath.regcwb [1])
);

DFFPOSX1 _12171_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf115),
    .D(_0_[2]),
    .Q(\datapath.regcwb [2])
);

DFFPOSX1 _12172_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf114),
    .D(_0_[3]),
    .Q(\datapath.regcwb [3])
);

DFFPOSX1 _12173_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf113),
    .D(_0_[4]),
    .Q(\datapath.regcwb [4])
);

DFFPOSX1 _12174_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf112),
    .D(_0_[5]),
    .Q(\datapath.regcwb [5])
);

DFFPOSX1 _12175_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf111),
    .D(_0_[6]),
    .Q(\datapath.regcwb [6])
);

DFFPOSX1 _12176_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf110),
    .D(_0_[7]),
    .Q(\datapath.regcwb [7])
);

DFFPOSX1 _12177_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf109),
    .D(_0_[8]),
    .Q(\datapath.regcwb [8])
);

DFFPOSX1 _12178_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf108),
    .D(_0_[9]),
    .Q(\datapath.regcwb [9])
);

DFFPOSX1 _12179_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf107),
    .D(_0_[10]),
    .Q(\datapath.regcwb [10])
);

DFFPOSX1 _12180_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf106),
    .D(_0_[11]),
    .Q(\datapath.regcwb [11])
);

DFFPOSX1 _12181_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf105),
    .D(_0_[12]),
    .Q(\datapath.regcwb [12])
);

DFFPOSX1 _12182_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf104),
    .D(_0_[13]),
    .Q(\datapath.regcwb [13])
);

DFFPOSX1 _12183_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf103),
    .D(_0_[14]),
    .Q(\datapath.regcwb [14])
);

DFFPOSX1 _12184_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf102),
    .D(_0_[15]),
    .Q(\datapath.regcwb [15])
);

DFFPOSX1 _12185_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf101),
    .D(_0_[16]),
    .Q(\datapath.regcwb [16])
);

DFFPOSX1 _12186_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf100),
    .D(_0_[17]),
    .Q(\datapath.regcwb [17])
);

DFFPOSX1 _12187_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf99),
    .D(_0_[18]),
    .Q(\datapath.regcwb [18])
);

DFFPOSX1 _12188_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf98),
    .D(_0_[19]),
    .Q(\datapath.regcwb [19])
);

DFFPOSX1 _12189_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf97),
    .D(_0_[20]),
    .Q(\datapath.regcwb [20])
);

DFFPOSX1 _12190_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf96),
    .D(_0_[21]),
    .Q(\datapath.regcwb [21])
);

DFFPOSX1 _12191_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf95),
    .D(_0_[22]),
    .Q(\datapath.regcwb [22])
);

DFFPOSX1 _12192_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf94),
    .D(_0_[23]),
    .Q(\datapath.regcwb [23])
);

DFFPOSX1 _12193_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf93),
    .D(_0_[24]),
    .Q(\datapath.regcwb [24])
);

DFFPOSX1 _12194_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf92),
    .D(_0_[25]),
    .Q(\datapath.regcwb [25])
);

DFFPOSX1 _12195_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf91),
    .D(_0_[26]),
    .Q(\datapath.regcwb [26])
);

DFFPOSX1 _12196_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf90),
    .D(_0_[27]),
    .Q(\datapath.regcwb [27])
);

DFFPOSX1 _12197_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf89),
    .D(_0_[28]),
    .Q(\datapath.regcwb [28])
);

DFFPOSX1 _12198_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf88),
    .D(_0_[29]),
    .Q(\datapath.regcwb [29])
);

DFFPOSX1 _12199_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf87),
    .D(_0_[30]),
    .Q(\datapath.regcwb [30])
);

DFFPOSX1 _12200_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf86),
    .D(_0_[31]),
    .Q(\datapath.regcwb [31])
);

DFFPOSX1 _12201_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf85),
    .D(\datapath._52_ ),
    .Q(\datapath.regwbtrap )
);

DFFPOSX1 _12202_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf84),
    .D(\datapath.excpt_cause [0]),
    .Q(\datapath.csr.csr_mcause [0])
);

DFFPOSX1 _12203_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf83),
    .D(\datapath.excpt_cause [1]),
    .Q(\datapath.csr.csr_mcause [1])
);

DFFPOSX1 _12204_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf82),
    .D(\datapath.excpt_cause [2]),
    .Q(\datapath.csr.csr_mcause [2])
);

DFFPOSX1 _12205_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf81),
    .D(\datapath.excpt_cause [3]),
    .Q(\datapath.csr.csr_mcause [3])
);

DFFPOSX1 _12206_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf80),
    .D(\datapath._51_ ),
    .Q(\datapath.regmret )
);

DFFPOSX1 _12207_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf79),
    .D(\datapath._50_ ),
    .Q(\datapath.regcsrtrap )
);

DFFPOSX1 _12208_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf78),
    .D(\datapath._49_ [0]),
    .Q(\datapath.wbinstr [0])
);

DFFPOSX1 _12209_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf77),
    .D(\datapath._49_ [1]),
    .Q(\datapath.wbinstr [1])
);

DFFPOSX1 _12210_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf76),
    .D(\datapath._49_ [2]),
    .Q(\datapath.wbinstr [2])
);

DFFPOSX1 _12211_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf75),
    .D(\datapath._49_ [3]),
    .Q(\datapath.wbinstr [3])
);

DFFPOSX1 _12212_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf74),
    .D(\datapath._49_ [4]),
    .Q(\datapath.wbinstr [4])
);

DFFPOSX1 _12213_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf73),
    .D(\datapath._49_ [5]),
    .Q(\datapath.wbinstr [5])
);

DFFPOSX1 _12214_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf72),
    .D(\datapath._49_ [6]),
    .Q(\datapath.wbinstr [6])
);

DFFPOSX1 _12215_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf71),
    .D(\datapath._49_ [7]),
    .Q(\datapath.wbinstr [7])
);

DFFPOSX1 _12216_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf70),
    .D(\datapath._49_ [8]),
    .Q(\datapath.wbinstr [8])
);

DFFPOSX1 _12217_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf69),
    .D(\datapath._49_ [9]),
    .Q(\datapath.wbinstr [9])
);

DFFPOSX1 _12218_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf68),
    .D(\datapath._49_ [10]),
    .Q(\datapath.wbinstr [10])
);

DFFPOSX1 _12219_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf67),
    .D(\datapath._49_ [11]),
    .Q(\datapath.wbinstr [11])
);

DFFPOSX1 _12220_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf66),
    .D(\datapath._49_ [12]),
    .Q(\datapath.wbinstr [12])
);

DFFPOSX1 _12221_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf65),
    .D(\datapath._49_ [13]),
    .Q(\datapath.wbinstr [13])
);

DFFPOSX1 _12222_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf64),
    .D(\datapath._49_ [14]),
    .Q(\datapath.wbinstr [14])
);

DFFPOSX1 _12223_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf63),
    .D(\datapath.mempc_4 [0]),
    .Q(\datapath.wbpc_4 [0])
);

DFFPOSX1 _12224_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf62),
    .D(\datapath.mempc_4 [1]),
    .Q(\datapath.wbpc_4 [1])
);

DFFPOSX1 _12225_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf61),
    .D(\datapath.mempc_4 [2]),
    .Q(\datapath.wbpc_4 [2])
);

DFFPOSX1 _12226_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf60),
    .D(\datapath.mempc_4 [3]),
    .Q(\datapath.wbpc_4 [3])
);

DFFPOSX1 _12227_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf59),
    .D(\datapath.mempc_4 [4]),
    .Q(\datapath.wbpc_4 [4])
);

DFFPOSX1 _12228_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf58),
    .D(\datapath.mempc_4 [5]),
    .Q(\datapath.wbpc_4 [5])
);

DFFPOSX1 _12229_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf57),
    .D(\datapath.mempc_4 [6]),
    .Q(\datapath.wbpc_4 [6])
);

DFFPOSX1 _12230_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf56),
    .D(\datapath.mempc_4 [7]),
    .Q(\datapath.wbpc_4 [7])
);

DFFPOSX1 _12231_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf55),
    .D(\datapath.mempc_4 [8]),
    .Q(\datapath.wbpc_4 [8])
);

DFFPOSX1 _12232_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf54),
    .D(\datapath.mempc_4 [9]),
    .Q(\datapath.wbpc_4 [9])
);

DFFPOSX1 _12233_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf53),
    .D(\datapath.mempc_4 [10]),
    .Q(\datapath.wbpc_4 [10])
);

DFFPOSX1 _12234_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf52),
    .D(\datapath.mempc_4 [11]),
    .Q(\datapath.wbpc_4 [11])
);

DFFPOSX1 _12235_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf51),
    .D(\datapath.mempc_4 [12]),
    .Q(\datapath.wbpc_4 [12])
);

DFFPOSX1 _12236_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf50),
    .D(\datapath.mempc_4 [13]),
    .Q(\datapath.wbpc_4 [13])
);

DFFPOSX1 _12237_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf49),
    .D(\datapath.mempc_4 [14]),
    .Q(\datapath.wbpc_4 [14])
);

DFFPOSX1 _12238_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf48),
    .D(\datapath.mempc_4 [15]),
    .Q(\datapath.wbpc_4 [15])
);

DFFPOSX1 _12239_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf47),
    .D(\datapath.mempc_4 [16]),
    .Q(\datapath.wbpc_4 [16])
);

DFFPOSX1 _12240_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf46),
    .D(\datapath.mempc_4 [17]),
    .Q(\datapath.wbpc_4 [17])
);

DFFPOSX1 _12241_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf45),
    .D(\datapath.mempc_4 [18]),
    .Q(\datapath.wbpc_4 [18])
);

DFFPOSX1 _12242_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf44),
    .D(\datapath.mempc_4 [19]),
    .Q(\datapath.wbpc_4 [19])
);

DFFPOSX1 _12243_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf43),
    .D(\datapath.mempc_4 [20]),
    .Q(\datapath.wbpc_4 [20])
);

DFFPOSX1 _12244_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf42),
    .D(\datapath.mempc_4 [21]),
    .Q(\datapath.wbpc_4 [21])
);

DFFPOSX1 _12245_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf41),
    .D(\datapath.mempc_4 [22]),
    .Q(\datapath.wbpc_4 [22])
);

DFFPOSX1 _12246_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf40),
    .D(\datapath.mempc_4 [23]),
    .Q(\datapath.wbpc_4 [23])
);

DFFPOSX1 _12247_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf39),
    .D(\datapath.mempc_4 [24]),
    .Q(\datapath.wbpc_4 [24])
);

DFFPOSX1 _12248_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf38),
    .D(\datapath.mempc_4 [25]),
    .Q(\datapath.wbpc_4 [25])
);

DFFPOSX1 _12249_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf37),
    .D(\datapath.mempc_4 [26]),
    .Q(\datapath.wbpc_4 [26])
);

DFFPOSX1 _12250_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf36),
    .D(\datapath.mempc_4 [27]),
    .Q(\datapath.wbpc_4 [27])
);

DFFPOSX1 _12251_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf35),
    .D(\datapath.mempc_4 [28]),
    .Q(\datapath.wbpc_4 [28])
);

DFFPOSX1 _12252_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf34),
    .D(\datapath.mempc_4 [29]),
    .Q(\datapath.wbpc_4 [29])
);

DFFPOSX1 _12253_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf33),
    .D(\datapath.mempc_4 [30]),
    .Q(\datapath.wbpc_4 [30])
);

DFFPOSX1 _12254_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf32),
    .D(\datapath.mempc_4 [31]),
    .Q(\datapath.wbpc_4 [31])
);

DFFPOSX1 _12255_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf31),
    .D(\datapath.mempc [2]),
    .Q(\datapath.csr.csr_mepc [2])
);

DFFPOSX1 _12256_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf30),
    .D(\datapath.mempc [3]),
    .Q(\datapath.csr.csr_mepc [3])
);

DFFPOSX1 _12257_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf29),
    .D(\datapath.mempc [4]),
    .Q(\datapath.csr.csr_mepc [4])
);

DFFPOSX1 _12258_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf28),
    .D(\datapath.mempc [5]),
    .Q(\datapath.csr.csr_mepc [5])
);

DFFPOSX1 _12259_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf27),
    .D(\datapath.mempc [6]),
    .Q(\datapath.csr.csr_mepc [6])
);

DFFPOSX1 _12260_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf26),
    .D(\datapath.mempc [7]),
    .Q(\datapath.csr.csr_mepc [7])
);

DFFPOSX1 _12261_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf25),
    .D(\datapath.mempc [8]),
    .Q(\datapath.csr.csr_mepc [8])
);

DFFPOSX1 _12262_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf24),
    .D(\datapath.mempc [9]),
    .Q(\datapath.csr.csr_mepc [9])
);

DFFPOSX1 _12263_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf23),
    .D(\datapath.mempc [10]),
    .Q(\datapath.csr.csr_mepc [10])
);

DFFPOSX1 _12264_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf22),
    .D(\datapath.mempc [11]),
    .Q(\datapath.csr.csr_mepc [11])
);

DFFPOSX1 _12265_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf21),
    .D(\datapath.mempc [12]),
    .Q(\datapath.csr.csr_mepc [12])
);

DFFPOSX1 _12266_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf20),
    .D(\datapath.mempc [13]),
    .Q(\datapath.csr.csr_mepc [13])
);

DFFPOSX1 _12267_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf19),
    .D(\datapath.mempc [14]),
    .Q(\datapath.csr.csr_mepc [14])
);

DFFPOSX1 _12268_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf18),
    .D(\datapath.mempc [15]),
    .Q(\datapath.csr.csr_mepc [15])
);

DFFPOSX1 _12269_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf17),
    .D(\datapath.mempc [16]),
    .Q(\datapath.csr.csr_mepc [16])
);

DFFPOSX1 _12270_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf16),
    .D(\datapath.mempc [17]),
    .Q(\datapath.csr.csr_mepc [17])
);

DFFPOSX1 _12271_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf15),
    .D(\datapath.mempc [18]),
    .Q(\datapath.csr.csr_mepc [18])
);

DFFPOSX1 _12272_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf14),
    .D(\datapath.mempc [19]),
    .Q(\datapath.csr.csr_mepc [19])
);

DFFPOSX1 _12273_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf13),
    .D(\datapath.mempc [20]),
    .Q(\datapath.csr.csr_mepc [20])
);

DFFPOSX1 _12274_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf12),
    .D(\datapath.mempc [21]),
    .Q(\datapath.csr.csr_mepc [21])
);

DFFPOSX1 _12275_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf11),
    .D(\datapath.mempc [22]),
    .Q(\datapath.csr.csr_mepc [22])
);

DFFPOSX1 _12276_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf10),
    .D(\datapath.mempc [23]),
    .Q(\datapath.csr.csr_mepc [23])
);

DFFPOSX1 _12277_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf9),
    .D(\datapath.mempc [24]),
    .Q(\datapath.csr.csr_mepc [24])
);

DFFPOSX1 _12278_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf8),
    .D(\datapath.mempc [25]),
    .Q(\datapath.csr.csr_mepc [25])
);

DFFPOSX1 _12279_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf7),
    .D(\datapath.mempc [26]),
    .Q(\datapath.csr.csr_mepc [26])
);

DFFPOSX1 _12280_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf6),
    .D(\datapath.mempc [27]),
    .Q(\datapath.csr.csr_mepc [27])
);

DFFPOSX1 _12281_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf5),
    .D(\datapath.mempc [28]),
    .Q(\datapath.csr.csr_mepc [28])
);

DFFPOSX1 _12282_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf4),
    .D(\datapath.mempc [29]),
    .Q(\datapath.csr.csr_mepc [29])
);

DFFPOSX1 _12283_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf3),
    .D(\datapath.mempc [30]),
    .Q(\datapath.csr.csr_mepc [30])
);

DFFPOSX1 _12284_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf2),
    .D(\datapath.mempc [31]),
    .Q(\datapath.csr.csr_mepc [31])
);

\$_DLATCH_P_  _12285_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[0]),
    .E(_251_),
    .Q(\datapath.rs2bypass [0])
);

\$_DLATCH_P_  _12286_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[1]),
    .E(_251_),
    .Q(\datapath.rs2bypass [1])
);

\$_DLATCH_P_  _12287_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[2]),
    .E(_251_),
    .Q(\datapath.rs2bypass [2])
);

\$_DLATCH_P_  _12288_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[3]),
    .E(_251_),
    .Q(\datapath.rs2bypass [3])
);

\$_DLATCH_P_  _12289_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[4]),
    .E(_251_),
    .Q(\datapath.rs2bypass [4])
);

\$_DLATCH_P_  _12290_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[5]),
    .E(_251_),
    .Q(\datapath.rs2bypass [5])
);

\$_DLATCH_P_  _12291_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[6]),
    .E(_251_),
    .Q(\datapath.rs2bypass [6])
);

\$_DLATCH_P_  _12292_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[7]),
    .E(_251_),
    .Q(\datapath.rs2bypass [7])
);

\$_DLATCH_P_  _12293_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[8]),
    .E(_251_),
    .Q(\datapath.rs2bypass [8])
);

\$_DLATCH_P_  _12294_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[9]),
    .E(_251_),
    .Q(\datapath.rs2bypass [9])
);

\$_DLATCH_P_  _12295_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[10]),
    .E(_251_),
    .Q(\datapath.rs2bypass [10])
);

\$_DLATCH_P_  _12296_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[11]),
    .E(_251_),
    .Q(\datapath.rs2bypass [11])
);

\$_DLATCH_P_  _12297_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[12]),
    .E(_251_),
    .Q(\datapath.rs2bypass [12])
);

\$_DLATCH_P_  _12298_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[13]),
    .E(_251_),
    .Q(\datapath.rs2bypass [13])
);

\$_DLATCH_P_  _12299_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[14]),
    .E(_251_),
    .Q(\datapath.rs2bypass [14])
);

\$_DLATCH_P_  _12300_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[15]),
    .E(_251_),
    .Q(\datapath.rs2bypass [15])
);

\$_DLATCH_P_  _12301_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[16]),
    .E(_251_),
    .Q(\datapath.rs2bypass [16])
);

\$_DLATCH_P_  _12302_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[17]),
    .E(_251_),
    .Q(\datapath.rs2bypass [17])
);

\$_DLATCH_P_  _12303_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[18]),
    .E(_251_),
    .Q(\datapath.rs2bypass [18])
);

\$_DLATCH_P_  _12304_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[19]),
    .E(_251_),
    .Q(\datapath.rs2bypass [19])
);

\$_DLATCH_P_  _12305_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[20]),
    .E(_251_),
    .Q(\datapath.rs2bypass [20])
);

\$_DLATCH_P_  _12306_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[21]),
    .E(_251_),
    .Q(\datapath.rs2bypass [21])
);

\$_DLATCH_P_  _12307_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[22]),
    .E(_251_),
    .Q(\datapath.rs2bypass [22])
);

\$_DLATCH_P_  _12308_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[23]),
    .E(_251_),
    .Q(\datapath.rs2bypass [23])
);

\$_DLATCH_P_  _12309_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[24]),
    .E(_251_),
    .Q(\datapath.rs2bypass [24])
);

\$_DLATCH_P_  _12310_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[25]),
    .E(_251_),
    .Q(\datapath.rs2bypass [25])
);

\$_DLATCH_P_  _12311_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[26]),
    .E(_251_),
    .Q(\datapath.rs2bypass [26])
);

\$_DLATCH_P_  _12312_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[27]),
    .E(_251_),
    .Q(\datapath.rs2bypass [27])
);

\$_DLATCH_P_  _12313_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[28]),
    .E(_251_),
    .Q(\datapath.rs2bypass [28])
);

\$_DLATCH_P_  _12314_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[29]),
    .E(_251_),
    .Q(\datapath.rs2bypass [29])
);

\$_DLATCH_P_  _12315_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[30]),
    .E(_251_),
    .Q(\datapath.rs2bypass [30])
);

\$_DLATCH_P_  _12316_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_250_[31]),
    .E(_251_),
    .Q(\datapath.rs2bypass [31])
);

\$_DLATCH_P_  _12317_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[0]),
    .E(_252_),
    .Q(\datapath.bbypass [0])
);

\$_DLATCH_P_  _12318_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[1]),
    .E(_252_),
    .Q(\datapath.bbypass [1])
);

\$_DLATCH_P_  _12319_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[2]),
    .E(_252_),
    .Q(\datapath.bbypass [2])
);

\$_DLATCH_P_  _12320_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[3]),
    .E(_252_),
    .Q(\datapath.bbypass [3])
);

\$_DLATCH_P_  _12321_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[4]),
    .E(_252_),
    .Q(\datapath.bbypass [4])
);

\$_DLATCH_P_  _12322_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[5]),
    .E(_252_),
    .Q(\datapath.bbypass [5])
);

\$_DLATCH_P_  _12323_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[6]),
    .E(_252_),
    .Q(\datapath.bbypass [6])
);

\$_DLATCH_P_  _12324_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[7]),
    .E(_252_),
    .Q(\datapath.bbypass [7])
);

\$_DLATCH_P_  _12325_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[8]),
    .E(_252_),
    .Q(\datapath.bbypass [8])
);

\$_DLATCH_P_  _12326_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[9]),
    .E(_252_),
    .Q(\datapath.bbypass [9])
);

\$_DLATCH_P_  _12327_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[10]),
    .E(_252_),
    .Q(\datapath.bbypass [10])
);

\$_DLATCH_P_  _12328_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[11]),
    .E(_252_),
    .Q(\datapath.bbypass [11])
);

\$_DLATCH_P_  _12329_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[12]),
    .E(_252_),
    .Q(\datapath.bbypass [12])
);

\$_DLATCH_P_  _12330_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[13]),
    .E(_252_),
    .Q(\datapath.bbypass [13])
);

\$_DLATCH_P_  _12331_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[14]),
    .E(_252_),
    .Q(\datapath.bbypass [14])
);

\$_DLATCH_P_  _12332_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[15]),
    .E(_252_),
    .Q(\datapath.bbypass [15])
);

\$_DLATCH_P_  _12333_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[16]),
    .E(_252_),
    .Q(\datapath.bbypass [16])
);

\$_DLATCH_P_  _12334_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[17]),
    .E(_252_),
    .Q(\datapath.bbypass [17])
);

\$_DLATCH_P_  _12335_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[18]),
    .E(_252_),
    .Q(\datapath.bbypass [18])
);

\$_DLATCH_P_  _12336_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[19]),
    .E(_252_),
    .Q(\datapath.bbypass [19])
);

\$_DLATCH_P_  _12337_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[20]),
    .E(_252_),
    .Q(\datapath.bbypass [20])
);

\$_DLATCH_P_  _12338_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[21]),
    .E(_252_),
    .Q(\datapath.bbypass [21])
);

\$_DLATCH_P_  _12339_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[22]),
    .E(_252_),
    .Q(\datapath.bbypass [22])
);

\$_DLATCH_P_  _12340_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[23]),
    .E(_252_),
    .Q(\datapath.bbypass [23])
);

\$_DLATCH_P_  _12341_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[24]),
    .E(_252_),
    .Q(\datapath.bbypass [24])
);

\$_DLATCH_P_  _12342_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[25]),
    .E(_252_),
    .Q(\datapath.bbypass [25])
);

\$_DLATCH_P_  _12343_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[26]),
    .E(_252_),
    .Q(\datapath.bbypass [26])
);

\$_DLATCH_P_  _12344_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[27]),
    .E(_252_),
    .Q(\datapath.bbypass [27])
);

\$_DLATCH_P_  _12345_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[28]),
    .E(_252_),
    .Q(\datapath.bbypass [28])
);

\$_DLATCH_P_  _12346_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[29]),
    .E(_252_),
    .Q(\datapath.bbypass [29])
);

\$_DLATCH_P_  _12347_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[30]),
    .E(_252_),
    .Q(\datapath.bbypass [30])
);

\$_DLATCH_P_  _12348_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_249_[31]),
    .E(_252_),
    .Q(\datapath.bbypass [31])
);

\$_DLATCH_P_  _12349_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[0]),
    .E(_253_),
    .Q(\datapath.abypass [0])
);

\$_DLATCH_P_  _12350_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[1]),
    .E(_253_),
    .Q(\datapath.abypass [1])
);

\$_DLATCH_P_  _12351_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[2]),
    .E(_253_),
    .Q(\datapath.abypass [2])
);

\$_DLATCH_P_  _12352_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[3]),
    .E(_253_),
    .Q(\datapath.abypass [3])
);

\$_DLATCH_P_  _12353_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[4]),
    .E(_253_),
    .Q(\datapath.abypass [4])
);

\$_DLATCH_P_  _12354_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[5]),
    .E(_253_),
    .Q(\datapath.abypass [5])
);

\$_DLATCH_P_  _12355_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[6]),
    .E(_253_),
    .Q(\datapath.abypass [6])
);

\$_DLATCH_P_  _12356_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[7]),
    .E(_253_),
    .Q(\datapath.abypass [7])
);

\$_DLATCH_P_  _12357_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[8]),
    .E(_253_),
    .Q(\datapath.abypass [8])
);

\$_DLATCH_P_  _12358_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[9]),
    .E(_253_),
    .Q(\datapath.abypass [9])
);

\$_DLATCH_P_  _12359_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[10]),
    .E(_253_),
    .Q(\datapath.abypass [10])
);

\$_DLATCH_P_  _12360_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[11]),
    .E(_253_),
    .Q(\datapath.abypass [11])
);

\$_DLATCH_P_  _12361_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[12]),
    .E(_253_),
    .Q(\datapath.abypass [12])
);

\$_DLATCH_P_  _12362_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[13]),
    .E(_253_),
    .Q(\datapath.abypass [13])
);

\$_DLATCH_P_  _12363_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[14]),
    .E(_253_),
    .Q(\datapath.abypass [14])
);

\$_DLATCH_P_  _12364_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[15]),
    .E(_253_),
    .Q(\datapath.abypass [15])
);

\$_DLATCH_P_  _12365_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[16]),
    .E(_253_),
    .Q(\datapath.abypass [16])
);

\$_DLATCH_P_  _12366_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[17]),
    .E(_253_),
    .Q(\datapath.abypass [17])
);

\$_DLATCH_P_  _12367_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[18]),
    .E(_253_),
    .Q(\datapath.abypass [18])
);

\$_DLATCH_P_  _12368_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[19]),
    .E(_253_),
    .Q(\datapath.abypass [19])
);

\$_DLATCH_P_  _12369_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[20]),
    .E(_253_),
    .Q(\datapath.abypass [20])
);

\$_DLATCH_P_  _12370_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[21]),
    .E(_253_),
    .Q(\datapath.abypass [21])
);

\$_DLATCH_P_  _12371_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[22]),
    .E(_253_),
    .Q(\datapath.abypass [22])
);

\$_DLATCH_P_  _12372_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[23]),
    .E(_253_),
    .Q(\datapath.abypass [23])
);

\$_DLATCH_P_  _12373_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[24]),
    .E(_253_),
    .Q(\datapath.abypass [24])
);

\$_DLATCH_P_  _12374_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[25]),
    .E(_253_),
    .Q(\datapath.abypass [25])
);

\$_DLATCH_P_  _12375_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[26]),
    .E(_253_),
    .Q(\datapath.abypass [26])
);

\$_DLATCH_P_  _12376_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[27]),
    .E(_253_),
    .Q(\datapath.abypass [27])
);

\$_DLATCH_P_  _12377_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[28]),
    .E(_253_),
    .Q(\datapath.abypass [28])
);

\$_DLATCH_P_  _12378_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[29]),
    .E(_253_),
    .Q(\datapath.abypass [29])
);

\$_DLATCH_P_  _12379_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[30]),
    .E(_253_),
    .Q(\datapath.abypass [30])
);

\$_DLATCH_P_  _12380_ (
    .gnd(gnd),
    .vdd(vdd),
    .D(_248_[31]),
    .E(_253_),
    .Q(\datapath.abypass [31])
);

NAND2X1 _12381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [31]),
    .B(\datapath.alu.b [31]),
    .Y(_1620_)
);

INVX2 _12382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1620_),
    .Y(_1630_)
);

INVX2 _12383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [31]),
    .Y(_1641_)
);

INVX2 _12384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [31]),
    .Y(_1652_)
);

NAND2X1 _12385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1641_),
    .B(_1652_),
    .Y(_1663_)
);

INVX2 _12386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1663_),
    .Y(_1674_)
);

NAND2X1 _12387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [23]),
    .B(\datapath.alu.b [23]),
    .Y(_1684_)
);

INVX4 _12388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [23]),
    .Y(_1695_)
);

INVX2 _12389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [23]),
    .Y(_1706_)
);

NAND2X1 _12390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1695_),
    .B(_1706_),
    .Y(_1717_)
);

NAND2X1 _12391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1684_),
    .B(_1717_),
    .Y(_1727_)
);

INVX4 _12392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [22]),
    .Y(_1738_)
);

INVX2 _12393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [22]),
    .Y(_1749_)
);

NAND2X1 _12394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1738_),
    .B(_1749_),
    .Y(_1760_)
);

NAND2X1 _12395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [22]),
    .B(\datapath.alu.b [22]),
    .Y(_1770_)
);

NAND2X1 _12396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1770_),
    .B(_1760_),
    .Y(_1781_)
);

NAND2X1 _12397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1727_),
    .B(_1781_),
    .Y(_1792_)
);

NAND2X1 _12398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [21]),
    .B(\datapath.alu.b [21]),
    .Y(_1802_)
);

INVX2 _12399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1802_),
    .Y(_1813_)
);

NOR2X1 _12400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [21]),
    .B(\datapath.alu.b [21]),
    .Y(_1824_)
);

INVX2 _12401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [20]),
    .Y(_1835_)
);

INVX1 _12402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [20]),
    .Y(_1846_)
);

NAND2X1 _12403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1835_),
    .B(_1846_),
    .Y(_1856_)
);

NAND2X1 _12404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [20]),
    .B(\datapath.alu.b [20]),
    .Y(_1867_)
);

NAND2X1 _12405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1867_),
    .B(_1856_),
    .Y(_1878_)
);

OAI21X1 _12406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1813_),
    .B(_1824_),
    .C(_1878_),
    .Y(_1889_)
);

NOR2X1 _12407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1792_),
    .B(_1889_),
    .Y(_1899_)
);

INVX4 _12408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [19]),
    .Y(_1910_)
);

INVX1 _12409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [19]),
    .Y(_1921_)
);

NOR2X1 _12410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1910_),
    .B(_1921_),
    .Y(_1932_)
);

NOR2X1 _12411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [19]),
    .B(\datapath.alu.b [19]),
    .Y(_1942_)
);

NOR2X1 _12412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [18]),
    .B(\datapath.alu.b [18]),
    .Y(_1953_)
);

INVX4 _12413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [18]),
    .Y(_1964_)
);

INVX2 _12414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [18]),
    .Y(_1974_)
);

NOR2X1 _12415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1964_),
    .B(_1974_),
    .Y(_1985_)
);

OAI22X1 _12416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1932_),
    .B(_1942_),
    .C(_1953_),
    .D(_1985_),
    .Y(_1996_)
);

NAND2X1 _12417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [17]),
    .B(\datapath.alu.b [17]),
    .Y(_2007_)
);

INVX2 _12418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [17]),
    .Y(_2017_)
);

INVX1 _12419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [17]),
    .Y(_2028_)
);

NAND2X1 _12420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2017_),
    .B(_2028_),
    .Y(_2039_)
);

NAND2X1 _12421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2007_),
    .B(_2039_),
    .Y(_2050_)
);

NOR2X1 _12422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [16]),
    .B(\datapath.alu.b [16]),
    .Y(_2060_)
);

INVX4 _12423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [16]),
    .Y(_2071_)
);

INVX2 _12424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [16]),
    .Y(_2082_)
);

NOR2X1 _12425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2071_),
    .B(_2082_),
    .Y(_2092_)
);

OAI21X1 _12426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2060_),
    .B(_2092_),
    .C(_2050_),
    .Y(_2103_)
);

NOR2X1 _12427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1996_),
    .B(_2103_),
    .Y(_2114_)
);

NAND2X1 _12428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2114_),
    .B(_1899_),
    .Y(_2124_)
);

INVX1 _12429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [30]),
    .Y(_2135_)
);

INVX1 _12430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [30]),
    .Y(_2146_)
);

NAND2X1 _12431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2135_),
    .B(_2146_),
    .Y(_2157_)
);

NAND2X1 _12432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [30]),
    .B(\datapath.alu.b [30]),
    .Y(_2168_)
);

NAND2X1 _12433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2168_),
    .B(_2157_),
    .Y(_2178_)
);

OAI21X1 _12434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1674_),
    .B(_1630_),
    .C(_2178_),
    .Y(_2189_)
);

NAND2X1 _12435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [29]),
    .B(\datapath.alu.b [29]),
    .Y(_2200_)
);

INVX1 _12436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2200_),
    .Y(_2210_)
);

INVX2 _12437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [29]),
    .Y(_2221_)
);

INVX1 _12438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [29]),
    .Y(_2232_)
);

NAND2X1 _12439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2221_),
    .B(_2232_),
    .Y(_2243_)
);

INVX2 _12440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2243_),
    .Y(_2253_)
);

INVX2 _12441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [28]),
    .Y(_2264_)
);

INVX1 _12442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [28]),
    .Y(_2274_)
);

NAND2X1 _12443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2264_),
    .B(_2274_),
    .Y(_2285_)
);

NAND2X1 _12444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [28]),
    .B(\datapath.alu.b [28]),
    .Y(_2296_)
);

NAND2X1 _12445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2296_),
    .B(_2285_),
    .Y(_2307_)
);

OAI21X1 _12446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2253_),
    .B(_2210_),
    .C(_2307_),
    .Y(_2317_)
);

NOR2X1 _12447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2189_),
    .B(_2317_),
    .Y(_2328_)
);

NAND2X1 _12448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [27]),
    .B(\datapath.alu.b [27]),
    .Y(_2339_)
);

INVX2 _12449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [27]),
    .Y(_2349_)
);

INVX2 _12450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [27]),
    .Y(_2360_)
);

NAND2X1 _12451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2349_),
    .B(_2360_),
    .Y(_2371_)
);

NAND2X1 _12452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2339_),
    .B(_2371_),
    .Y(_2381_)
);

INVX2 _12453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [26]),
    .Y(_2392_)
);

INVX1 _12454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [26]),
    .Y(_2403_)
);

NAND2X1 _12455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2392_),
    .B(_2403_),
    .Y(_2413_)
);

NAND2X1 _12456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [26]),
    .B(\datapath.alu.b [26]),
    .Y(_2424_)
);

NAND2X1 _12457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2424_),
    .B(_2413_),
    .Y(_2430_)
);

NAND2X1 _12458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2381_),
    .B(_2430_),
    .Y(_2431_)
);

NAND2X1 _12459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [25]),
    .B(\datapath.alu.b [25]),
    .Y(_2432_)
);

INVX2 _12460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [25]),
    .Y(_2433_)
);

INVX1 _12461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [25]),
    .Y(_2434_)
);

NAND2X1 _12462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2433_),
    .B(_2434_),
    .Y(_2435_)
);

NAND2X1 _12463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2432_),
    .B(_2435_),
    .Y(_2436_)
);

NOR2X1 _12464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [24]),
    .B(\datapath.alu.b [24]),
    .Y(_2437_)
);

NAND2X1 _12465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [24]),
    .B(\datapath.alu.b [24]),
    .Y(_2438_)
);

INVX2 _12466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2438_),
    .Y(_2439_)
);

OAI21X1 _12467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_2439_),
    .C(_2436_),
    .Y(_2440_)
);

NOR2X1 _12468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2431_),
    .B(_2440_),
    .Y(_2441_)
);

NAND2X1 _12469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2441_),
    .B(_2328_),
    .Y(_2442_)
);

NOR2X1 _12470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2124_),
    .B(_2442_),
    .Y(_2443_)
);

NAND2X1 _12471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [15]),
    .B(\datapath.alu.b [15]),
    .Y(_2444_)
);

INVX2 _12472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [15]),
    .Y(_2445_)
);

INVX2 _12473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [15]),
    .Y(_2446_)
);

NAND2X1 _12474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2445_),
    .B(_2446_),
    .Y(_2447_)
);

NAND2X1 _12475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2444_),
    .B(_2447_),
    .Y(_2448_)
);

XNOR2X1 _12476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [14]),
    .B(\datapath.alu.b [14]),
    .Y(_2449_)
);

NAND2X1 _12477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2449_),
    .B(_2448_),
    .Y(_2450_)
);

INVX4 _12478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [12]),
    .Y(_2451_)
);

INVX4 _12479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [13]),
    .Y(_2452_)
);

AOI22X1 _12480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2451_),
    .B(\datapath.alu.b [12]),
    .C(_2452_),
    .D(\datapath.alu.b [13]),
    .Y(_2453_)
);

INVX2 _12481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [13]),
    .Y(_2454_)
);

NAND2X1 _12482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [13]),
    .B(_2454_),
    .Y(_2455_)
);

INVX1 _12483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [12]),
    .Y(_2456_)
);

NAND2X1 _12484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [12]),
    .B(_2456_),
    .Y(_2457_)
);

NAND3X1 _12485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2455_),
    .B(_2457_),
    .C(_2453_),
    .Y(_2458_)
);

NOR2X1 _12486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2458_),
    .B(_2450_),
    .Y(_2459_)
);

NAND2X1 _12487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [11]),
    .B(\datapath.alu.b [11]),
    .Y(_2460_)
);

INVX2 _12488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [11]),
    .Y(_2461_)
);

INVX2 _12489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [11]),
    .Y(_2462_)
);

NAND2X1 _12490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2461_),
    .B(_2462_),
    .Y(_2463_)
);

NAND2X1 _12491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2460_),
    .B(_2463_),
    .Y(_2464_)
);

XNOR2X1 _12492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [10]),
    .B(\datapath.alu.b [10]),
    .Y(_2465_)
);

NAND2X1 _12493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465_),
    .B(_2464_),
    .Y(_2466_)
);

XNOR2X1 _12494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [9]),
    .B(\datapath.alu.b [9]),
    .Y(_2467_)
);

XNOR2X1 _12495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [8]),
    .B(\datapath.alu.b [8]),
    .Y(_2468_)
);

NAND2X1 _12496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2467_),
    .B(_2468_),
    .Y(_2469_)
);

NOR2X1 _12497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2469_),
    .B(_2466_),
    .Y(_2470_)
);

NAND2X1 _12498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2459_),
    .B(_2470_),
    .Y(_2471_)
);

XNOR2X1 _12499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [7]),
    .B(\datapath.alu.b [7]),
    .Y(_2472_)
);

XNOR2X1 _12500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [6]),
    .B(\datapath.alu.b [6]),
    .Y(_2473_)
);

NAND2X1 _12501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2472_),
    .B(_2473_),
    .Y(_2474_)
);

INVX2 _12502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [4]),
    .Y(_2475_)
);

INVX4 _12503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [5]),
    .Y(_2476_)
);

AOI22X1 _12504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2475_),
    .B(\datapath.alu.b_4_bF$buf4 ),
    .C(_2476_),
    .D(\datapath.alu.b [5]),
    .Y(_2477_)
);

INVX2 _12505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [5]),
    .Y(_2478_)
);

NAND2X1 _12506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [5]),
    .B(_2478_),
    .Y(_2479_)
);

INVX8 _12507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_4_bF$buf3 ),
    .Y(_2480_)
);

NAND2X1 _12508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [4]),
    .B(_2480__bF$buf5),
    .Y(_2481_)
);

NAND3X1 _12509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2479_),
    .B(_2481_),
    .C(_2477_),
    .Y(_2482_)
);

NOR2X1 _12510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2474_),
    .B(_2482_),
    .Y(_2483_)
);

NAND2X1 _12511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf6 ),
    .B(\datapath.alu.a [3]),
    .Y(_2484_)
);

INVX1 _12512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2484_),
    .Y(_2485_)
);

NOR2X1 _12513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf5 ),
    .B(\datapath.alu.a [3]),
    .Y(_2486_)
);

XNOR2X1 _12514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf7 ),
    .B(\datapath.alu.a [2]),
    .Y(_2487_)
);

OAI21X1 _12515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2485_),
    .B(_2486_),
    .C(_2487_),
    .Y(_2488_)
);

INVX8 _12516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf6 ),
    .Y(_2489_)
);

NAND2X1 _12517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [1]),
    .B(_2489__bF$buf7),
    .Y(_2490_)
);

INVX4 _12518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf10 ),
    .Y(_2491_)
);

NAND2X1 _12519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [0]),
    .B(_2491_),
    .Y(_2492_)
);

NOR2X1 _12520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [1]),
    .B(_2489__bF$buf6),
    .Y(_2493_)
);

OAI21X1 _12521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2493_),
    .B(_2492_),
    .C(_2490_),
    .Y(_2494_)
);

INVX8 _12522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf6 ),
    .Y(_2495_)
);

NOR2X1 _12523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [2]),
    .B(_2495__bF$buf6),
    .Y(_2496_)
);

INVX8 _12524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf4 ),
    .Y(_2497_)
);

NOR2X1 _12525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [3]),
    .B(_2497__bF$buf6),
    .Y(_2498_)
);

NAND2X1 _12526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [3]),
    .B(_2497__bF$buf5),
    .Y(_2499_)
);

AOI21X1 _12527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2499_),
    .B(_2496_),
    .C(_2498_),
    .Y(_2500_)
);

OAI21X1 _12528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2488_),
    .B(_2494_),
    .C(_2500_),
    .Y(_2501_)
);

INVX4 _12529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [7]),
    .Y(_2502_)
);

INVX2 _12530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [7]),
    .Y(_2503_)
);

INVX4 _12531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [6]),
    .Y(_2504_)
);

NAND2X1 _12532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [6]),
    .B(_2504_),
    .Y(_2505_)
);

OAI21X1 _12533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [7]),
    .B(_2503_),
    .C(_2505_),
    .Y(_2506_)
);

OAI21X1 _12534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2502_),
    .B(\datapath.alu.b [7]),
    .C(_2506_),
    .Y(_2507_)
);

NOR2X1 _12535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [5]),
    .B(_2476_),
    .Y(_2508_)
);

OR2X2 _12536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2477_),
    .B(_2508_),
    .Y(_2509_)
);

OAI21X1 _12537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2509_),
    .B(_2474_),
    .C(_2507_),
    .Y(_2510_)
);

AOI21X1 _12538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2483_),
    .B(_2501_),
    .C(_2510_),
    .Y(_2511_)
);

INVX2 _12539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [9]),
    .Y(_2512_)
);

NOR2X1 _12540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [9]),
    .B(_2512_),
    .Y(_2513_)
);

NAND2X1 _12541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [9]),
    .B(_2512_),
    .Y(_2514_)
);

INVX2 _12542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [8]),
    .Y(_2515_)
);

NOR2X1 _12543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [8]),
    .B(_2515_),
    .Y(_2516_)
);

OAI21X1 _12544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2513_),
    .B(_2516_),
    .C(_2514_),
    .Y(_2517_)
);

INVX2 _12545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [10]),
    .Y(_2518_)
);

NOR2X1 _12546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [10]),
    .B(_2518_),
    .Y(_2519_)
);

NOR2X1 _12547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [11]),
    .B(_2462_),
    .Y(_2520_)
);

NOR2X1 _12548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [11]),
    .B(_2461_),
    .Y(_2521_)
);

INVX1 _12549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2521_),
    .Y(_2522_)
);

AOI21X1 _12550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519_),
    .B(_2522_),
    .C(_2520_),
    .Y(_2523_)
);

OAI21X1 _12551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2466_),
    .B(_2517_),
    .C(_2523_),
    .Y(_2524_)
);

NAND2X1 _12552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [13]),
    .B(_2452_),
    .Y(_2525_)
);

INVX1 _12553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2525_),
    .Y(_2526_)
);

NAND2X1 _12554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [12]),
    .B(_2451_),
    .Y(_2527_)
);

INVX1 _12555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2527_),
    .Y(_2528_)
);

OAI21X1 _12556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2528_),
    .B(_2526_),
    .C(_2455_),
    .Y(_2529_)
);

INVX2 _12557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [14]),
    .Y(_2530_)
);

NAND2X1 _12558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [14]),
    .B(_2530_),
    .Y(_2531_)
);

INVX2 _12559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2531_),
    .Y(_2532_)
);

NOR2X1 _12560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [15]),
    .B(_2445_),
    .Y(_2533_)
);

INVX1 _12561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2533_),
    .Y(_2534_)
);

NOR2X1 _12562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [15]),
    .B(_2446_),
    .Y(_2535_)
);

OAI21X1 _12563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2532_),
    .B(_2535_),
    .C(_2534_),
    .Y(_2536_)
);

OAI21X1 _12564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2529_),
    .B(_2450_),
    .C(_2536_),
    .Y(_2537_)
);

AOI21X1 _12565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2459_),
    .B(_2524_),
    .C(_2537_),
    .Y(_2538_)
);

OAI21X1 _12566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2511_),
    .B(_2471_),
    .C(_2538_),
    .Y(_2539_)
);

NOR2X1 _12567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [17]),
    .B(_2028_),
    .Y(_2540_)
);

NOR2X1 _12568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [16]),
    .B(_2082_),
    .Y(_2541_)
);

NAND2X1 _12569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [17]),
    .B(_2028_),
    .Y(_2542_)
);

OAI21X1 _12570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2540_),
    .B(_2541_),
    .C(_2542_),
    .Y(_2543_)
);

NAND2X1 _12571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [19]),
    .B(_1910_),
    .Y(_2544_)
);

OAI21X1 _12572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [18]),
    .B(_1974_),
    .C(_2544_),
    .Y(_2545_)
);

OAI21X1 _12573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1910_),
    .B(\datapath.alu.b [19]),
    .C(_2545_),
    .Y(_2546_)
);

OAI21X1 _12574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1996_),
    .B(_2543_),
    .C(_2546_),
    .Y(_2547_)
);

INVX1 _12575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [21]),
    .Y(_2548_)
);

NOR2X1 _12576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [21]),
    .B(_2548_),
    .Y(_2549_)
);

NOR2X1 _12577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [20]),
    .B(_1846_),
    .Y(_2550_)
);

INVX2 _12578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [21]),
    .Y(_2551_)
);

NOR2X1 _12579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [21]),
    .B(_2551_),
    .Y(_2552_)
);

INVX1 _12580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2552_),
    .Y(_2553_)
);

OAI21X1 _12581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2549_),
    .B(_2550_),
    .C(_2553_),
    .Y(_2554_)
);

NOR2X1 _12582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [22]),
    .B(_1749_),
    .Y(_2555_)
);

NOR2X1 _12583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [23]),
    .B(_1706_),
    .Y(_2556_)
);

AOI21X1 _12584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2555_),
    .B(_1727_),
    .C(_2556_),
    .Y(_2557_)
);

OAI21X1 _12585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1792_),
    .B(_2554_),
    .C(_2557_),
    .Y(_2558_)
);

AOI21X1 _12586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2547_),
    .B(_1899_),
    .C(_2558_),
    .Y(_2559_)
);

NOR2X1 _12587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [25]),
    .B(_2434_),
    .Y(_2560_)
);

INVX1 _12588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [24]),
    .Y(_2561_)
);

NOR2X1 _12589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [24]),
    .B(_2561_),
    .Y(_2562_)
);

NAND2X1 _12590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [25]),
    .B(_2434_),
    .Y(_2563_)
);

OAI21X1 _12591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560_),
    .B(_2562_),
    .C(_2563_),
    .Y(_2564_)
);

NAND2X1 _12592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [27]),
    .B(_2360_),
    .Y(_2565_)
);

NOR2X1 _12593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [26]),
    .B(_2403_),
    .Y(_2566_)
);

NOR2X1 _12594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [27]),
    .B(_2360_),
    .Y(_2567_)
);

OAI21X1 _12595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2566_),
    .B(_2567_),
    .C(_2565_),
    .Y(_2568_)
);

OAI21X1 _12596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2431_),
    .B(_2564_),
    .C(_2568_),
    .Y(_2569_)
);

NAND2X1 _12597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [29]),
    .B(_2232_),
    .Y(_2570_)
);

NOR2X1 _12598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [29]),
    .B(_2232_),
    .Y(_2571_)
);

NOR2X1 _12599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [28]),
    .B(_2274_),
    .Y(_2572_)
);

OAI21X1 _12600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2571_),
    .B(_2572_),
    .C(_2570_),
    .Y(_2573_)
);

NAND2X1 _12601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1620_),
    .B(_1663_),
    .Y(_2574_)
);

NOR2X1 _12602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [31]),
    .B(_1652_),
    .Y(_2575_)
);

NOR2X1 _12603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [30]),
    .B(_2146_),
    .Y(_2576_)
);

AOI21X1 _12604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2576_),
    .B(_2574_),
    .C(_2575_),
    .Y(_2577_)
);

OAI21X1 _12605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2189_),
    .B(_2573_),
    .C(_2577_),
    .Y(_2578_)
);

AOI21X1 _12606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2328_),
    .B(_2569_),
    .C(_2578_),
    .Y(_2579_)
);

OAI21X1 _12607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2559_),
    .B(_2442_),
    .C(_2579_),
    .Y(_2580_)
);

AOI21X1 _12608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2443_),
    .B(_2539_),
    .C(_2580_),
    .Y(_2581_)
);

OAI21X1 _12609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1630_),
    .B(_1674_),
    .C(_2581_),
    .Y(_2582_)
);

AND2X2 _12610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1899_),
    .B(_2114_),
    .Y(_2583_)
);

AND2X2 _12611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2328_),
    .B(_2441_),
    .Y(_2584_)
);

NAND2X1 _12612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2583_),
    .B(_2584_),
    .Y(_2585_)
);

INVX2 _12613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [14]),
    .Y(_2586_)
);

NAND2X1 _12614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [14]),
    .B(_2586_),
    .Y(_2587_)
);

NAND2X1 _12615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2531_),
    .B(_2587_),
    .Y(_2588_)
);

AOI21X1 _12616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2444_),
    .B(_2447_),
    .C(_2588_),
    .Y(_2589_)
);

NAND2X1 _12617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2525_),
    .B(_2455_),
    .Y(_2590_)
);

NAND2X1 _12618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2527_),
    .B(_2457_),
    .Y(_2591_)
);

NOR2X1 _12619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2590_),
    .B(_2591_),
    .Y(_2592_)
);

NAND2X1 _12620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2589_),
    .B(_2592_),
    .Y(_2593_)
);

XOR2X1 _12621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [10]),
    .B(\datapath.alu.b [10]),
    .Y(_2594_)
);

AOI21X1 _12622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2460_),
    .B(_2463_),
    .C(_2594_),
    .Y(_2595_)
);

INVX2 _12623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [9]),
    .Y(_2596_)
);

NAND2X1 _12624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [9]),
    .B(_2596_),
    .Y(_2597_)
);

NAND2X1 _12625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2597_),
    .B(_2514_),
    .Y(_2598_)
);

INVX4 _12626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [8]),
    .Y(_2599_)
);

NAND2X1 _12627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [8]),
    .B(_2599_),
    .Y(_2600_)
);

NAND2X1 _12628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [8]),
    .B(_2515_),
    .Y(_2601_)
);

NAND2X1 _12629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2600_),
    .B(_2601_),
    .Y(_2602_)
);

NOR2X1 _12630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2598_),
    .B(_2602_),
    .Y(_2603_)
);

NAND2X1 _12631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2595_),
    .B(_2603_),
    .Y(_2604_)
);

NOR2X1 _12632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2604_),
    .B(_2593_),
    .Y(_2605_)
);

XOR2X1 _12633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf3 ),
    .B(\datapath.alu.a [3]),
    .Y(_2606_)
);

XOR2X1 _12634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf5 ),
    .B(\datapath.alu.a [2]),
    .Y(_2607_)
);

NOR2X1 _12635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2606_),
    .B(_2607_),
    .Y(_2608_)
);

XOR2X1 _12636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf5 ),
    .B(\datapath.alu.a [1]),
    .Y(_2609_)
);

NOR2X1 _12637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf9 ),
    .B(\datapath.alu.a [0]),
    .Y(_2610_)
);

NAND2X1 _12638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf8 ),
    .B(\datapath.alu.a [0]),
    .Y(_2611_)
);

INVX2 _12639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2611_),
    .Y(_2612_)
);

NOR2X1 _12640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2610_),
    .B(_2612_),
    .Y(_2613_)
);

NOR2X1 _12641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2609_),
    .B(_2613_),
    .Y(_2614_)
);

AND2X2 _12642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2614_),
    .B(_2608_),
    .Y(_2615_)
);

NAND3X1 _12643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2483_),
    .B(_2615_),
    .C(_2605_),
    .Y(_2616_)
);

NOR2X1 _12644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2616_),
    .B(_2585_),
    .Y(_2617_)
);

INVX1 _12645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.funsel [1]),
    .Y(_2618_)
);

NOR2X1 _12646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.funsel [0]),
    .B(_2618_),
    .Y(_2619_)
);

NOR2X1 _12647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.funsel [2]),
    .B(_2575_),
    .Y(_2620_)
);

NAND2X1 _12648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2619_),
    .B(_2620_),
    .Y(_2621_)
);

NOR2X1 _12649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2621_),
    .B(_2617_),
    .Y(_2622_)
);

NAND2X1 _12650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.funsel [0]),
    .B(\datapath.alu.funsel [1]),
    .Y(_2623_)
);

NOR2X1 _12651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.funsel [2]),
    .B(_2623_),
    .Y(_2624_)
);

OAI21X1 _12652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2585_),
    .B(_2616_),
    .C(_2624_),
    .Y(_2625_)
);

INVX2 _12653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [2]),
    .Y(_2626_)
);

NAND2X1 _12654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf7 ),
    .B(\datapath.alu.a [3]),
    .Y(_2627_)
);

OAI21X1 _12655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2626_),
    .B(\datapath.alu.b_0_bF$buf6 ),
    .C(_2627_),
    .Y(_2628_)
);

NOR2X1 _12656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf5),
    .B(_2628_),
    .Y(_2629_)
);

INVX2 _12657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [0]),
    .Y(_2630_)
);

NAND2X1 _12658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf5 ),
    .B(\datapath.alu.a [1]),
    .Y(_2631_)
);

OAI21X1 _12659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2630_),
    .B(\datapath.alu.b_0_bF$buf4 ),
    .C(_2631_),
    .Y(_2632_)
);

NOR2X1 _12660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf4 ),
    .B(_2632_),
    .Y(_2633_)
);

OAI21X1 _12661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2629_),
    .B(_2633_),
    .C(_2495__bF$buf5),
    .Y(_2634_)
);

NAND2X1 _12662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [6]),
    .B(_2491_),
    .Y(_2635_)
);

NAND2X1 _12663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf3 ),
    .B(\datapath.alu.a [7]),
    .Y(_2636_)
);

NAND3X1 _12664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf3 ),
    .B(_2636_),
    .C(_2635_),
    .Y(_2637_)
);

NAND2X1 _12665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf2 ),
    .B(\datapath.alu.a [5]),
    .Y(_2638_)
);

OAI21X1 _12666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2475_),
    .B(\datapath.alu.b_0_bF$buf1 ),
    .C(_2638_),
    .Y(_2639_)
);

OAI21X1 _12667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf2 ),
    .B(_2639_),
    .C(_2637_),
    .Y(_2640_)
);

NAND2X1 _12668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf4 ),
    .B(_2640_),
    .Y(_2641_)
);

NAND3X1 _12669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf4),
    .B(_2634_),
    .C(_2641_),
    .Y(_2642_)
);

NAND2X1 _12670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf0 ),
    .B(\datapath.alu.a [15]),
    .Y(_2643_)
);

OAI21X1 _12671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2530_),
    .B(\datapath.alu.b_0_bF$buf10 ),
    .C(_2643_),
    .Y(_2644_)
);

NAND2X1 _12672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf9 ),
    .B(\datapath.alu.a [13]),
    .Y(_2645_)
);

OAI21X1 _12673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2451_),
    .B(\datapath.alu.b_0_bF$buf8 ),
    .C(_2645_),
    .Y(_2646_)
);

MUX2X1 _12674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2646_),
    .B(_2644_),
    .S(_2489__bF$buf4),
    .Y(_2647_)
);

INVX2 _12675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [10]),
    .Y(_2648_)
);

NAND2X1 _12676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf7 ),
    .B(\datapath.alu.a [11]),
    .Y(_2649_)
);

OAI21X1 _12677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648_),
    .B(\datapath.alu.b_0_bF$buf6 ),
    .C(_2649_),
    .Y(_2650_)
);

NAND2X1 _12678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf5 ),
    .B(\datapath.alu.a [9]),
    .Y(_2651_)
);

OAI21X1 _12679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2599_),
    .B(\datapath.alu.b_0_bF$buf4 ),
    .C(_2651_),
    .Y(_2652_)
);

MUX2X1 _12680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2652_),
    .B(_2650_),
    .S(_2489__bF$buf3),
    .Y(_2653_)
);

MUX2X1 _12681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2653_),
    .B(_2647_),
    .S(_2495__bF$buf4),
    .Y(_2654_)
);

NAND2X1 _12682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf2 ),
    .B(_2654_),
    .Y(_2655_)
);

INVX1 _12683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.funsel [2]),
    .Y(_2656_)
);

NAND2X1 _12684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.funsel [0]),
    .B(_2618_),
    .Y(_2657_)
);

NOR2X1 _12685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2656_),
    .B(_2657_),
    .Y(_2658_)
);

NAND2X1 _12686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf4),
    .B(_2658_),
    .Y(_2659_)
);

AOI21X1 _12687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2655_),
    .B(_2642_),
    .C(_2659_),
    .Y(_2660_)
);

MUX2X1 _12688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [31]),
    .B(\datapath.alu.a [30]),
    .S(\datapath.alu.b_0_bF$buf3 ),
    .Y(_2661_)
);

MUX2X1 _12689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [29]),
    .B(\datapath.alu.a [28]),
    .S(\datapath.alu.b_0_bF$buf2 ),
    .Y(_2662_)
);

MUX2X1 _12690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2662_),
    .B(_2661_),
    .S(_2489__bF$buf2),
    .Y(_2663_)
);

MUX2X1 _12691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [27]),
    .B(\datapath.alu.a [26]),
    .S(\datapath.alu.b_0_bF$buf1 ),
    .Y(_2664_)
);

MUX2X1 _12692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [25]),
    .B(\datapath.alu.a [24]),
    .S(\datapath.alu.b_0_bF$buf0 ),
    .Y(_2665_)
);

MUX2X1 _12693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2665_),
    .B(_2664_),
    .S(_2489__bF$buf1),
    .Y(_2666_)
);

MUX2X1 _12694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2666_),
    .B(_2663_),
    .S(_2495__bF$buf3),
    .Y(_2667_)
);

MUX2X1 _12695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [23]),
    .B(\datapath.alu.a [22]),
    .S(\datapath.alu.b_0_bF$buf10 ),
    .Y(_2668_)
);

MUX2X1 _12696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [21]),
    .B(\datapath.alu.a [20]),
    .S(\datapath.alu.b_0_bF$buf9 ),
    .Y(_2669_)
);

MUX2X1 _12697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2669_),
    .B(_2668_),
    .S(_2489__bF$buf0),
    .Y(_2670_)
);

MUX2X1 _12698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [19]),
    .B(\datapath.alu.a [18]),
    .S(\datapath.alu.b_0_bF$buf8 ),
    .Y(_2671_)
);

MUX2X1 _12699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [17]),
    .B(\datapath.alu.a [16]),
    .S(\datapath.alu.b_0_bF$buf7 ),
    .Y(_2672_)
);

MUX2X1 _12700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2672_),
    .B(_2671_),
    .S(_2489__bF$buf7),
    .Y(_2673_)
);

MUX2X1 _12701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2673_),
    .B(_2670_),
    .S(_2495__bF$buf2),
    .Y(_2674_)
);

MUX2X1 _12702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2674_),
    .B(_2667_),
    .S(_2497__bF$buf3),
    .Y(_2675_)
);

INVX2 _12703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2658_),
    .Y(_2676_)
);

NOR2X1 _12704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf3),
    .B(_2676_),
    .Y(_2677_)
);

AND2X2 _12705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2675_),
    .B(_2677_),
    .Y(_2678_)
);

NOR2X1 _12706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.funsel [3]),
    .B(_2656_),
    .Y(_2679_)
);

NAND2X1 _12707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2619_),
    .B(_2679_),
    .Y(_2680_)
);

NOR2X1 _12708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2610_),
    .B(_2680__bF$buf3),
    .Y(_2681_)
);

NOR2X1 _12709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.funsel [1]),
    .B(\datapath.alu.funsel [2]),
    .Y(_2682_)
);

INVX2 _12710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2682_),
    .Y(_2683_)
);

INVX1 _12711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.funsel [0]),
    .Y(_2684_)
);

NAND2X1 _12712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.funsel [3]),
    .B(_2684_),
    .Y(_2685_)
);

INVX2 _12713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.funsel [3]),
    .Y(_2686_)
);

NOR2X1 _12714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.funsel [0]),
    .B(\datapath.alu.funsel [1]),
    .Y(_2687_)
);

NAND3X1 _12715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686_),
    .B(\datapath.alu.funsel [2]),
    .C(_2687_),
    .Y(_2688_)
);

OAI21X1 _12716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2683_),
    .B(_2685_),
    .C(_2688__bF$buf3),
    .Y(_2689_)
);

AND2X2 _12717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2689_),
    .B(_2613_),
    .Y(_2690_)
);

INVX1 _12718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2623_),
    .Y(_2691_)
);

NAND2X1 _12719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2691_),
    .B(_2679_),
    .Y(_2692_)
);

AND2X2 _12720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.funsel [3]),
    .B(\datapath.alu.funsel [2]),
    .Y(_2693_)
);

NAND2X1 _12721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2687_),
    .B(_2693_),
    .Y(_2694_)
);

OAI22X1 _12722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2630_),
    .B(_2694_),
    .C(_2692_),
    .D(_2611_),
    .Y(_2695_)
);

NOR3X1 _12723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2681_),
    .B(_2695_),
    .C(_2690_),
    .Y(_2696_)
);

OR2X2 _12724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2492_),
    .B(\datapath.alu.b_1_bF$buf1 ),
    .Y(_2697_)
);

NOR3X1 _12725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf1 ),
    .B(\datapath.alu.b_2_bF$buf3 ),
    .C(_2697_),
    .Y(_2698_)
);

NAND2X1 _12726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.funsel [0]),
    .B(_2686_),
    .Y(_2699_)
);

OR2X2 _12727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2683_),
    .B(_2699_),
    .Y(_2700_)
);

NOR2X1 _12728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_4_bF$buf2 ),
    .B(_2700_),
    .Y(_2701_)
);

NAND3X1 _12729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2682_),
    .B(_2699_),
    .C(_2685_),
    .Y(_2702_)
);

INVX8 _12730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2702_),
    .Y(_2703_)
);

AOI22X1 _12731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2613_),
    .B(_2703__bF$buf3),
    .C(_2698_),
    .D(_2701_),
    .Y(_2704_)
);

NAND2X1 _12732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.funsel [3]),
    .B(\datapath.alu.funsel [2]),
    .Y(_2705_)
);

NOR2X1 _12733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2623_),
    .B(_2705_),
    .Y(_2706_)
);

INVX8 _12734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2706__bF$buf3),
    .Y(_2707_)
);

NAND2X1 _12735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2693_),
    .B(_2619_),
    .Y(_2708_)
);

OAI21X1 _12736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2707_),
    .B(\datapath.alu.a [0]),
    .C(_2708__bF$buf3),
    .Y(_2709_)
);

NAND2X1 _12737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf6 ),
    .B(_2709_),
    .Y(_2710_)
);

NAND3X1 _12738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2704_),
    .B(_2710_),
    .C(_2696_),
    .Y(_2711_)
);

NOR3X1 _12739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2711_),
    .B(_2678_),
    .C(_2660_),
    .Y(_2712_)
);

OAI21X1 _12740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2581_),
    .B(_2625_),
    .C(_2712_),
    .Y(_2713_)
);

AOI21X1 _12741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2582_),
    .B(_2622_),
    .C(_2713_),
    .Y(_2714_)
);

INVX2 _12742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2714_),
    .Y(\datapath.alu.condtrue )
);

NAND2X1 _12743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.funsel [2]),
    .B(_2686_),
    .Y(_2715_)
);

NOR2X1 _12744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2657_),
    .B(_2715_),
    .Y(_2716_)
);

NOR2X1 _12745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2705_),
    .B(_2657_),
    .Y(_2717_)
);

NAND2X1 _12746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf5 ),
    .B(\datapath.alu.a [24]),
    .Y(_2718_)
);

OAI21X1 _12747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1695_),
    .B(\datapath.alu.b_0_bF$buf4 ),
    .C(_2718_),
    .Y(_2719_)
);

NAND2X1 _12748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf3 ),
    .B(\datapath.alu.a [22]),
    .Y(_2720_)
);

OAI21X1 _12749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551_),
    .B(\datapath.alu.b_0_bF$buf2 ),
    .C(_2720_),
    .Y(_2721_)
);

MUX2X1 _12750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2721_),
    .B(_2719_),
    .S(_2489__bF$buf6),
    .Y(_2722_)
);

MUX2X1 _12751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [20]),
    .B(\datapath.alu.a [19]),
    .S(\datapath.alu.b_0_bF$buf1 ),
    .Y(_2723_)
);

NAND2X1 _12752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf0 ),
    .B(_2723_),
    .Y(_2724_)
);

NAND2X1 _12753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf0 ),
    .B(\datapath.alu.a [18]),
    .Y(_2725_)
);

OAI21X1 _12754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2017_),
    .B(\datapath.alu.b_0_bF$buf10 ),
    .C(_2725_),
    .Y(_2726_)
);

OAI21X1 _12755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf6 ),
    .B(_2726_),
    .C(_2724_),
    .Y(_2727_)
);

MUX2X1 _12756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2727_),
    .B(_2722_),
    .S(_2495__bF$buf1),
    .Y(_2728_)
);

NAND2X1 _12757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf2),
    .B(_2728_),
    .Y(_2729_)
);

NAND2X1 _12758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf9 ),
    .B(\datapath.alu.a [28]),
    .Y(_2730_)
);

OAI21X1 _12759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2349_),
    .B(\datapath.alu.b_0_bF$buf8 ),
    .C(_2730_),
    .Y(_2731_)
);

NAND2X1 _12760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf7 ),
    .B(\datapath.alu.a [26]),
    .Y(_2732_)
);

OAI21X1 _12761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2433_),
    .B(\datapath.alu.b_0_bF$buf6 ),
    .C(_2732_),
    .Y(_2733_)
);

MUX2X1 _12762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2733_),
    .B(_2731_),
    .S(_2489__bF$buf5),
    .Y(_2734_)
);

NOR2X1 _12763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf2 ),
    .B(_2734_),
    .Y(_2735_)
);

NAND2X1 _12764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf5 ),
    .B(\datapath.alu.a [30]),
    .Y(_2736_)
);

OAI21X1 _12765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2221_),
    .B(\datapath.alu.b_0_bF$buf4 ),
    .C(_2736_),
    .Y(_2737_)
);

NAND2X1 _12766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf4),
    .B(_2737_),
    .Y(_2738_)
);

OAI21X1 _12767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf3),
    .B(_1641_),
    .C(_2738_),
    .Y(_2739_)
);

AOI21X1 _12768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf1 ),
    .B(_2739_),
    .C(_2735_),
    .Y(_2740_)
);

OAI21X1 _12769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2740_),
    .B(_2497__bF$buf1),
    .C(_2729_),
    .Y(_2741_)
);

NOR2X1 _12770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf3 ),
    .B(_1641_),
    .Y(_2742_)
);

MUX2X1 _12771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2737_),
    .B(_2742_),
    .S(_2489__bF$buf2),
    .Y(_2743_)
);

INVX1 _12772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2743_),
    .Y(_2744_)
);

AOI21X1 _12773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf0 ),
    .B(_2744_),
    .C(_2735_),
    .Y(_2745_)
);

OAI21X1 _12774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2745_),
    .B(_2497__bF$buf0),
    .C(_2729_),
    .Y(_2746_)
);

AOI22X1 _12775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2741_),
    .B(_2717_),
    .C(_2716_),
    .D(_2746_),
    .Y(_2747_)
);

INVX1 _12776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2747_),
    .Y(_2748_)
);

NAND2X1 _12777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf2 ),
    .B(\datapath.alu.a [8]),
    .Y(_2749_)
);

OAI21X1 _12778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2502_),
    .B(\datapath.alu.b_0_bF$buf1 ),
    .C(_2749_),
    .Y(_2750_)
);

NAND2X1 _12779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf0 ),
    .B(\datapath.alu.a [6]),
    .Y(_2751_)
);

OAI21X1 _12780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2476_),
    .B(\datapath.alu.b_0_bF$buf10 ),
    .C(_2751_),
    .Y(_2752_)
);

MUX2X1 _12781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2752_),
    .B(_2750_),
    .S(_2489__bF$buf1),
    .Y(_2753_)
);

INVX2 _12782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [1]),
    .Y(_2754_)
);

NAND2X1 _12783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf9 ),
    .B(\datapath.alu.a [2]),
    .Y(_2755_)
);

OAI21X1 _12784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2754_),
    .B(\datapath.alu.b_0_bF$buf8 ),
    .C(_2755_),
    .Y(_2756_)
);

NOR2X1 _12785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf5 ),
    .B(_2756_),
    .Y(_2757_)
);

INVX2 _12786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [3]),
    .Y(_2758_)
);

NAND2X1 _12787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf7 ),
    .B(\datapath.alu.a [4]),
    .Y(_2759_)
);

OAI21X1 _12788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2758_),
    .B(\datapath.alu.b_0_bF$buf6 ),
    .C(_2759_),
    .Y(_2760_)
);

OAI21X1 _12789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2760_),
    .B(_2489__bF$buf0),
    .C(_2495__bF$buf0),
    .Y(_2761_)
);

OAI22X1 _12790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2761_),
    .B(_2757_),
    .C(_2753_),
    .D(_2495__bF$buf6),
    .Y(_2762_)
);

MUX2X1 _12791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [16]),
    .B(\datapath.alu.a [15]),
    .S(\datapath.alu.b_0_bF$buf5 ),
    .Y(_2763_)
);

NAND2X1 _12792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf4 ),
    .B(_2763_),
    .Y(_2764_)
);

NAND2X1 _12793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf4 ),
    .B(\datapath.alu.a [14]),
    .Y(_2765_)
);

OAI21X1 _12794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2452_),
    .B(\datapath.alu.b_0_bF$buf3 ),
    .C(_2765_),
    .Y(_2766_)
);

OAI21X1 _12795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf3 ),
    .B(_2766_),
    .C(_2764_),
    .Y(_2767_)
);

INVX1 _12796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2767_),
    .Y(_2768_)
);

NAND2X1 _12797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf2 ),
    .B(\datapath.alu.a [12]),
    .Y(_2769_)
);

OAI21X1 _12798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2461_),
    .B(\datapath.alu.b_0_bF$buf1 ),
    .C(_2769_),
    .Y(_2770_)
);

NAND2X1 _12799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf0 ),
    .B(\datapath.alu.a [10]),
    .Y(_2771_)
);

OAI21X1 _12800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2596_),
    .B(\datapath.alu.b_0_bF$buf10 ),
    .C(_2771_),
    .Y(_2772_)
);

MUX2X1 _12801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2772_),
    .B(_2770_),
    .S(_2489__bF$buf7),
    .Y(_2773_)
);

NAND2X1 _12802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495__bF$buf5),
    .B(_2773_),
    .Y(_2774_)
);

OAI21X1 _12803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2768_),
    .B(_2495__bF$buf4),
    .C(_2774_),
    .Y(_2775_)
);

AOI21X1 _12804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf0 ),
    .B(_2775_),
    .C(_2659_),
    .Y(_2776_)
);

OAI21X1 _12805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf6 ),
    .B(_2762_),
    .C(_2776_),
    .Y(_2777_)
);

NOR2X1 _12806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf2 ),
    .B(_2754_),
    .Y(_2778_)
);

OAI21X1 _12807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2778_),
    .B(_2493_),
    .C(_2611_),
    .Y(_2779_)
);

XNOR2X1 _12808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf1 ),
    .B(\datapath.alu.a [1]),
    .Y(_2780_)
);

NAND2X1 _12809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2612_),
    .B(_2780_),
    .Y(_2781_)
);

AOI21X1 _12810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2781_),
    .B(_2779_),
    .C(_2702_),
    .Y(_2782_)
);

INVX1 _12811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2782_),
    .Y(_2783_)
);

OAI21X1 _12812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2692_),
    .B(_2489__bF$buf6),
    .C(_2694_),
    .Y(_2784_)
);

NAND2X1 _12813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf5),
    .B(_2754_),
    .Y(_2785_)
);

NAND2X1 _12814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf0 ),
    .B(\datapath.alu.a [1]),
    .Y(_2786_)
);

INVX1 _12815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2786_),
    .Y(_2787_)
);

OAI21X1 _12816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2688__bF$buf2),
    .B(_2787_),
    .C(_2680__bF$buf2),
    .Y(_2788_)
);

AOI22X1 _12817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2785_),
    .B(_2788_),
    .C(_2784_),
    .D(\datapath.alu.a [1]),
    .Y(_2789_)
);

AND2X2 _12818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2789_),
    .B(_2783_),
    .Y(_2790_)
);

OAI21X1 _12819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2754_),
    .B(\datapath.alu.b_0_bF$buf9 ),
    .C(_2611_),
    .Y(_2791_)
);

NAND2X1 _12820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf4),
    .B(_2791_),
    .Y(_2792_)
);

OR2X2 _12821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2792_),
    .B(\datapath.alu.b_2_bF$buf7 ),
    .Y(_2793_)
);

NOR2X1 _12822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf5 ),
    .B(_2793_),
    .Y(_2794_)
);

NAND2X1 _12823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf8 ),
    .B(_2630_),
    .Y(_2795_)
);

NOR2X1 _12824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2795_),
    .B(_2780_),
    .Y(_2796_)
);

NOR2X1 _12825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [0]),
    .B(_2491_),
    .Y(_2797_)
);

OR2X2 _12826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2683_),
    .B(_2685_),
    .Y(_2798_)
);

INVX8 _12827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2798_),
    .Y(_2799_)
);

OAI21X1 _12828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2609_),
    .B(_2797_),
    .C(_2799__bF$buf3),
    .Y(_2800_)
);

NAND2X1 _12829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.funsel [1]),
    .B(_2684_),
    .Y(_2801_)
);

NOR2X1 _12830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2705_),
    .B(_2801_),
    .Y(_2802_)
);

AOI22X1 _12831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2493_),
    .B(_2706__bF$buf2),
    .C(_2802_),
    .D(\datapath.alu.b_1_bF$buf6 ),
    .Y(_2803_)
);

OAI21X1 _12832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2800_),
    .B(_2796_),
    .C(_2803_),
    .Y(_2804_)
);

AOI21X1 _12833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2701_),
    .B(_2794_),
    .C(_2804_),
    .Y(_2805_)
);

NAND3X1 _12834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2805_),
    .B(_2790_),
    .C(_2777_),
    .Y(_2806_)
);

AOI21X1 _12835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_4_bF$buf1 ),
    .B(_2748_),
    .C(_2806_),
    .Y(_2807_)
);

INVX2 _12836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2807_),
    .Y(\datapath.alu.c [1])
);

INVX4 _12837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2716_),
    .Y(_2808_)
);

INVX4 _12838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2717_),
    .Y(_2809_)
);

INVX4 _12839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [24]),
    .Y(_2810_)
);

NAND2X1 _12840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf7 ),
    .B(\datapath.alu.a [25]),
    .Y(_2811_)
);

OAI21X1 _12841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2810_),
    .B(\datapath.alu.b_0_bF$buf6 ),
    .C(_2811_),
    .Y(_2812_)
);

NAND2X1 _12842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf5 ),
    .B(\datapath.alu.a [23]),
    .Y(_2813_)
);

OAI21X1 _12843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1738_),
    .B(\datapath.alu.b_0_bF$buf4 ),
    .C(_2813_),
    .Y(_2814_)
);

MUX2X1 _12844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2814_),
    .B(_2812_),
    .S(_2489__bF$buf3),
    .Y(_2815_)
);

NAND2X1 _12845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf3 ),
    .B(\datapath.alu.a [21]),
    .Y(_2816_)
);

OAI21X1 _12846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1835_),
    .B(\datapath.alu.b_0_bF$buf2 ),
    .C(_2816_),
    .Y(_2817_)
);

NAND2X1 _12847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf1 ),
    .B(\datapath.alu.a [19]),
    .Y(_2818_)
);

OAI21X1 _12848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1964_),
    .B(\datapath.alu.b_0_bF$buf0 ),
    .C(_2818_),
    .Y(_2819_)
);

MUX2X1 _12849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2819_),
    .B(_2817_),
    .S(_2489__bF$buf2),
    .Y(_2820_)
);

MUX2X1 _12850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2820_),
    .B(_2815_),
    .S(_2495__bF$buf3),
    .Y(_2821_)
);

NAND2X1 _12851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf10 ),
    .B(\datapath.alu.a [29]),
    .Y(_2822_)
);

OAI21X1 _12852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2264_),
    .B(\datapath.alu.b_0_bF$buf9 ),
    .C(_2822_),
    .Y(_2823_)
);

NAND2X1 _12853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf8 ),
    .B(\datapath.alu.a [27]),
    .Y(_2824_)
);

OAI21X1 _12854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2392_),
    .B(\datapath.alu.b_0_bF$buf7 ),
    .C(_2824_),
    .Y(_2825_)
);

MUX2X1 _12855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825_),
    .B(_2823_),
    .S(_2489__bF$buf1),
    .Y(_2826_)
);

NAND2X1 _12856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf6 ),
    .B(\datapath.alu.a [31]),
    .Y(_2827_)
);

OAI21X1 _12857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2135_),
    .B(\datapath.alu.b_0_bF$buf5 ),
    .C(_2827_),
    .Y(_2828_)
);

MUX2X1 _12858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2828_),
    .B(\datapath.alu.a [31]),
    .S(_2489__bF$buf0),
    .Y(_2829_)
);

MUX2X1 _12859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2826_),
    .B(_2829_),
    .S(_2495__bF$buf2),
    .Y(_2830_)
);

MUX2X1 _12860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2821_),
    .B(_2830_),
    .S(_2497__bF$buf6),
    .Y(_2831_)
);

NAND2X1 _12861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf7),
    .B(_2828_),
    .Y(_2832_)
);

MUX2X1 _12862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2826_),
    .B(_2832_),
    .S(_2495__bF$buf1),
    .Y(_2833_)
);

MUX2X1 _12863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2821_),
    .B(_2833_),
    .S(_2497__bF$buf5),
    .Y(_2834_)
);

OAI22X1 _12864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2831_),
    .B(_2809_),
    .C(_2808_),
    .D(_2834_),
    .Y(_2835_)
);

NAND2X1 _12865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf4 ),
    .B(\datapath.alu.a [17]),
    .Y(_2836_)
);

OAI21X1 _12866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2071_),
    .B(\datapath.alu.b_0_bF$buf3 ),
    .C(_2836_),
    .Y(_2837_)
);

NOR2X1 _12867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf6),
    .B(_2837_),
    .Y(_2838_)
);

NOR2X1 _12868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf5 ),
    .B(_2644_),
    .Y(_2839_)
);

OAI21X1 _12869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2838_),
    .B(_2839_),
    .C(\datapath.alu.b_2_bF$buf6 ),
    .Y(_2840_)
);

NOR2X1 _12870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf5),
    .B(_2646_),
    .Y(_2841_)
);

NOR2X1 _12871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf4 ),
    .B(_2650_),
    .Y(_2842_)
);

OAI21X1 _12872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2841_),
    .B(_2842_),
    .C(_2495__bF$buf0),
    .Y(_2843_)
);

AOI21X1 _12873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2843_),
    .B(_2840_),
    .C(_2497__bF$buf4),
    .Y(_2844_)
);

OAI21X1 _12874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2504_),
    .B(\datapath.alu.b_0_bF$buf2 ),
    .C(_2636_),
    .Y(_2845_)
);

MUX2X1 _12875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2652_),
    .B(_2845_),
    .S(\datapath.alu.b_1_bF$buf3 ),
    .Y(_2846_)
);

MUX2X1 _12876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2639_),
    .B(_2628_),
    .S(\datapath.alu.b_1_bF$buf2 ),
    .Y(_2847_)
);

MUX2X1 _12877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2847_),
    .B(_2846_),
    .S(_2495__bF$buf6),
    .Y(_2848_)
);

OAI21X1 _12878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2848_),
    .B(\datapath.alu.b_3_bF$buf4 ),
    .C(_2658_),
    .Y(_2849_)
);

OAI21X1 _12879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2630_),
    .B(\datapath.alu.b_0_bF$buf1 ),
    .C(\datapath.alu.b_1_bF$buf1 ),
    .Y(_2850_)
);

OAI21X1 _12880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2626_),
    .B(\datapath.alu.b_0_bF$buf0 ),
    .C(_2631_),
    .Y(_2851_)
);

OAI21X1 _12881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2851_),
    .B(\datapath.alu.b_1_bF$buf0 ),
    .C(_2850_),
    .Y(_2852_)
);

NOR2X1 _12882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf5 ),
    .B(_2852_),
    .Y(_2853_)
);

NOR2X1 _12883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf3 ),
    .B(_2700_),
    .Y(_2854_)
);

AOI21X1 _12884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2854_),
    .B(_2853_),
    .C(_2677_),
    .Y(_2855_)
);

OAI21X1 _12885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2849_),
    .B(_2844_),
    .C(_2855_),
    .Y(_2856_)
);

OAI21X1 _12886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2835_),
    .B(_2480__bF$buf2),
    .C(_2856_),
    .Y(_2857_)
);

NAND2X1 _12887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf6 ),
    .B(_2754_),
    .Y(_2858_)
);

AOI21X1 _12888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2858_),
    .B(_2795_),
    .C(_2778_),
    .Y(_2859_)
);

AOI21X1 _12889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2607_),
    .B(_2859_),
    .C(_2798_),
    .Y(_2860_)
);

OAI21X1 _12890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2607_),
    .B(_2859_),
    .C(_2860_),
    .Y(_2861_)
);

OAI21X1 _12891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2780_),
    .B(_2611_),
    .C(_2786_),
    .Y(_2862_)
);

OAI21X1 _12892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2862_),
    .B(_2607_),
    .C(_2703__bF$buf2),
    .Y(_2863_)
);

AOI21X1 _12893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2607_),
    .B(_2862_),
    .C(_2863_),
    .Y(_2864_)
);

NOR2X1 _12894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2623_),
    .B(_2715_),
    .Y(_2865_)
);

NAND2X1 _12895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf4 ),
    .B(\datapath.alu.a [2]),
    .Y(_2866_)
);

INVX2 _12896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2866_),
    .Y(_2867_)
);

AOI22X1 _12897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2496_),
    .B(_2706__bF$buf1),
    .C(_2865__bF$buf3),
    .D(_2867_),
    .Y(_2868_)
);

INVX8 _12898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2694_),
    .Y(_2869_)
);

AOI22X1 _12899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf3 ),
    .B(_2802_),
    .C(_2869__bF$buf3),
    .D(\datapath.alu.a [2]),
    .Y(_2870_)
);

OAI21X1 _12900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2688__bF$buf1),
    .B(_2867_),
    .C(_2680__bF$buf1),
    .Y(_2871_)
);

OAI21X1 _12901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf2 ),
    .B(\datapath.alu.a [2]),
    .C(_2871_),
    .Y(_2872_)
);

NAND3X1 _12902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2868_),
    .B(_2870_),
    .C(_2872_),
    .Y(_2873_)
);

NOR2X1 _12903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2864_),
    .B(_2873_),
    .Y(_2874_)
);

AND2X2 _12904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2874_),
    .B(_2861_),
    .Y(_2875_)
);

NAND2X1 _12905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2875_),
    .B(_2857_),
    .Y(\datapath.alu.c [2])
);

XNOR2X1 _12906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf2 ),
    .B(\datapath.alu.a [3]),
    .Y(_2876_)
);

NAND2X1 _12907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [2]),
    .B(_2495__bF$buf5),
    .Y(_2877_)
);

OAI21X1 _12908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2859_),
    .B(_2496_),
    .C(_2877_),
    .Y(_2878_)
);

OAI21X1 _12909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2878_),
    .B(_2876_),
    .C(_2799__bF$buf2),
    .Y(_2879_)
);

AOI21X1 _12910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2876_),
    .B(_2878_),
    .C(_2879_),
    .Y(_2880_)
);

AOI21X1 _12911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2607_),
    .B(_2862_),
    .C(_2867_),
    .Y(_2881_)
);

OAI21X1 _12912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2881_),
    .B(_2876_),
    .C(_2703__bF$buf1),
    .Y(_2882_)
);

AOI21X1 _12913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2876_),
    .B(_2881_),
    .C(_2882_),
    .Y(_2883_)
);

INVX4 _12914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2701_),
    .Y(_2884_)
);

OAI21X1 _12915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2758_),
    .B(\datapath.alu.b_0_bF$buf10 ),
    .C(_2755_),
    .Y(_2885_)
);

MUX2X1 _12916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2885_),
    .B(_2791_),
    .S(_2489__bF$buf4),
    .Y(_2886_)
);

INVX1 _12917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2886_),
    .Y(_2887_)
);

NAND3X1 _12918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf3),
    .B(_2495__bF$buf4),
    .C(_2887_),
    .Y(_2888_)
);

NAND2X1 _12919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2498_),
    .B(_2706__bF$buf0),
    .Y(_2889_)
);

OAI21X1 _12920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2758_),
    .B(_2694_),
    .C(_2889_),
    .Y(_2890_)
);

OAI22X1 _12921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2876_),
    .B(_2688__bF$buf0),
    .C(_2708__bF$buf2),
    .D(_2497__bF$buf2),
    .Y(_2891_)
);

OAI22X1 _12922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2692_),
    .B(_2484_),
    .C(_2680__bF$buf0),
    .D(_2486_),
    .Y(_2892_)
);

NOR3X1 _12923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2891_),
    .B(_2890_),
    .C(_2892_),
    .Y(_2893_)
);

OAI21X1 _12924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884_),
    .B(_2888_),
    .C(_2893_),
    .Y(_2894_)
);

NOR3X1 _12925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2880_),
    .B(_2894_),
    .C(_2883_),
    .Y(_2895_)
);

MUX2X1 _12926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2752_),
    .B(_2760_),
    .S(\datapath.alu.b_1_bF$buf5 ),
    .Y(_2896_)
);

MUX2X1 _12927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2772_),
    .B(_2750_),
    .S(\datapath.alu.b_1_bF$buf4 ),
    .Y(_2897_)
);

MUX2X1 _12928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2897_),
    .B(_2896_),
    .S(\datapath.alu.b_2_bF$buf1 ),
    .Y(_2898_)
);

NAND2X1 _12929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf9 ),
    .B(\datapath.alu.a [16]),
    .Y(_2899_)
);

OAI21X1 _12930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2445_),
    .B(\datapath.alu.b_0_bF$buf8 ),
    .C(_2899_),
    .Y(_2900_)
);

MUX2X1 _12931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2900_),
    .B(_2726_),
    .S(_2489__bF$buf3),
    .Y(_2901_)
);

MUX2X1 _12932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2770_),
    .B(_2766_),
    .S(_2489__bF$buf2),
    .Y(_2902_)
);

MUX2X1 _12933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2902_),
    .B(_2901_),
    .S(_2495__bF$buf3),
    .Y(_2903_)
);

MUX2X1 _12934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2903_),
    .B(_2898_),
    .S(\datapath.alu.b_3_bF$buf1 ),
    .Y(_2904_)
);

MUX2X1 _12935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2733_),
    .B(_2719_),
    .S(\datapath.alu.b_1_bF$buf3 ),
    .Y(_2905_)
);

NAND2X1 _12936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf7 ),
    .B(\datapath.alu.a [20]),
    .Y(_2906_)
);

OAI21X1 _12937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1910_),
    .B(\datapath.alu.b_0_bF$buf6 ),
    .C(_2906_),
    .Y(_2907_)
);

MUX2X1 _12938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2907_),
    .B(_2721_),
    .S(_2489__bF$buf1),
    .Y(_2908_)
);

MUX2X1 _12939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2908_),
    .B(_2905_),
    .S(_2495__bF$buf2),
    .Y(_2909_)
);

MUX2X1 _12940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2737_),
    .B(_2731_),
    .S(\datapath.alu.b_1_bF$buf2 ),
    .Y(_2910_)
);

NAND2X1 _12941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf0 ),
    .B(\datapath.alu.a [31]),
    .Y(_2911_)
);

OAI21X1 _12942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2910_),
    .B(\datapath.alu.b_2_bF$buf7 ),
    .C(_2911_),
    .Y(_2912_)
);

MUX2X1 _12943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2909_),
    .B(_2912_),
    .S(_2497__bF$buf1),
    .Y(_2913_)
);

MUX2X1 _12944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2904_),
    .B(_2913_),
    .S(_2480__bF$buf1),
    .Y(_2914_)
);

NAND2X1 _12945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [31]),
    .B(_2491_),
    .Y(_2915_)
);

NOR2X1 _12946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf1 ),
    .B(_2915_),
    .Y(_2916_)
);

NAND2X1 _12947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf6 ),
    .B(_2916_),
    .Y(_2917_)
);

OAI21X1 _12948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf5 ),
    .B(_2910_),
    .C(_2917_),
    .Y(_2918_)
);

MUX2X1 _12949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2918_),
    .B(_2909_),
    .S(\datapath.alu.b_3_bF$buf0 ),
    .Y(_2919_)
);

MUX2X1 _12950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2919_),
    .B(_2904_),
    .S(\datapath.alu.b_4_bF$buf0 ),
    .Y(_2920_)
);

AOI22X1 _12951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2717_),
    .B(_2914_),
    .C(_2920_),
    .D(_2716_),
    .Y(_2921_)
);

NAND2X1 _12952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2895_),
    .B(_2921_),
    .Y(\datapath.alu.c [3])
);

MUX2X1 _12953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2812_),
    .B(_2825_),
    .S(_2489__bF$buf0),
    .Y(_2922_)
);

NAND2X1 _12954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf4 ),
    .B(_2922_),
    .Y(_2923_)
);

MUX2X1 _12955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2817_),
    .B(_2814_),
    .S(_2489__bF$buf7),
    .Y(_2924_)
);

NAND2X1 _12956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495__bF$buf1),
    .B(_2924_),
    .Y(_2925_)
);

NAND3X1 _12957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf0),
    .B(_2923_),
    .C(_2925_),
    .Y(_2926_)
);

INVX1 _12958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2911_),
    .Y(_2927_)
);

MUX2X1 _12959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2823_),
    .B(_2828_),
    .S(_2489__bF$buf6),
    .Y(_2928_)
);

NOR2X1 _12960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf3 ),
    .B(_2928_),
    .Y(_2929_)
);

OAI21X1 _12961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2929_),
    .B(_2927_),
    .C(\datapath.alu.b_3_bF$buf6 ),
    .Y(_2930_)
);

AOI21X1 _12962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2926_),
    .B(_2930_),
    .C(_2809_),
    .Y(_2931_)
);

NAND2X1 _12963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf5 ),
    .B(_2929_),
    .Y(_2932_)
);

AOI21X1 _12964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2932_),
    .B(_2926_),
    .C(_2808_),
    .Y(_2933_)
);

OAI21X1 _12965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2931_),
    .B(_2933_),
    .C(\datapath.alu.b_4_bF$buf4 ),
    .Y(_2934_)
);

NOR2X1 _12966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [4]),
    .B(_2480__bF$buf0),
    .Y(_2935_)
);

NOR2X1 _12967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_4_bF$buf3 ),
    .B(_2475_),
    .Y(_2936_)
);

AOI21X1 _12968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2612_),
    .B(_2609_),
    .C(_2787_),
    .Y(_2937_)
);

NOR2X1 _12969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf2 ),
    .B(_2626_),
    .Y(_2938_)
);

OAI21X1 _12970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2496_),
    .B(_2938_),
    .C(_2606_),
    .Y(_2939_)
);

OAI21X1 _12971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2486_),
    .B(_2866_),
    .C(_2484_),
    .Y(_2940_)
);

INVX1 _12972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2940_),
    .Y(_2941_)
);

OAI21X1 _12973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2937_),
    .B(_2939_),
    .C(_2941_),
    .Y(_2942_)
);

OAI21X1 _12974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2935_),
    .B(_2936_),
    .C(_2942_),
    .Y(_2943_)
);

NOR2X1 _12975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2935_),
    .B(_2936_),
    .Y(_2944_)
);

NOR2X1 _12976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2876_),
    .B(_2487_),
    .Y(_2945_)
);

AOI21X1 _12977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2945_),
    .B(_2862_),
    .C(_2940_),
    .Y(_2946_)
);

AOI21X1 _12978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2944_),
    .B(_2946_),
    .C(_2702_),
    .Y(_2947_)
);

NAND2X1 _12979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2943_),
    .B(_2947_),
    .Y(_2948_)
);

NAND2X1 _12980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [10]),
    .B(_2491_),
    .Y(_2949_)
);

NAND3X1 _12981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf0 ),
    .B(_2649_),
    .C(_2949_),
    .Y(_2950_)
);

NAND2X1 _12982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [8]),
    .B(_2491_),
    .Y(_2951_)
);

NAND3X1 _12983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf5),
    .B(_2651_),
    .C(_2951_),
    .Y(_2952_)
);

AOI21X1 _12984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2950_),
    .B(_2952_),
    .C(_2495__bF$buf0),
    .Y(_2953_)
);

NAND2X1 _12985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [4]),
    .B(_2491_),
    .Y(_2954_)
);

NAND3X1 _12986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf4),
    .B(_2638_),
    .C(_2954_),
    .Y(_2955_)
);

AOI21X1 _12987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2637_),
    .B(_2955_),
    .C(\datapath.alu.b_2_bF$buf1 ),
    .Y(_2956_)
);

OAI21X1 _12988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2956_),
    .B(_2953_),
    .C(_2497__bF$buf6),
    .Y(_2957_)
);

MUX2X1 _12989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [15]),
    .B(\datapath.alu.a [14]),
    .S(\datapath.alu.b_0_bF$buf5 ),
    .Y(_2958_)
);

MUX2X1 _12990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [13]),
    .B(\datapath.alu.a [12]),
    .S(\datapath.alu.b_0_bF$buf4 ),
    .Y(_2959_)
);

MUX2X1 _12991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2959_),
    .B(_2958_),
    .S(_2489__bF$buf3),
    .Y(_2960_)
);

MUX2X1 _12992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2673_),
    .B(_2960_),
    .S(\datapath.alu.b_2_bF$buf0 ),
    .Y(_2961_)
);

AOI21X1 _12993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf4 ),
    .B(_2961_),
    .C(_2659_),
    .Y(_2962_)
);

MUX2X1 _12994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [1]),
    .B(\datapath.alu.a [2]),
    .S(\datapath.alu.b_0_bF$buf3 ),
    .Y(_2963_)
);

MUX2X1 _12995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [3]),
    .B(\datapath.alu.a [4]),
    .S(\datapath.alu.b_0_bF$buf2 ),
    .Y(_2964_)
);

MUX2X1 _12996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2964_),
    .B(_2963_),
    .S(_2489__bF$buf2),
    .Y(_2965_)
);

OAI21X1 _12997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2492_),
    .B(\datapath.alu.b_1_bF$buf6 ),
    .C(\datapath.alu.b_2_bF$buf7 ),
    .Y(_2966_)
);

OAI21X1 _12998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2965_),
    .B(\datapath.alu.b_2_bF$buf6 ),
    .C(_2966_),
    .Y(_2967_)
);

NOR2X1 _12999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf3 ),
    .B(_2967_),
    .Y(_2968_)
);

AOI22X1 _13000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2701_),
    .B(_2968_),
    .C(_2962_),
    .D(_2957_),
    .Y(_2969_)
);

AND2X2 _13001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2969_),
    .B(_2948_),
    .Y(_2970_)
);

NOR2X1 _13002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf2 ),
    .B(_2758_),
    .Y(_2971_)
);

AOI21X1 _13003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2938_),
    .B(_2876_),
    .C(_2971_),
    .Y(_2972_)
);

OAI21X1 _13004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2488_),
    .B(_2859_),
    .C(_2972_),
    .Y(_2973_)
);

NAND2X1 _13005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2944_),
    .B(_2973_),
    .Y(_2974_)
);

INVX1 _13006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2944_),
    .Y(_2975_)
);

OAI21X1 _13007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2493_),
    .B(_2797_),
    .C(_2490_),
    .Y(_2976_)
);

OAI21X1 _13008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2606_),
    .B(_2877_),
    .C(_2499_),
    .Y(_2977_)
);

AOI21X1 _13009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2976_),
    .B(_2608_),
    .C(_2977_),
    .Y(_2978_)
);

AOI21X1 _13010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2975_),
    .B(_2978_),
    .C(_2798_),
    .Y(_2979_)
);

NOR2X1 _13011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf5),
    .B(_2475_),
    .Y(_2980_)
);

AOI22X1 _13012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2935_),
    .B(_2706__bF$buf3),
    .C(_2865__bF$buf2),
    .D(_2980_),
    .Y(_2981_)
);

OAI21X1 _13013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2688__bF$buf3),
    .B(_2980_),
    .C(_2680__bF$buf3),
    .Y(_2982_)
);

OAI21X1 _13014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_4_bF$buf2 ),
    .B(\datapath.alu.a [4]),
    .C(_2982_),
    .Y(_2983_)
);

AOI22X1 _13015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_4_bF$buf1 ),
    .B(_2802_),
    .C(_2869__bF$buf2),
    .D(\datapath.alu.a [4]),
    .Y(_2984_)
);

NAND3X1 _13016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2981_),
    .B(_2984_),
    .C(_2983_),
    .Y(_2985_)
);

AOI21X1 _13017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2974_),
    .B(_2979_),
    .C(_2985_),
    .Y(_2986_)
);

NAND3X1 _13018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2986_),
    .B(_2934_),
    .C(_2970_),
    .Y(\datapath.alu.c [4])
);

XOR2X1 _13019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [5]),
    .B(\datapath.alu.b [5]),
    .Y(_2987_)
);

AOI21X1 _13020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2944_),
    .B(_2973_),
    .C(_2936_),
    .Y(_2988_)
);

AOI21X1 _13021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2987_),
    .B(_2988_),
    .C(_2798_),
    .Y(_2989_)
);

OAI21X1 _13022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2987_),
    .B(_2988_),
    .C(_2989_),
    .Y(_2990_)
);

MUX2X1 _13023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2734_),
    .B(_2722_),
    .S(\datapath.alu.b_2_bF$buf5 ),
    .Y(_2991_)
);

OAI21X1 _13024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf4 ),
    .B(\datapath.alu.b_1_bF$buf5 ),
    .C(\datapath.alu.a [31]),
    .Y(_2992_)
);

OAI21X1 _13025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2738_),
    .B(\datapath.alu.b_2_bF$buf3 ),
    .C(_2992_),
    .Y(_2993_)
);

MUX2X1 _13026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2991_),
    .B(_2993_),
    .S(_2497__bF$buf5),
    .Y(_2994_)
);

NOR2X1 _13027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf2 ),
    .B(_2743_),
    .Y(_2995_)
);

MUX2X1 _13028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2991_),
    .B(_2995_),
    .S(_2497__bF$buf4),
    .Y(_2996_)
);

OAI22X1 _13029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2994_),
    .B(_2809_),
    .C(_2808_),
    .D(_2996_),
    .Y(_2997_)
);

NOR2X1 _13030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2476_),
    .B(_2478_),
    .Y(_2998_)
);

OAI21X1 _13031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2688__bF$buf2),
    .B(_2998_),
    .C(_2680__bF$buf2),
    .Y(_2999_)
);

OAI21X1 _13032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [5]),
    .B(\datapath.alu.b [5]),
    .C(_2999_),
    .Y(_3000_)
);

NAND2X1 _13033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [5]),
    .B(_2476_),
    .Y(_3001_)
);

INVX1 _13034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2998_),
    .Y(_3002_)
);

OAI22X1 _13035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2692_),
    .B(_3002_),
    .C(_2707_),
    .D(_3001_),
    .Y(_3003_)
);

OAI22X1 _13036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2476_),
    .B(_2694_),
    .C(_2708__bF$buf1),
    .D(_2478_),
    .Y(_3004_)
);

NOR2X1 _13037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3004_),
    .B(_3003_),
    .Y(_3005_)
);

NAND2X1 _13038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3000_),
    .B(_3005_),
    .Y(_3006_)
);

AOI21X1 _13039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_4_bF$buf0 ),
    .B(_2997_),
    .C(_3006_),
    .Y(_3007_)
);

INVX1 _13040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2980_),
    .Y(_3008_)
);

OAI21X1 _13041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2946_),
    .B(_2944_),
    .C(_3008_),
    .Y(_3009_)
);

OR2X2 _13042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3009_),
    .B(_2987_),
    .Y(_3010_)
);

AOI21X1 _13043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2987_),
    .B(_3009_),
    .C(_2702_),
    .Y(_3011_)
);

NAND2X1 _13044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf1 ),
    .B(_2727_),
    .Y(_3012_)
);

NAND2X1 _13045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495__bF$buf6),
    .B(_2767_),
    .Y(_3013_)
);

AOI21X1 _13046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3012_),
    .B(_3013_),
    .C(_2497__bF$buf3),
    .Y(_3014_)
);

INVX2 _13047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2659_),
    .Y(_3015_)
);

MUX2X1 _13048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2773_),
    .B(_2753_),
    .S(\datapath.alu.b_2_bF$buf0 ),
    .Y(_3016_)
);

OAI21X1 _13049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3016_),
    .B(\datapath.alu.b_3_bF$buf1 ),
    .C(_3015_),
    .Y(_3017_)
);

MUX2X1 _13050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [4]),
    .B(\datapath.alu.a [5]),
    .S(\datapath.alu.b_0_bF$buf1 ),
    .Y(_3018_)
);

NAND2X1 _13051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf1),
    .B(_3018_),
    .Y(_3019_)
);

OAI21X1 _13052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf0),
    .B(_2885_),
    .C(_3019_),
    .Y(_3020_)
);

MUX2X1 _13053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3020_),
    .B(_2792_),
    .S(_2495__bF$buf5),
    .Y(_3021_)
);

NAND2X1 _13054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf2),
    .B(_3021_),
    .Y(_3022_)
);

OAI22X1 _13055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3014_),
    .B(_3017_),
    .C(_3022_),
    .D(_2884_),
    .Y(_3023_)
);

AOI21X1 _13056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3011_),
    .B(_3010_),
    .C(_3023_),
    .Y(_3024_)
);

NAND3X1 _13057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3007_),
    .B(_2990_),
    .C(_3024_),
    .Y(\datapath.alu.c [5])
);

XOR2X1 _13058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [6]),
    .B(\datapath.alu.b [6]),
    .Y(_3025_)
);

AOI21X1 _13059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2980_),
    .B(_2987_),
    .C(_2998_),
    .Y(_3026_)
);

OAI21X1 _13060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2935_),
    .B(_2936_),
    .C(_2987_),
    .Y(_3027_)
);

OAI21X1 _13061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2946_),
    .B(_3027_),
    .C(_3026_),
    .Y(_3028_)
);

OAI21X1 _13062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3028_),
    .B(_3025_),
    .C(_2703__bF$buf0),
    .Y(_3029_)
);

AOI21X1 _13063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3025_),
    .B(_3028_),
    .C(_3029_),
    .Y(_3030_)
);

OAI21X1 _13064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2508_),
    .B(_2936_),
    .C(_3001_),
    .Y(_3031_)
);

OAI21X1 _13065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2978_),
    .B(_2482_),
    .C(_3031_),
    .Y(_3032_)
);

OAI21X1 _13066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3032_),
    .B(_2473_),
    .C(_2799__bF$buf1),
    .Y(_3033_)
);

AOI21X1 _13067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2473_),
    .B(_3032_),
    .C(_3033_),
    .Y(_3034_)
);

NAND2X1 _13068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf7 ),
    .B(_2826_),
    .Y(_3035_)
);

NAND2X1 _13069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495__bF$buf4),
    .B(_2815_),
    .Y(_3036_)
);

NAND3X1 _13070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf1),
    .B(_3035_),
    .C(_3036_),
    .Y(_3037_)
);

INVX1 _13071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2992_),
    .Y(_3038_)
);

NOR2X1 _13072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf6 ),
    .B(_2832_),
    .Y(_3039_)
);

OAI21X1 _13073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3039_),
    .B(_3038_),
    .C(\datapath.alu.b_3_bF$buf0 ),
    .Y(_3040_)
);

AOI21X1 _13074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3040_),
    .B(_3037_),
    .C(_2809_),
    .Y(_3041_)
);

NAND2X1 _13075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf6 ),
    .B(_3039_),
    .Y(_3042_)
);

AOI21X1 _13076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3042_),
    .B(_3037_),
    .C(_2808_),
    .Y(_3043_)
);

OAI21X1 _13077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3041_),
    .B(_3043_),
    .C(\datapath.alu.b_4_bF$buf4 ),
    .Y(_3044_)
);

NAND2X1 _13078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495__bF$buf3),
    .B(_2846_),
    .Y(_3045_)
);

OAI21X1 _13079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2841_),
    .B(_2842_),
    .C(\datapath.alu.b_2_bF$buf5 ),
    .Y(_3046_)
);

NAND2X1 _13080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3045_),
    .B(_3046_),
    .Y(_3047_)
);

NOR2X1 _13081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf5 ),
    .B(_3047_),
    .Y(_3048_)
);

NAND2X1 _13082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf4 ),
    .B(_2820_),
    .Y(_3049_)
);

OAI21X1 _13083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2838_),
    .B(_2839_),
    .C(_2495__bF$buf2),
    .Y(_3050_)
);

NAND2X1 _13084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3049_),
    .B(_3050_),
    .Y(_3051_)
);

NOR2X1 _13085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf0),
    .B(_3051_),
    .Y(_3052_)
);

OAI21X1 _13086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3052_),
    .B(_3048_),
    .C(_3015_),
    .Y(_3053_)
);

NAND2X1 _13087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf3 ),
    .B(_2852_),
    .Y(_3054_)
);

OAI21X1 _13088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2504_),
    .B(\datapath.alu.b_0_bF$buf0 ),
    .C(_2638_),
    .Y(_3055_)
);

NAND2X1 _13089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf7),
    .B(_3055_),
    .Y(_3056_)
);

OAI21X1 _13090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2475_),
    .B(\datapath.alu.b_0_bF$buf10 ),
    .C(_2627_),
    .Y(_3057_)
);

NAND2X1 _13091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf4 ),
    .B(_3057_),
    .Y(_3058_)
);

NAND3X1 _13092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495__bF$buf1),
    .B(_3056_),
    .C(_3058_),
    .Y(_3059_)
);

NAND3X1 _13093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf6),
    .B(_3059_),
    .C(_3054_),
    .Y(_3060_)
);

NOR2X1 _13094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884_),
    .B(_3060_),
    .Y(_3061_)
);

INVX2 _13095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [6]),
    .Y(_3062_)
);

OAI22X1 _13096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2504_),
    .B(_2694_),
    .C(_2708__bF$buf0),
    .D(_3062_),
    .Y(_3063_)
);

NOR2X1 _13097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2504_),
    .B(_3062_),
    .Y(_3064_)
);

INVX1 _13098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3064_),
    .Y(_3065_)
);

OAI22X1 _13099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2692_),
    .B(_3065_),
    .C(_2707_),
    .D(_2505_),
    .Y(_3066_)
);

NOR2X1 _13100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3063_),
    .B(_3066_),
    .Y(_3067_)
);

OAI21X1 _13101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2688__bF$buf1),
    .B(_3064_),
    .C(_2680__bF$buf1),
    .Y(_3068_)
);

OAI21X1 _13102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [6]),
    .B(\datapath.alu.b [6]),
    .C(_3068_),
    .Y(_3069_)
);

NAND2X1 _13103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3069_),
    .B(_3067_),
    .Y(_3070_)
);

NOR2X1 _13104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3070_),
    .B(_3061_),
    .Y(_3071_)
);

NAND3X1 _13105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3053_),
    .B(_3071_),
    .C(_3044_),
    .Y(_3072_)
);

NOR3X1 _13106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3030_),
    .B(_3034_),
    .C(_3072_),
    .Y(_3073_)
);

INVX2 _13107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3073_),
    .Y(\datapath.alu.c [6])
);

XOR2X1 _13108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [7]),
    .B(\datapath.alu.b [7]),
    .Y(_3074_)
);

INVX1 _13109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3026_),
    .Y(_3075_)
);

INVX1 _13110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3027_),
    .Y(_3076_)
);

AOI21X1 _13111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3076_),
    .B(_2942_),
    .C(_3075_),
    .Y(_3077_)
);

OAI21X1 _13112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3077_),
    .B(_2473_),
    .C(_3065_),
    .Y(_3078_)
);

OAI21X1 _13113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3078_),
    .B(_3074_),
    .C(_2703__bF$buf3),
    .Y(_3079_)
);

AOI21X1 _13114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3074_),
    .B(_3078_),
    .C(_3079_),
    .Y(_3080_)
);

NOR2X1 _13115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [6]),
    .B(_2504_),
    .Y(_3081_)
);

AOI21X1 _13116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2505_),
    .B(_3032_),
    .C(_3081_),
    .Y(_3082_)
);

AND2X2 _13117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3082_),
    .B(_3074_),
    .Y(_3083_)
);

OAI21X1 _13118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3082_),
    .B(_3074_),
    .C(_2799__bF$buf0),
    .Y(_3084_)
);

MUX2X1 _13119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2910_),
    .B(_2905_),
    .S(\datapath.alu.b_2_bF$buf2 ),
    .Y(_3085_)
);

NOR2X1 _13120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf5),
    .B(_1641_),
    .Y(_3086_)
);

AOI21X1 _13121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf4),
    .B(_3085_),
    .C(_3086_),
    .Y(_3087_)
);

AND2X2 _13122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2916_),
    .B(_2495__bF$buf0),
    .Y(_3088_)
);

MUX2X1 _13123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3085_),
    .B(_3088_),
    .S(_2497__bF$buf3),
    .Y(_3089_)
);

OAI22X1 _13124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3087_),
    .B(_2809_),
    .C(_2808_),
    .D(_3089_),
    .Y(_3090_)
);

MUX2X1 _13125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [18]),
    .B(\datapath.alu.a [17]),
    .S(\datapath.alu.b_0_bF$buf9 ),
    .Y(_3091_)
);

MUX2X1 _13126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2763_),
    .B(_3091_),
    .S(_2489__bF$buf6),
    .Y(_3092_)
);

MUX2X1 _13127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [22]),
    .B(\datapath.alu.a [21]),
    .S(\datapath.alu.b_0_bF$buf8 ),
    .Y(_3093_)
);

MUX2X1 _13128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2723_),
    .B(_3093_),
    .S(_2489__bF$buf5),
    .Y(_3094_)
);

MUX2X1 _13129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3094_),
    .B(_3092_),
    .S(\datapath.alu.b_2_bF$buf1 ),
    .Y(_3095_)
);

NAND2X1 _13130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf4 ),
    .B(_3095_),
    .Y(_3096_)
);

MUX2X1 _13131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [8]),
    .B(\datapath.alu.a [7]),
    .S(\datapath.alu.b_0_bF$buf7 ),
    .Y(_3097_)
);

MUX2X1 _13132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [10]),
    .B(\datapath.alu.a [9]),
    .S(\datapath.alu.b_0_bF$buf6 ),
    .Y(_3098_)
);

MUX2X1 _13133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3098_),
    .B(_3097_),
    .S(\datapath.alu.b_1_bF$buf3 ),
    .Y(_3099_)
);

MUX2X1 _13134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [14]),
    .B(\datapath.alu.a [13]),
    .S(\datapath.alu.b_0_bF$buf5 ),
    .Y(_3100_)
);

MUX2X1 _13135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [12]),
    .B(\datapath.alu.a [11]),
    .S(\datapath.alu.b_0_bF$buf4 ),
    .Y(_3101_)
);

MUX2X1 _13136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3101_),
    .B(_3100_),
    .S(_2489__bF$buf4),
    .Y(_3102_)
);

MUX2X1 _13137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3102_),
    .B(_3099_),
    .S(\datapath.alu.b_2_bF$buf0 ),
    .Y(_3103_)
);

NAND2X1 _13138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf2),
    .B(_3103_),
    .Y(_3104_)
);

NAND3X1 _13139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3015_),
    .B(_3096_),
    .C(_3104_),
    .Y(_3105_)
);

NAND2X1 _13140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf2 ),
    .B(_3018_),
    .Y(_3106_)
);

OAI21X1 _13141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2502_),
    .B(\datapath.alu.b_0_bF$buf3 ),
    .C(_2751_),
    .Y(_3107_)
);

OAI21X1 _13142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf1 ),
    .B(_3107_),
    .C(_3106_),
    .Y(_3108_)
);

MUX2X1 _13143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3108_),
    .B(_2886_),
    .S(_2495__bF$buf6),
    .Y(_3109_)
);

NAND3X1 _13144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf1),
    .B(_2701_),
    .C(_3109_),
    .Y(_3110_)
);

OAI21X1 _13145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2707_),
    .B(\datapath.alu.a [7]),
    .C(_2708__bF$buf3),
    .Y(_3111_)
);

NAND2X1 _13146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2502_),
    .B(_2503_),
    .Y(_3112_)
);

NOR2X1 _13147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2801_),
    .B(_2715_),
    .Y(_3113_)
);

INVX8 _13148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2688__bF$buf0),
    .Y(_3114_)
);

AOI22X1 _13149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3112_),
    .B(_3113_),
    .C(_3114_),
    .D(_3074_),
    .Y(_3115_)
);

AOI21X1 _13150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [7]),
    .B(_2865__bF$buf1),
    .C(_2869__bF$buf1),
    .Y(_3116_)
);

OAI21X1 _13151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3116_),
    .B(_2502_),
    .C(_3115_),
    .Y(_3117_)
);

AOI21X1 _13152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [7]),
    .B(_3111_),
    .C(_3117_),
    .Y(_3118_)
);

NAND3X1 _13153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3110_),
    .B(_3118_),
    .C(_3105_),
    .Y(_3119_)
);

AOI21X1 _13154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_4_bF$buf3 ),
    .B(_3090_),
    .C(_3119_),
    .Y(_3120_)
);

OAI21X1 _13155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3083_),
    .B(_3084_),
    .C(_3120_),
    .Y(_3121_)
);

NOR2X1 _13156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3080_),
    .B(_3121_),
    .Y(_3122_)
);

INVX2 _13157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3122_),
    .Y(\datapath.alu.c [7])
);

NAND2X1 _13158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3074_),
    .B(_3025_),
    .Y(_3123_)
);

NOR2X1 _13159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3123_),
    .B(_3027_),
    .Y(_3124_)
);

NOR2X1 _13160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2502_),
    .B(_2503_),
    .Y(_3125_)
);

AOI21X1 _13161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3112_),
    .B(_3064_),
    .C(_3125_),
    .Y(_3126_)
);

OAI21X1 _13162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3026_),
    .B(_3123_),
    .C(_3126_),
    .Y(_3127_)
);

AOI21X1 _13163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3124_),
    .B(_2942_),
    .C(_3127_),
    .Y(_3128_)
);

AOI21X1 _13164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2468_),
    .B(_3128_),
    .C(_2702_),
    .Y(_3129_)
);

OAI21X1 _13165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2468_),
    .B(_3128_),
    .C(_3129_),
    .Y(_3130_)
);

MUX2X1 _13166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2922_),
    .B(_2928_),
    .S(_2495__bF$buf5),
    .Y(_3131_)
);

AOI22X1 _13167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2717_),
    .B(_3086_),
    .C(_3131_),
    .D(_2497__bF$buf0),
    .Y(_3132_)
);

NOR3X1 _13168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf4),
    .B(_2676_),
    .C(_3132_),
    .Y(_3133_)
);

NOR2X1 _13169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2599_),
    .B(_2515_),
    .Y(_3134_)
);

AOI22X1 _13170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2516_),
    .B(_2706__bF$buf2),
    .C(_2865__bF$buf0),
    .D(_3134_),
    .Y(_3135_)
);

AOI22X1 _13171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [8]),
    .B(_2802_),
    .C(_2869__bF$buf0),
    .D(\datapath.alu.a [8]),
    .Y(_3136_)
);

NAND2X1 _13172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3135_),
    .B(_3136_),
    .Y(_3137_)
);

OAI21X1 _13173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2599_),
    .B(_2515_),
    .C(_3114_),
    .Y(_3138_)
);

AOI22X1 _13174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2599_),
    .B(_2515_),
    .C(_3138_),
    .D(_2680__bF$buf0),
    .Y(_3139_)
);

NOR3X1 _13175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3137_),
    .B(_3139_),
    .C(_3133_),
    .Y(_3140_)
);

OR2X2 _13176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2482_),
    .B(_2474_),
    .Y(_3141_)
);

NOR2X1 _13177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3074_),
    .B(_3025_),
    .Y(_3142_)
);

OAI21X1 _13178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2987_),
    .B(_2481_),
    .C(_2479_),
    .Y(_3143_)
);

NAND2X1 _13179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [6]),
    .B(_3062_),
    .Y(_3144_)
);

NOR2X1 _13180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [7]),
    .B(_2502_),
    .Y(_3145_)
);

INVX1 _13181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3145_),
    .Y(_3146_)
);

OAI21X1 _13182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3074_),
    .B(_3144_),
    .C(_3146_),
    .Y(_3147_)
);

AOI21X1 _13183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3142_),
    .B(_3143_),
    .C(_3147_),
    .Y(_3148_)
);

OAI21X1 _13184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3141_),
    .B(_2978_),
    .C(_3148_),
    .Y(_3149_)
);

NAND2X1 _13185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2468_),
    .B(_3149_),
    .Y(_3150_)
);

AOI21X1 _13186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3081_),
    .B(_2472_),
    .C(_3145_),
    .Y(_3151_)
);

OAI21X1 _13187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2474_),
    .B(_3031_),
    .C(_3151_),
    .Y(_3152_)
);

AOI21X1 _13188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2483_),
    .B(_2973_),
    .C(_3152_),
    .Y(_3153_)
);

AOI21X1 _13189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2602_),
    .B(_3153_),
    .C(_2798_),
    .Y(_3154_)
);

MUX2X1 _13190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3057_),
    .B(_2851_),
    .S(_2489__bF$buf3),
    .Y(_3155_)
);

OAI21X1 _13191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2599_),
    .B(\datapath.alu.b_0_bF$buf2 ),
    .C(_2636_),
    .Y(_3156_)
);

MUX2X1 _13192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3156_),
    .B(_3055_),
    .S(_2489__bF$buf2),
    .Y(_3157_)
);

MUX2X1 _13193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3157_),
    .B(_3155_),
    .S(_2495__bF$buf4),
    .Y(_3158_)
);

OAI21X1 _13194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2697_),
    .B(\datapath.alu.b_2_bF$buf7 ),
    .C(\datapath.alu.b_3_bF$buf3 ),
    .Y(_3159_)
);

OAI21X1 _13195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3158_),
    .B(\datapath.alu.b_3_bF$buf2 ),
    .C(_3159_),
    .Y(_3160_)
);

MUX2X1 _13196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2837_),
    .B(_2819_),
    .S(_2489__bF$buf1),
    .Y(_3161_)
);

MUX2X1 _13197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3161_),
    .B(_2924_),
    .S(_2495__bF$buf3),
    .Y(_3162_)
);

MUX2X1 _13198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3162_),
    .B(_2654_),
    .S(\datapath.alu.b_3_bF$buf1 ),
    .Y(_3163_)
);

OAI22X1 _13199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3160_),
    .B(_2884_),
    .C(_3163_),
    .D(_2659_),
    .Y(_3164_)
);

AOI21X1 _13200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3150_),
    .B(_3154_),
    .C(_3164_),
    .Y(_3165_)
);

NAND3X1 _13201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3130_),
    .B(_3165_),
    .C(_3140_),
    .Y(\datapath.alu.c [8])
);

OR2X2 _13202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3027_),
    .B(_3123_),
    .Y(_3166_)
);

INVX1 _13203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3127_),
    .Y(_3167_)
);

OAI21X1 _13204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2946_),
    .B(_3166_),
    .C(_3167_),
    .Y(_3168_)
);

AOI21X1 _13205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2602_),
    .B(_3168_),
    .C(_3134_),
    .Y(_3169_)
);

AOI21X1 _13206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2467_),
    .B(_3169_),
    .C(_2702_),
    .Y(_3170_)
);

OAI21X1 _13207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2467_),
    .B(_3169_),
    .C(_3170_),
    .Y(_3171_)
);

INVX1 _13208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3086_),
    .Y(_3172_)
);

OAI21X1 _13209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2740_),
    .B(\datapath.alu.b_3_bF$buf0 ),
    .C(_3172_),
    .Y(_3173_)
);

NOR2X1 _13210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf6 ),
    .B(_2808_),
    .Y(_3174_)
);

INVX1 _13211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3174_),
    .Y(_3175_)
);

NOR2X1 _13212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3175_),
    .B(_2745_),
    .Y(_3176_)
);

AOI21X1 _13213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2717_),
    .B(_3173_),
    .C(_3176_),
    .Y(_3177_)
);

OAI21X1 _13214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2792_),
    .B(\datapath.alu.b_2_bF$buf6 ),
    .C(\datapath.alu.b_3_bF$buf5 ),
    .Y(_3178_)
);

MUX2X1 _13215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [8]),
    .B(\datapath.alu.a [9]),
    .S(\datapath.alu.b_0_bF$buf1 ),
    .Y(_3179_)
);

NAND2X1 _13216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf0),
    .B(_3179_),
    .Y(_3180_)
);

OAI21X1 _13217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf7),
    .B(_3107_),
    .C(_3180_),
    .Y(_3181_)
);

MUX2X1 _13218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3181_),
    .B(_3020_),
    .S(_2495__bF$buf2),
    .Y(_3182_)
);

OAI21X1 _13219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3182_),
    .B(\datapath.alu.b_3_bF$buf4 ),
    .C(_3178_),
    .Y(_3183_)
);

NOR2X1 _13220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884_),
    .B(_3183_),
    .Y(_3184_)
);

NOR2X1 _13221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2596_),
    .B(_2512_),
    .Y(_3185_)
);

OAI21X1 _13222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2688__bF$buf3),
    .B(_3185_),
    .C(_2680__bF$buf3),
    .Y(_3186_)
);

OAI21X1 _13223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [9]),
    .B(\datapath.alu.b [9]),
    .C(_3186_),
    .Y(_3187_)
);

AOI22X1 _13224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2513_),
    .B(_2706__bF$buf1),
    .C(_2865__bF$buf3),
    .D(_3185_),
    .Y(_3188_)
);

NAND2X1 _13225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [9]),
    .B(_2869__bF$buf3),
    .Y(_3189_)
);

NAND3X1 _13226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3188_),
    .B(_3189_),
    .C(_3187_),
    .Y(_3190_)
);

NOR2X1 _13227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3190_),
    .B(_3184_),
    .Y(_3191_)
);

OAI21X1 _13228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf3),
    .B(_3177_),
    .C(_3191_),
    .Y(_3192_)
);

OAI21X1 _13229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3153_),
    .B(_2516_),
    .C(_2601_),
    .Y(_3193_)
);

NOR2X1 _13230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2467_),
    .B(_3193_),
    .Y(_3194_)
);

INVX2 _13231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2601_),
    .Y(_3195_)
);

AOI21X1 _13232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2467_),
    .B(_3195_),
    .C(_2798_),
    .Y(_3196_)
);

OAI21X1 _13233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3153_),
    .B(_2469_),
    .C(_3196_),
    .Y(_3197_)
);

OAI21X1 _13234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2728_),
    .B(_2497__bF$buf6),
    .C(_3015_),
    .Y(_3198_)
);

AOI21X1 _13235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf5),
    .B(_2775_),
    .C(_3198_),
    .Y(_3199_)
);

AOI21X1 _13236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [9]),
    .B(_2802_),
    .C(_3199_),
    .Y(_3200_)
);

OAI21X1 _13237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3197_),
    .B(_3194_),
    .C(_3200_),
    .Y(_3201_)
);

NOR2X1 _13238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3192_),
    .B(_3201_),
    .Y(_3202_)
);

NAND2X1 _13239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3171_),
    .B(_3202_),
    .Y(\datapath.alu.c [9])
);

AOI21X1 _13240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3134_),
    .B(_2598_),
    .C(_3185_),
    .Y(_3203_)
);

NAND2X1 _13241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2945_),
    .B(_2862_),
    .Y(_3204_)
);

AOI21X1 _13242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2941_),
    .B(_3204_),
    .C(_3166_),
    .Y(_3205_)
);

NOR2X1 _13243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2467_),
    .B(_2468_),
    .Y(_3206_)
);

OAI21X1 _13244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3205_),
    .B(_3127_),
    .C(_3206_),
    .Y(_3207_)
);

NAND3X1 _13245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2594_),
    .B(_3203_),
    .C(_3207_),
    .Y(_3208_)
);

OAI21X1 _13246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3195_),
    .B(_2516_),
    .C(_2598_),
    .Y(_3209_)
);

OAI21X1 _13247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3128_),
    .B(_3209_),
    .C(_3203_),
    .Y(_3210_)
);

NAND2X1 _13248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465_),
    .B(_3210_),
    .Y(_3211_)
);

AOI21X1 _13249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3208_),
    .B(_3211_),
    .C(_2702_),
    .Y(_3212_)
);

NAND2X1 _13250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2603_),
    .B(_3149_),
    .Y(_3213_)
);

INVX1 _13251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2514_),
    .Y(_3214_)
);

AOI21X1 _13252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2597_),
    .B(_3195_),
    .C(_3214_),
    .Y(_3215_)
);

AOI21X1 _13253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3215_),
    .B(_3213_),
    .C(_2594_),
    .Y(_3216_)
);

OAI21X1 _13254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3153_),
    .B(_2469_),
    .C(_3215_),
    .Y(_3217_)
);

OAI21X1 _13255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3217_),
    .B(_2465_),
    .C(_2799__bF$buf3),
    .Y(_3218_)
);

NOR2X1 _13256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3216_),
    .B(_3218_),
    .Y(_3219_)
);

AOI21X1 _13257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf4),
    .B(_2830_),
    .C(_3086_),
    .Y(_3220_)
);

NAND2X1 _13258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2833_),
    .B(_3174_),
    .Y(_3221_)
);

OAI21X1 _13259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3220_),
    .B(_2809_),
    .C(_3221_),
    .Y(_3222_)
);

NAND2X1 _13260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_4_bF$buf2 ),
    .B(_3222_),
    .Y(_3223_)
);

NAND3X1 _13261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf3),
    .B(_2843_),
    .C(_2840_),
    .Y(_3224_)
);

NAND2X1 _13262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf3 ),
    .B(_2821_),
    .Y(_3225_)
);

AOI21X1 _13263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3225_),
    .B(_3224_),
    .C(_2659_),
    .Y(_3226_)
);

INVX1 _13264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3226_),
    .Y(_3227_)
);

NOR2X1 _13265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648_),
    .B(_2518_),
    .Y(_3228_)
);

OAI21X1 _13266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2688__bF$buf2),
    .B(_3228_),
    .C(_2680__bF$buf2),
    .Y(_3229_)
);

OAI21X1 _13267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [10]),
    .B(\datapath.alu.b [10]),
    .C(_3229_),
    .Y(_3230_)
);

AOI22X1 _13268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2865__bF$buf2),
    .B(_3228_),
    .C(\datapath.alu.b [10]),
    .D(_2802_),
    .Y(_3231_)
);

AOI22X1 _13269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519_),
    .B(_2706__bF$buf0),
    .C(_2869__bF$buf2),
    .D(\datapath.alu.a [10]),
    .Y(_3232_)
);

NAND3X1 _13270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3231_),
    .B(_3232_),
    .C(_3230_),
    .Y(_3233_)
);

NAND2X1 _13271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf2 ),
    .B(_2853_),
    .Y(_3234_)
);

NAND3X1 _13272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf5 ),
    .B(_3056_),
    .C(_3058_),
    .Y(_3235_)
);

OAI21X1 _13273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648_),
    .B(\datapath.alu.b_0_bF$buf0 ),
    .C(_2651_),
    .Y(_3236_)
);

NAND2X1 _13274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf6),
    .B(_3236_),
    .Y(_3237_)
);

NAND2X1 _13275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf0 ),
    .B(_3156_),
    .Y(_3238_)
);

NAND3X1 _13276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495__bF$buf1),
    .B(_3237_),
    .C(_3238_),
    .Y(_3239_)
);

NAND3X1 _13277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf2),
    .B(_3235_),
    .C(_3239_),
    .Y(_3240_)
);

AOI21X1 _13278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3234_),
    .B(_3240_),
    .C(_2884_),
    .Y(_3241_)
);

NOR2X1 _13279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3233_),
    .B(_3241_),
    .Y(_1591_)
);

NAND3X1 _13280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3227_),
    .B(_1591_),
    .C(_3223_),
    .Y(_1592_)
);

NOR3X1 _13281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3219_),
    .B(_1592_),
    .C(_3212_),
    .Y(_1593_)
);

INVX2 _13282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1593_),
    .Y(\datapath.alu.c [10])
);

AND2X2 _13283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2463_),
    .B(_2460_),
    .Y(_1594_)
);

NAND2X1 _13284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [10]),
    .B(_2518_),
    .Y(_1595_)
);

INVX4 _13285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1595_),
    .Y(_1596_)
);

OAI21X1 _13286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519_),
    .B(_1596_),
    .C(_3210_),
    .Y(_1597_)
);

OAI21X1 _13287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648_),
    .B(_2518_),
    .C(_1597_),
    .Y(_1598_)
);

OAI21X1 _13288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1598_),
    .B(_1594_),
    .C(_2703__bF$buf2),
    .Y(_1599_)
);

AOI21X1 _13289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1594_),
    .B(_1598_),
    .C(_1599_),
    .Y(_1600_)
);

NOR3X1 _13290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2464_),
    .B(_1596_),
    .C(_3216_),
    .Y(_1601_)
);

OAI21X1 _13291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3216_),
    .B(_1596_),
    .C(_2464_),
    .Y(_1602_)
);

NAND2X1 _13292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2799__bF$buf2),
    .B(_1602_),
    .Y(_1603_)
);

NOR2X1 _13293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf1),
    .B(_2909_),
    .Y(_1604_)
);

NOR2X1 _13294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2659_),
    .B(_1604_),
    .Y(_1605_)
);

OAI21X1 _13295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf1 ),
    .B(_2903_),
    .C(_1605_),
    .Y(_1606_)
);

OAI21X1 _13296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462_),
    .B(_2708__bF$buf2),
    .C(_1606_),
    .Y(_1607_)
);

AOI21X1 _13297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf0),
    .B(_2912_),
    .C(_3086_),
    .Y(_1608_)
);

NAND2X1 _13298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3174_),
    .B(_2918_),
    .Y(_1609_)
);

OAI21X1 _13299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1608_),
    .B(_2809_),
    .C(_1609_),
    .Y(_1610_)
);

NAND2X1 _13300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_4_bF$buf1 ),
    .B(_1610_),
    .Y(_1611_)
);

NAND2X1 _13301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf4 ),
    .B(_3108_),
    .Y(_1612_)
);

OAI21X1 _13302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2461_),
    .B(\datapath.alu.b_0_bF$buf10 ),
    .C(_2771_),
    .Y(_1613_)
);

NAND2X1 _13303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf5),
    .B(_1613_),
    .Y(_1614_)
);

OAI21X1 _13304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf4),
    .B(_3179_),
    .C(_1614_),
    .Y(_1615_)
);

OAI21X1 _13305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf3 ),
    .B(_1615_),
    .C(_1612_),
    .Y(_1616_)
);

NAND3X1 _13306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf0 ),
    .B(_2495__bF$buf0),
    .C(_2887_),
    .Y(_1617_)
);

OAI21X1 _13307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1616_),
    .B(\datapath.alu.b_3_bF$buf6 ),
    .C(_1617_),
    .Y(_1618_)
);

NAND2X1 _13308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2701_),
    .B(_1618_),
    .Y(_1619_)
);

INVX2 _13309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2460_),
    .Y(_1621_)
);

OAI21X1 _13310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1621_),
    .B(_2688__bF$buf1),
    .C(_2680__bF$buf1),
    .Y(_1622_)
);

AOI22X1 _13311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2520_),
    .B(_2706__bF$buf3),
    .C(_2865__bF$buf1),
    .D(_1621_),
    .Y(_1623_)
);

OAI21X1 _13312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2461_),
    .B(_2694_),
    .C(_1623_),
    .Y(_1624_)
);

AOI21X1 _13313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2463_),
    .B(_1622_),
    .C(_1624_),
    .Y(_1625_)
);

NAND3X1 _13314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1625_),
    .B(_1619_),
    .C(_1611_),
    .Y(_1626_)
);

NOR2X1 _13315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1607_),
    .B(_1626_),
    .Y(_1627_)
);

OAI21X1 _13316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1603_),
    .B(_1601_),
    .C(_1627_),
    .Y(_1628_)
);

NOR2X1 _13317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1628_),
    .B(_1600_),
    .Y(_1629_)
);

INVX2 _13318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1629_),
    .Y(\datapath.alu.c [11])
);

OAI21X1 _13319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [9]),
    .B(\datapath.alu.b [9]),
    .C(_3134_),
    .Y(_1631_)
);

OAI21X1 _13320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2596_),
    .B(_2512_),
    .C(_1631_),
    .Y(_1632_)
);

NOR2X1 _13321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465_),
    .B(_2464_),
    .Y(_1633_)
);

AOI21X1 _13322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2463_),
    .B(_3228_),
    .C(_1621_),
    .Y(_1634_)
);

INVX1 _13323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1634_),
    .Y(_1635_)
);

AOI21X1 _13324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1633_),
    .B(_1632_),
    .C(_1635_),
    .Y(_1636_)
);

OAI21X1 _13325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519_),
    .B(_1596_),
    .C(_1594_),
    .Y(_1637_)
);

NOR2X1 _13326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3209_),
    .B(_1637_),
    .Y(_1638_)
);

OAI21X1 _13327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3205_),
    .B(_3127_),
    .C(_1638_),
    .Y(_1639_)
);

NAND3X1 _13328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2591_),
    .B(_1636_),
    .C(_1639_),
    .Y(_1640_)
);

INVX2 _13329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2591_),
    .Y(_1642_)
);

NAND2X1 _13330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3206_),
    .B(_1633_),
    .Y(_1643_)
);

OAI21X1 _13331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3128_),
    .B(_1643_),
    .C(_1636_),
    .Y(_1644_)
);

NAND2X1 _13332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1642_),
    .B(_1644_),
    .Y(_1645_)
);

AOI21X1 _13333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1640_),
    .B(_1645_),
    .C(_2702_),
    .Y(_1646_)
);

OAI21X1 _13334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2513_),
    .B(_2601_),
    .C(_2514_),
    .Y(_1647_)
);

OAI21X1 _13335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2520_),
    .B(_1595_),
    .C(_2522_),
    .Y(_1648_)
);

AOI21X1 _13336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1647_),
    .B(_2595_),
    .C(_1648_),
    .Y(_1649_)
);

OAI21X1 _13337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3153_),
    .B(_2604_),
    .C(_1649_),
    .Y(_1650_)
);

OAI21X1 _13338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1650_),
    .B(_1642_),
    .C(_2799__bF$buf1),
    .Y(_1651_)
);

AOI21X1 _13339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1642_),
    .B(_1650_),
    .C(_1651_),
    .Y(_1653_)
);

OAI21X1 _13340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2929_),
    .B(_2927_),
    .C(_2497__bF$buf6),
    .Y(_1654_)
);

AOI21X1 _13341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3172_),
    .B(_1654_),
    .C(_2809_),
    .Y(_1655_)
);

AND2X2 _13342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3174_),
    .B(_2929_),
    .Y(_1656_)
);

OAI21X1 _13343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1655_),
    .B(_1656_),
    .C(\datapath.alu.b_4_bF$buf0 ),
    .Y(_1657_)
);

MUX2X1 _13344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3161_),
    .B(_2647_),
    .S(\datapath.alu.b_2_bF$buf2 ),
    .Y(_1658_)
);

NAND2X1 _13345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf5),
    .B(_1658_),
    .Y(_1659_)
);

NAND3X1 _13346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf5 ),
    .B(_2923_),
    .C(_2925_),
    .Y(_1660_)
);

AOI21X1 _13347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1660_),
    .B(_1659_),
    .C(_2676_),
    .Y(_1661_)
);

NAND2X1 _13348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495__bF$buf6),
    .B(_3155_),
    .Y(_1662_)
);

NAND3X1 _13349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf4 ),
    .B(_2966_),
    .C(_1662_),
    .Y(_1664_)
);

NAND2X1 _13350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf1 ),
    .B(_3157_),
    .Y(_1665_)
);

OAI21X1 _13351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2451_),
    .B(\datapath.alu.b_0_bF$buf9 ),
    .C(_2649_),
    .Y(_1666_)
);

NAND2X1 _13352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf3),
    .B(_1666_),
    .Y(_1667_)
);

NAND2X1 _13353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf6 ),
    .B(_3236_),
    .Y(_1668_)
);

NAND3X1 _13354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495__bF$buf5),
    .B(_1667_),
    .C(_1668_),
    .Y(_1669_)
);

NAND3X1 _13355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf4),
    .B(_1669_),
    .C(_1665_),
    .Y(_1670_)
);

AOI21X1 _13356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1664_),
    .B(_1670_),
    .C(_2700_),
    .Y(_1671_)
);

OAI21X1 _13357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1661_),
    .B(_1671_),
    .C(_2480__bF$buf2),
    .Y(_1672_)
);

NOR2X1 _13358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2451_),
    .B(_2456_),
    .Y(_1673_)
);

AOI22X1 _13359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2528_),
    .B(_2706__bF$buf2),
    .C(_2865__bF$buf0),
    .D(_1673_),
    .Y(_1675_)
);

AOI22X1 _13360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [12]),
    .B(_2802_),
    .C(_2869__bF$buf1),
    .D(\datapath.alu.a [12]),
    .Y(_1676_)
);

NAND2X1 _13361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1675_),
    .B(_1676_),
    .Y(_1677_)
);

NAND2X1 _13362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2451_),
    .B(_2456_),
    .Y(_1678_)
);

OAI21X1 _13363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2688__bF$buf0),
    .B(_1673_),
    .C(_2680__bF$buf0),
    .Y(_1679_)
);

AOI21X1 _13364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1678_),
    .B(_1679_),
    .C(_1677_),
    .Y(_1680_)
);

NAND3X1 _13365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1672_),
    .B(_1680_),
    .C(_1657_),
    .Y(_1681_)
);

NOR3X1 _13366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1653_),
    .B(_1681_),
    .C(_1646_),
    .Y(_1682_)
);

INVX2 _13367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1682_),
    .Y(\datapath.alu.c [12])
);

OAI21X1 _13368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1637_),
    .B(_3203_),
    .C(_1634_),
    .Y(_1683_)
);

AOI21X1 _13369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1638_),
    .B(_3168_),
    .C(_1683_),
    .Y(_1685_)
);

INVX1 _13370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1673_),
    .Y(_1686_)
);

OAI21X1 _13371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_),
    .B(_1642_),
    .C(_1686_),
    .Y(_1687_)
);

OAI21X1 _13372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1687_),
    .B(_2590_),
    .C(_2703__bF$buf1),
    .Y(_1688_)
);

AOI21X1 _13373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2590_),
    .B(_1687_),
    .C(_1688_),
    .Y(_1689_)
);

NAND2X1 _13374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1642_),
    .B(_1650_),
    .Y(_1690_)
);

AOI21X1 _13375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2457_),
    .B(_1690_),
    .C(_2590_),
    .Y(_1691_)
);

INVX1 _13376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2590_),
    .Y(_1692_)
);

OAI21X1 _13377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2451_),
    .B(\datapath.alu.b [12]),
    .C(_1690_),
    .Y(_1693_)
);

OAI21X1 _13378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1693_),
    .B(_1692_),
    .C(_2799__bF$buf0),
    .Y(_1694_)
);

AOI21X1 _13379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf3),
    .B(_2993_),
    .C(_3086_),
    .Y(_1696_)
);

NAND2X1 _13380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2995_),
    .B(_3174_),
    .Y(_1697_)
);

OAI21X1 _13381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1696_),
    .B(_2809_),
    .C(_1697_),
    .Y(_1698_)
);

OR2X2 _13382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2991_),
    .B(_2497__bF$buf2),
    .Y(_1699_)
);

OAI21X1 _13383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2768_),
    .B(\datapath.alu.b_2_bF$buf0 ),
    .C(_3012_),
    .Y(_1700_)
);

AOI21X1 _13384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf1),
    .B(_1700_),
    .C(_2659_),
    .Y(_1701_)
);

OAI21X1 _13385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2707_),
    .B(\datapath.alu.a [13]),
    .C(_2708__bF$buf1),
    .Y(_1702_)
);

NAND2X1 _13386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2452_),
    .B(_2454_),
    .Y(_1703_)
);

NOR2X1 _13387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2452_),
    .B(_2454_),
    .Y(_1704_)
);

OAI21X1 _13388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2688__bF$buf3),
    .B(_1704_),
    .C(_2680__bF$buf3),
    .Y(_1705_)
);

AOI22X1 _13389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1703_),
    .B(_1705_),
    .C(_1702_),
    .D(\datapath.alu.b [13]),
    .Y(_1707_)
);

AOI21X1 _13390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [13]),
    .B(_2865__bF$buf3),
    .C(_2869__bF$buf0),
    .Y(_1708_)
);

OAI21X1 _13391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2452_),
    .B(_1708_),
    .C(_1707_),
    .Y(_1709_)
);

AOI21X1 _13392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1699_),
    .B(_1701_),
    .C(_1709_),
    .Y(_1710_)
);

NAND2X1 _13393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf8 ),
    .B(_2451_),
    .Y(_1711_)
);

OAI21X1 _13394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf7 ),
    .B(\datapath.alu.a [13]),
    .C(_1711_),
    .Y(_1712_)
);

NAND2X1 _13395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf5 ),
    .B(_1613_),
    .Y(_1713_)
);

OAI21X1 _13396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1712_),
    .B(\datapath.alu.b_1_bF$buf4 ),
    .C(_1713_),
    .Y(_1714_)
);

NAND2X1 _13397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495__bF$buf4),
    .B(_1714_),
    .Y(_1715_)
);

OAI21X1 _13398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495__bF$buf3),
    .B(_3181_),
    .C(_1715_),
    .Y(_1716_)
);

MUX2X1 _13399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1716_),
    .B(_3021_),
    .S(_2497__bF$buf0),
    .Y(_1718_)
);

OAI21X1 _13400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884_),
    .B(_1718_),
    .C(_1710_),
    .Y(_1719_)
);

AOI21X1 _13401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_4_bF$buf4 ),
    .B(_1698_),
    .C(_1719_),
    .Y(_1720_)
);

OAI21X1 _13402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1694_),
    .B(_1691_),
    .C(_1720_),
    .Y(_1721_)
);

NOR2X1 _13403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1689_),
    .B(_1721_),
    .Y(_1722_)
);

INVX2 _13404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1722_),
    .Y(\datapath.alu.c [13])
);

INVX2 _13405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2587_),
    .Y(_1723_)
);

NAND2X1 _13406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2590_),
    .B(_2591_),
    .Y(_1724_)
);

AOI21X1 _13407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1703_),
    .B(_1673_),
    .C(_1704_),
    .Y(_1725_)
);

OAI21X1 _13408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_),
    .B(_1724_),
    .C(_1725_),
    .Y(_1726_)
);

OAI21X1 _13409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2532_),
    .B(_1723_),
    .C(_1726_),
    .Y(_1728_)
);

INVX1 _13410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1726_),
    .Y(_1729_)
);

AOI21X1 _13411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2449_),
    .B(_1729_),
    .C(_2702_),
    .Y(_1730_)
);

AOI21X1 _13412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2455_),
    .B(_2457_),
    .C(_2526_),
    .Y(_1731_)
);

AOI21X1 _13413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2592_),
    .B(_1650_),
    .C(_1731_),
    .Y(_1732_)
);

AND2X2 _13414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1732_),
    .B(_2588_),
    .Y(_1733_)
);

OAI21X1 _13415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1732_),
    .B(_2588_),
    .C(_2799__bF$buf3),
    .Y(_1734_)
);

INVX2 _13416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2700_),
    .Y(_1735_)
);

NAND3X1 _13417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf3 ),
    .B(_3059_),
    .C(_3054_),
    .Y(_1736_)
);

NAND3X1 _13418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf7 ),
    .B(_3237_),
    .C(_3238_),
    .Y(_1737_)
);

NAND2X1 _13419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf6 ),
    .B(_2452_),
    .Y(_1739_)
);

OAI21X1 _13420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf5 ),
    .B(\datapath.alu.a [14]),
    .C(_1739_),
    .Y(_1740_)
);

NAND2X1 _13421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf3 ),
    .B(_1666_),
    .Y(_1741_)
);

OAI21X1 _13422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1740_),
    .B(\datapath.alu.b_1_bF$buf2 ),
    .C(_1741_),
    .Y(_1742_)
);

OAI21X1 _13423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1742_),
    .B(\datapath.alu.b_2_bF$buf6 ),
    .C(_1737_),
    .Y(_1743_)
);

OAI21X1 _13424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1743_),
    .B(\datapath.alu.b_3_bF$buf2 ),
    .C(_1736_),
    .Y(_1744_)
);

NAND2X1 _13425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1735_),
    .B(_1744_),
    .Y(_1745_)
);

NOR2X1 _13426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf1 ),
    .B(_3051_),
    .Y(_1746_)
);

NAND2X1 _13427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3035_),
    .B(_3036_),
    .Y(_1747_)
);

NOR2X1 _13428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf6),
    .B(_1747_),
    .Y(_1748_)
);

OAI21X1 _13429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1746_),
    .B(_1748_),
    .C(_2658_),
    .Y(_1750_)
);

NAND2X1 _13430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1745_),
    .B(_1750_),
    .Y(_1751_)
);

OAI21X1 _13431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3039_),
    .B(_3038_),
    .C(_2497__bF$buf5),
    .Y(_1752_)
);

OAI21X1 _13432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf4),
    .B(_1641_),
    .C(_1752_),
    .Y(_1753_)
);

AOI22X1 _13433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3039_),
    .B(_3174_),
    .C(_1753_),
    .D(_2717_),
    .Y(_1754_)
);

NOR2X1 _13434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2530_),
    .B(_2586_),
    .Y(_1755_)
);

OAI21X1 _13435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2688__bF$buf2),
    .B(_1755_),
    .C(_2680__bF$buf2),
    .Y(_1756_)
);

OAI21X1 _13436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [14]),
    .B(\datapath.alu.b [14]),
    .C(_1756_),
    .Y(_1757_)
);

OAI21X1 _13437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586_),
    .B(_2708__bF$buf0),
    .C(_1757_),
    .Y(_1758_)
);

AOI22X1 _13438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2532_),
    .B(_2706__bF$buf1),
    .C(_2865__bF$buf2),
    .D(_1755_),
    .Y(_1759_)
);

OAI21X1 _13439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2530_),
    .B(_2694_),
    .C(_1759_),
    .Y(_1761_)
);

NOR2X1 _13440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1761_),
    .B(_1758_),
    .Y(_1762_)
);

OAI21X1 _13441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1754_),
    .B(_2480__bF$buf1),
    .C(_1762_),
    .Y(_1763_)
);

AOI21X1 _13442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf0),
    .B(_1751_),
    .C(_1763_),
    .Y(_1764_)
);

OAI21X1 _13443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1733_),
    .B(_1734_),
    .C(_1764_),
    .Y(_1765_)
);

AOI21X1 _13444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1728_),
    .B(_1730_),
    .C(_1765_),
    .Y(_1766_)
);

INVX2 _13445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1766_),
    .Y(\datapath.alu.c [14])
);

INVX1 _13446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1755_),
    .Y(_1767_)
);

AOI21X1 _13447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1767_),
    .B(_1728_),
    .C(_2448_),
    .Y(_1768_)
);

AND2X2 _13448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2447_),
    .B(_2444_),
    .Y(_1769_)
);

OAI21X1 _13449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2530_),
    .B(_2586_),
    .C(_1728_),
    .Y(_1771_)
);

OAI21X1 _13450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1771_),
    .B(_1769_),
    .C(_2703__bF$buf0),
    .Y(_1772_)
);

OAI21X1 _13451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1732_),
    .B(_2588_),
    .C(_2587_),
    .Y(_1773_)
);

XNOR2X1 _13452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1773_),
    .B(_1769_),
    .Y(_1774_)
);

NAND2X1 _13453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf0 ),
    .B(_3085_),
    .Y(_1775_)
);

OAI21X1 _13454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf6 ),
    .B(_3095_),
    .C(_1775_),
    .Y(_1776_)
);

OAI21X1 _13455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2445_),
    .B(\datapath.alu.b_0_bF$buf4 ),
    .C(_2765_),
    .Y(_1777_)
);

NAND2X1 _13456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf2),
    .B(_1777_),
    .Y(_1778_)
);

OAI21X1 _13457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1712_),
    .B(_2489__bF$buf1),
    .C(_1778_),
    .Y(_1779_)
);

MUX2X1 _13458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1779_),
    .B(_1615_),
    .S(_2495__bF$buf2),
    .Y(_1780_)
);

NAND2X1 _13459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf5 ),
    .B(_3109_),
    .Y(_1782_)
);

OAI21X1 _13460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf4 ),
    .B(_1780_),
    .C(_1782_),
    .Y(_1783_)
);

AOI22X1 _13461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2658_),
    .B(_1776_),
    .C(_1783_),
    .D(_1735_),
    .Y(_1784_)
);

NAND2X1 _13462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [31]),
    .B(_2717_),
    .Y(_1785_)
);

NAND2X1 _13463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf3),
    .B(_3088_),
    .Y(_1786_)
);

OAI21X1 _13464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1786_),
    .B(_2808_),
    .C(_1785_),
    .Y(_1787_)
);

OAI21X1 _13465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2707_),
    .B(\datapath.alu.a [15]),
    .C(_2708__bF$buf3),
    .Y(_1788_)
);

NAND2X1 _13466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [15]),
    .B(_1788_),
    .Y(_1789_)
);

AOI22X1 _13467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2447_),
    .B(_3113_),
    .C(_3114_),
    .D(_1769_),
    .Y(_1790_)
);

OAI21X1 _13468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2692_),
    .B(_2446_),
    .C(_2694_),
    .Y(_1791_)
);

NAND2X1 _13469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [15]),
    .B(_1791_),
    .Y(_1793_)
);

NAND3X1 _13470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1790_),
    .B(_1793_),
    .C(_1789_),
    .Y(_1794_)
);

AOI21X1 _13471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_4_bF$buf3 ),
    .B(_1787_),
    .C(_1794_),
    .Y(_1795_)
);

OAI21X1 _13472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1784_),
    .B(\datapath.alu.b_4_bF$buf2 ),
    .C(_1795_),
    .Y(_1796_)
);

AOI21X1 _13473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2799__bF$buf2),
    .B(_1774_),
    .C(_1796_),
    .Y(_1797_)
);

OAI21X1 _13474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1768_),
    .B(_1772_),
    .C(_1797_),
    .Y(\datapath.alu.c [15])
);

XNOR2X1 _13475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [16]),
    .B(\datapath.alu.b [16]),
    .Y(_1798_)
);

OAI21X1 _13476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2532_),
    .B(_1723_),
    .C(_1769_),
    .Y(_1799_)
);

NOR2X1 _13477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1724_),
    .B(_1799_),
    .Y(_1800_)
);

NAND2X1 _13478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1638_),
    .B(_1800_),
    .Y(_1801_)
);

INVX1 _13479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2444_),
    .Y(_1803_)
);

AOI21X1 _13480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2447_),
    .B(_1755_),
    .C(_1803_),
    .Y(_1804_)
);

OAI21X1 _13481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1799_),
    .B(_1725_),
    .C(_1804_),
    .Y(_1805_)
);

AOI21X1 _13482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1800_),
    .B(_1683_),
    .C(_1805_),
    .Y(_1806_)
);

OAI21X1 _13483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3128_),
    .B(_1801_),
    .C(_1806_),
    .Y(_1807_)
);

XNOR2X1 _13484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1807_),
    .B(_1798_),
    .Y(_1808_)
);

AOI21X1 _13485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1596_),
    .B(_2464_),
    .C(_2521_),
    .Y(_1809_)
);

OAI21X1 _13486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3215_),
    .B(_2466_),
    .C(_1809_),
    .Y(_1810_)
);

OAI21X1 _13487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2451_),
    .B(\datapath.alu.b [12]),
    .C(_2455_),
    .Y(_1811_)
);

OAI21X1 _13488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [13]),
    .B(_2454_),
    .C(_1811_),
    .Y(_1812_)
);

AOI21X1 _13489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1723_),
    .B(_2448_),
    .C(_2533_),
    .Y(_1814_)
);

OAI21X1 _13490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1812_),
    .B(_2450_),
    .C(_1814_),
    .Y(_1815_)
);

AOI21X1 _13491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2459_),
    .B(_1810_),
    .C(_1815_),
    .Y(_1816_)
);

OAI21X1 _13492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2471_),
    .B(_3153_),
    .C(_1816_),
    .Y(_1817_)
);

NOR2X1 _13493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1798_),
    .B(_1817_),
    .Y(_1818_)
);

INVX1 _13494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1798_),
    .Y(_1819_)
);

OAI21X1 _13495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2535_),
    .B(_2587_),
    .C(_2534_),
    .Y(_1820_)
);

AOI21X1 _13496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1731_),
    .B(_2589_),
    .C(_1820_),
    .Y(_1821_)
);

OAI21X1 _13497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2593_),
    .B(_1649_),
    .C(_1821_),
    .Y(_1822_)
);

AOI21X1 _13498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2605_),
    .B(_3149_),
    .C(_1822_),
    .Y(_1823_)
);

OAI21X1 _13499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1823_),
    .B(_1819_),
    .C(_2799__bF$buf1),
    .Y(_1825_)
);

OR2X2 _13500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1785_),
    .B(_2480__bF$buf5),
    .Y(_1826_)
);

OAI21X1 _13501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2692_),
    .B(_2071_),
    .C(_2708__bF$buf2),
    .Y(_1827_)
);

NAND2X1 _13502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [16]),
    .B(_1827_),
    .Y(_1828_)
);

NOR3X1 _13503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2801_),
    .B(_2060_),
    .C(_2715_),
    .Y(_1829_)
);

AND2X2 _13504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2706__bF$buf0),
    .B(_2541_),
    .Y(_1830_)
);

OAI22X1 _13505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2694_),
    .B(_2071_),
    .C(_2688__bF$buf1),
    .D(_1798_),
    .Y(_1831_)
);

NOR3X1 _13506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1829_),
    .B(_1830_),
    .C(_1831_),
    .Y(_1832_)
);

NAND3X1 _13507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1832_),
    .B(_1828_),
    .C(_1826_),
    .Y(_1833_)
);

AOI21X1 _13508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3015_),
    .B(_2675_),
    .C(_1833_),
    .Y(_1834_)
);

NAND2X1 _13509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1667_),
    .B(_1668_),
    .Y(_1836_)
);

NAND2X1 _13510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf5 ),
    .B(_1836_),
    .Y(_1837_)
);

MUX2X1 _13511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2445_),
    .B(_2071_),
    .S(\datapath.alu.b_0_bF$buf3 ),
    .Y(_1838_)
);

OR2X2 _13512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1838_),
    .B(\datapath.alu.b_1_bF$buf1 ),
    .Y(_1839_)
);

NAND2X1 _13513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf0 ),
    .B(_1740_),
    .Y(_1840_)
);

NAND3X1 _13514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495__bF$buf1),
    .B(_1839_),
    .C(_1840_),
    .Y(_1841_)
);

AOI21X1 _13515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1841_),
    .B(_1837_),
    .C(\datapath.alu.b_3_bF$buf3 ),
    .Y(_1842_)
);

MUX2X1 _13516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [5]),
    .B(\datapath.alu.a [6]),
    .S(\datapath.alu.b_0_bF$buf2 ),
    .Y(_1843_)
);

MUX2X1 _13517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [7]),
    .B(\datapath.alu.a [8]),
    .S(\datapath.alu.b_0_bF$buf1 ),
    .Y(_1844_)
);

MUX2X1 _13518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1844_),
    .B(_1843_),
    .S(_2489__bF$buf0),
    .Y(_1845_)
);

MUX2X1 _13519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1845_),
    .B(_2965_),
    .S(_2495__bF$buf0),
    .Y(_1847_)
);

OAI21X1 _13520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1847_),
    .B(_2497__bF$buf2),
    .C(_2480__bF$buf4),
    .Y(_1848_)
);

NOR2X1 _13521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf4 ),
    .B(_2697_),
    .Y(_1849_)
);

NAND2X1 _13522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf1),
    .B(_1849_),
    .Y(_1850_)
);

AOI21X1 _13523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_4_bF$buf1 ),
    .B(_1850_),
    .C(_2700_),
    .Y(_1851_)
);

OAI21X1 _13524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1842_),
    .B(_1848_),
    .C(_1851_),
    .Y(_1852_)
);

AND2X2 _13525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1834_),
    .B(_1852_),
    .Y(_1853_)
);

OAI21X1 _13526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1825_),
    .B(_1818_),
    .C(_1853_),
    .Y(_1854_)
);

AOI21X1 _13527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2703__bF$buf3),
    .B(_1808_),
    .C(_1854_),
    .Y(_1855_)
);

INVX2 _13528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1855_),
    .Y(\datapath.alu.c [16])
);

INVX1 _13529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2050_),
    .Y(_1857_)
);

INVX1 _13530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2092_),
    .Y(_1858_)
);

NOR2X1 _13531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2449_),
    .B(_2448_),
    .Y(_1859_)
);

NAND3X1 _13532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2590_),
    .B(_2591_),
    .C(_1859_),
    .Y(_1860_)
);

NOR2X1 _13533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1643_),
    .B(_1860_),
    .Y(_1861_)
);

INVX1 _13534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1725_),
    .Y(_1862_)
);

INVX1 _13535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1804_),
    .Y(_1863_)
);

AOI21X1 _13536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1859_),
    .B(_1862_),
    .C(_1863_),
    .Y(_1864_)
);

OAI21X1 _13537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1636_),
    .B(_1860_),
    .C(_1864_),
    .Y(_1865_)
);

AOI21X1 _13538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1861_),
    .B(_3168_),
    .C(_1865_),
    .Y(_1866_)
);

OAI21X1 _13539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1866_),
    .B(_2060_),
    .C(_1858_),
    .Y(_1868_)
);

OAI21X1 _13540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1868_),
    .B(_1857_),
    .C(_2703__bF$buf2),
    .Y(_1869_)
);

AOI21X1 _13541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1857_),
    .B(_1868_),
    .C(_1869_),
    .Y(_1870_)
);

NAND2X1 _13542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [16]),
    .B(_2082_),
    .Y(_1871_)
);

OAI21X1 _13543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1823_),
    .B(_1819_),
    .C(_1871_),
    .Y(_1872_)
);

AND2X2 _13544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1872_),
    .B(_2050_),
    .Y(_1873_)
);

OAI21X1 _13545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1872_),
    .B(_2050_),
    .C(_2799__bF$buf0),
    .Y(_1874_)
);

NAND2X1 _13546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf3 ),
    .B(_1714_),
    .Y(_1875_)
);

NAND2X1 _13547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf0 ),
    .B(_2071_),
    .Y(_1876_)
);

OAI21X1 _13548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf10 ),
    .B(\datapath.alu.a [17]),
    .C(_1876_),
    .Y(_1877_)
);

NAND2X1 _13549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf7),
    .B(_1877_),
    .Y(_1879_)
);

OAI21X1 _13550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf6),
    .B(_1777_),
    .C(_1879_),
    .Y(_1880_)
);

OAI21X1 _13551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1880_),
    .B(\datapath.alu.b_2_bF$buf2 ),
    .C(_1875_),
    .Y(_1881_)
);

MUX2X1 _13552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1881_),
    .B(_3182_),
    .S(_2497__bF$buf0),
    .Y(_1882_)
);

OAI21X1 _13553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2700_),
    .B(_1882_),
    .C(_2747_),
    .Y(_1883_)
);

INVX1 _13554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2794_),
    .Y(_1884_)
);

OAI21X1 _13555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2707_),
    .B(\datapath.alu.a [17]),
    .C(_2708__bF$buf1),
    .Y(_1885_)
);

OAI22X1 _13556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2017_),
    .B(_2694_),
    .C(_2692_),
    .D(_2007_),
    .Y(_1886_)
);

OAI21X1 _13557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [17]),
    .B(\datapath.alu.b [17]),
    .C(_3113_),
    .Y(_1887_)
);

OAI21X1 _13558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2050_),
    .B(_2688__bF$buf0),
    .C(_1887_),
    .Y(_1888_)
);

NOR2X1 _13559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1886_),
    .B(_1888_),
    .Y(_1890_)
);

OAI21X1 _13560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf3),
    .B(_1785_),
    .C(_1890_),
    .Y(_1891_)
);

AOI21X1 _13561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [17]),
    .B(_1885_),
    .C(_1891_),
    .Y(_1892_)
);

NOR2X1 _13562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf2),
    .B(_2700_),
    .Y(_1893_)
);

INVX4 _13563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1893_),
    .Y(_1894_)
);

OAI21X1 _13564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1884_),
    .B(_1894_),
    .C(_1892_),
    .Y(_1895_)
);

AOI21X1 _13565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf1),
    .B(_1883_),
    .C(_1895_),
    .Y(_1896_)
);

OAI21X1 _13566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1873_),
    .B(_1874_),
    .C(_1896_),
    .Y(_1897_)
);

NOR2X1 _13567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1870_),
    .B(_1897_),
    .Y(_1898_)
);

INVX2 _13568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1898_),
    .Y(\datapath.alu.c [17])
);

NOR2X1 _13569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1953_),
    .B(_1985_),
    .Y(_1900_)
);

INVX4 _13570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1900_),
    .Y(_1901_)
);

NOR2X1 _13571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1798_),
    .B(_2050_),
    .Y(_1902_)
);

OAI21X1 _13572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2050_),
    .B(_1858_),
    .C(_2007_),
    .Y(_1903_)
);

AOI21X1 _13573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1902_),
    .B(_1807_),
    .C(_1903_),
    .Y(_1904_)
);

OR2X2 _13574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1904_),
    .B(_1901_),
    .Y(_1905_)
);

AOI21X1 _13575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1901_),
    .B(_1904_),
    .C(_2702_),
    .Y(_1906_)
);

OAI21X1 _13576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2540_),
    .B(_1871_),
    .C(_2542_),
    .Y(_1907_)
);

INVX1 _13577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1907_),
    .Y(_1908_)
);

OAI21X1 _13578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1823_),
    .B(_2103_),
    .C(_1908_),
    .Y(_1909_)
);

NOR2X1 _13579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1901_),
    .B(_1909_),
    .Y(_1911_)
);

NAND2X1 _13580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1901_),
    .B(_1909_),
    .Y(_1912_)
);

NAND2X1 _13581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2799__bF$buf3),
    .B(_1912_),
    .Y(_1913_)
);

AOI22X1 _13582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2865__bF$buf1),
    .B(_1985_),
    .C(\datapath.alu.a [18]),
    .D(_2869__bF$buf3),
    .Y(_1914_)
);

AOI21X1 _13583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1964_),
    .B(_2706__bF$buf3),
    .C(_2802_),
    .Y(_1915_)
);

OAI21X1 _13584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1974_),
    .B(_1915_),
    .C(_1914_),
    .Y(_1916_)
);

OAI22X1 _13585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1953_),
    .B(_2680__bF$buf1),
    .C(_1901_),
    .D(_2688__bF$buf3),
    .Y(_1917_)
);

NOR2X1 _13586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1917_),
    .B(_1916_),
    .Y(_1918_)
);

AND2X2 _13587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1918_),
    .B(_1826_),
    .Y(_1919_)
);

AND2X2 _13588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3235_),
    .B(_3239_),
    .Y(_1920_)
);

NAND2X1 _13589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf6 ),
    .B(_1838_),
    .Y(_1922_)
);

MUX2X1 _13590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2017_),
    .B(_1964_),
    .S(\datapath.alu.b_0_bF$buf9 ),
    .Y(_1923_)
);

INVX1 _13591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1923_),
    .Y(_1924_)
);

OAI21X1 _13592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1924_),
    .B(\datapath.alu.b_1_bF$buf5 ),
    .C(_1922_),
    .Y(_1925_)
);

MUX2X1 _13593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1925_),
    .B(_1742_),
    .S(_2495__bF$buf6),
    .Y(_1926_)
);

NAND2X1 _13594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf6),
    .B(_1926_),
    .Y(_1927_)
);

OAI21X1 _13595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf5),
    .B(_1920_),
    .C(_1927_),
    .Y(_1928_)
);

AND2X2 _13596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1928_),
    .B(_2480__bF$buf0),
    .Y(_1929_)
);

AOI21X1 _13597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2853_),
    .B(_2854_),
    .C(_2701_),
    .Y(_1930_)
);

OAI21X1 _13598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1929_),
    .B(_1930_),
    .C(_1919_),
    .Y(_1931_)
);

AOI21X1 _13599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf5),
    .B(_2835_),
    .C(_1931_),
    .Y(_1933_)
);

OAI21X1 _13600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1911_),
    .B(_1913_),
    .C(_1933_),
    .Y(_1934_)
);

AOI21X1 _13601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1905_),
    .B(_1906_),
    .C(_1934_),
    .Y(_1935_)
);

INVX2 _13602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1935_),
    .Y(\datapath.alu.c [18])
);

NOR2X1 _13603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1942_),
    .B(_1932_),
    .Y(_1936_)
);

INVX2 _13604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1936_),
    .Y(_1937_)
);

INVX1 _13605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1985_),
    .Y(_1938_)
);

OAI21X1 _13606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1904_),
    .B(_1901_),
    .C(_1938_),
    .Y(_1939_)
);

AND2X2 _13607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1939_),
    .B(_1937_),
    .Y(_1940_)
);

NOR2X1 _13608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1937_),
    .B(_1939_),
    .Y(_1941_)
);

OAI21X1 _13609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1940_),
    .B(_1941_),
    .C(_2703__bF$buf1),
    .Y(_1943_)
);

NOR2X1 _13610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [18]),
    .B(_1964_),
    .Y(_1944_)
);

INVX1 _13611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1944_),
    .Y(_1945_)
);

NAND2X1 _13612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1945_),
    .B(_1912_),
    .Y(_1946_)
);

AOI21X1 _13613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1937_),
    .B(_1946_),
    .C(_2798_),
    .Y(_1947_)
);

OAI21X1 _13614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1937_),
    .B(_1946_),
    .C(_1947_),
    .Y(_1948_)
);

OAI22X1 _13615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2809_),
    .B(_2913_),
    .C(_2919_),
    .D(_2808_),
    .Y(_1949_)
);

OAI21X1 _13616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2707_),
    .B(\datapath.alu.a [19]),
    .C(_2708__bF$buf0),
    .Y(_1950_)
);

OAI21X1 _13617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [19]),
    .B(\datapath.alu.b [19]),
    .C(_3113_),
    .Y(_1951_)
);

AOI22X1 _13618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1932_),
    .B(_2865__bF$buf0),
    .C(_3114_),
    .D(_1936_),
    .Y(_1952_)
);

NAND3X1 _13619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1951_),
    .B(_1952_),
    .C(_1826_),
    .Y(_1954_)
);

AOI21X1 _13620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [19]),
    .B(_1950_),
    .C(_1954_),
    .Y(_1955_)
);

OAI21X1 _13621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1910_),
    .B(_2694_),
    .C(_1955_),
    .Y(_1956_)
);

AOI21X1 _13622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf4),
    .B(_1949_),
    .C(_1956_),
    .Y(_1957_)
);

NAND2X1 _13623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf8 ),
    .B(_1964_),
    .Y(_1958_)
);

OAI21X1 _13624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf7 ),
    .B(\datapath.alu.a [19]),
    .C(_1958_),
    .Y(_1959_)
);

MUX2X1 _13625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1959_),
    .B(_1877_),
    .S(_2489__bF$buf5),
    .Y(_1960_)
);

MUX2X1 _13626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1960_),
    .B(_1779_),
    .S(_2495__bF$buf5),
    .Y(_1961_)
);

NOR2X1 _13627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf2 ),
    .B(_1961_),
    .Y(_1962_)
);

OAI21X1 _13628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1616_),
    .B(_2497__bF$buf4),
    .C(_2480__bF$buf3),
    .Y(_1963_)
);

AOI21X1 _13629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_4_bF$buf0 ),
    .B(_2888_),
    .C(_2700_),
    .Y(_1965_)
);

OAI21X1 _13630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1963_),
    .B(_1962_),
    .C(_1965_),
    .Y(_1966_)
);

AND2X2 _13631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1957_),
    .B(_1966_),
    .Y(_1967_)
);

NAND3X1 _13632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1967_),
    .B(_1943_),
    .C(_1948_),
    .Y(\datapath.alu.c [19])
);

INVX2 _13633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1878_),
    .Y(_1968_)
);

INVX1 _13634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1903_),
    .Y(_1969_)
);

NAND2X1 _13635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1936_),
    .B(_1900_),
    .Y(_1970_)
);

AOI21X1 _13636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1985_),
    .B(_1936_),
    .C(_1932_),
    .Y(_1971_)
);

OAI21X1 _13637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1969_),
    .B(_1970_),
    .C(_1971_),
    .Y(_1972_)
);

OAI21X1 _13638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3205_),
    .B(_3127_),
    .C(_1861_),
    .Y(_1973_)
);

INVX1 _13639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1970_),
    .Y(_1975_)
);

NAND2X1 _13640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1902_),
    .B(_1975_),
    .Y(_1976_)
);

AOI21X1 _13641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1806_),
    .B(_1973_),
    .C(_1976_),
    .Y(_1977_)
);

OAI21X1 _13642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1977_),
    .B(_1972_),
    .C(_1968_),
    .Y(_1978_)
);

INVX1 _13643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1976_),
    .Y(_1979_)
);

AOI21X1 _13644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1979_),
    .B(_1807_),
    .C(_1972_),
    .Y(_1980_)
);

NAND2X1 _13645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1878_),
    .B(_1980_),
    .Y(_1981_)
);

NAND3X1 _13646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2703__bF$buf0),
    .B(_1978_),
    .C(_1981_),
    .Y(_1982_)
);

INVX1 _13647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2114_),
    .Y(_1983_)
);

NOR2X1 _13648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [19]),
    .B(_1910_),
    .Y(_1984_)
);

AOI21X1 _13649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2544_),
    .B(_1944_),
    .C(_1984_),
    .Y(_1986_)
);

OAI21X1 _13650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1908_),
    .B(_1996_),
    .C(_1986_),
    .Y(_1987_)
);

INVX1 _13651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1987_),
    .Y(_1988_)
);

OAI21X1 _13652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1823_),
    .B(_1983_),
    .C(_1988_),
    .Y(_1989_)
);

AOI21X1 _13653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1878_),
    .B(_1989_),
    .C(_2798_),
    .Y(_1990_)
);

OAI21X1 _13654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1878_),
    .B(_1989_),
    .C(_1990_),
    .Y(_1991_)
);

OAI21X1 _13655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2707_),
    .B(\datapath.alu.a [20]),
    .C(_2708__bF$buf3),
    .Y(_1992_)
);

INVX1 _13656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1867_),
    .Y(_1993_)
);

AOI22X1 _13657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1993_),
    .B(_2865__bF$buf3),
    .C(_1968_),
    .D(_3114_),
    .Y(_1994_)
);

AOI22X1 _13658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1856_),
    .B(_3113_),
    .C(_2869__bF$buf2),
    .D(\datapath.alu.a [20]),
    .Y(_1995_)
);

NAND2X1 _13659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1995_),
    .B(_1994_),
    .Y(_1997_)
);

AOI21X1 _13660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [20]),
    .B(_1992_),
    .C(_1997_),
    .Y(_1998_)
);

OAI21X1 _13661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2931_),
    .B(_2933_),
    .C(_2480__bF$buf2),
    .Y(_1999_)
);

NAND3X1 _13662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1826_),
    .B(_1998_),
    .C(_1999_),
    .Y(_2000_)
);

NAND2X1 _13663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf4 ),
    .B(_1923_),
    .Y(_2001_)
);

NAND2X1 _13664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf6 ),
    .B(_1910_),
    .Y(_2002_)
);

OAI21X1 _13665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf5 ),
    .B(\datapath.alu.a [20]),
    .C(_2002_),
    .Y(_2003_)
);

OAI21X1 _13666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2003_),
    .B(\datapath.alu.b_1_bF$buf3 ),
    .C(_2001_),
    .Y(_2004_)
);

OAI21X1 _13667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf2 ),
    .B(_1838_),
    .C(_1840_),
    .Y(_2005_)
);

NAND2X1 _13668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf1 ),
    .B(_2005_),
    .Y(_2006_)
);

OAI21X1 _13669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf0 ),
    .B(_2004_),
    .C(_2006_),
    .Y(_2008_)
);

AND2X2 _13670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1665_),
    .B(_1669_),
    .Y(_2009_)
);

AOI21X1 _13671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf1 ),
    .B(_2009_),
    .C(\datapath.alu.b_4_bF$buf4 ),
    .Y(_2010_)
);

OAI21X1 _13672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2008_),
    .B(\datapath.alu.b_3_bF$buf0 ),
    .C(_2010_),
    .Y(_2011_)
);

NOR2X1 _13673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf1),
    .B(_2968_),
    .Y(_2012_)
);

NOR2X1 _13674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2700_),
    .B(_2012_),
    .Y(_2013_)
);

AOI21X1 _13675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2011_),
    .B(_2013_),
    .C(_2000_),
    .Y(_2014_)
);

NAND3X1 _13676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1991_),
    .B(_2014_),
    .C(_1982_),
    .Y(\datapath.alu.c [20])
);

NOR2X1 _13677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1824_),
    .B(_1813_),
    .Y(_2015_)
);

INVX2 _13678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2015_),
    .Y(_2016_)
);

INVX1 _13679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1971_),
    .Y(_2018_)
);

AOI21X1 _13680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1975_),
    .B(_1903_),
    .C(_2018_),
    .Y(_2019_)
);

OAI21X1 _13681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1866_),
    .B(_1976_),
    .C(_2019_),
    .Y(_2020_)
);

AOI21X1 _13682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1968_),
    .B(_2020_),
    .C(_1993_),
    .Y(_2021_)
);

OR2X2 _13683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2021_),
    .B(_2016_),
    .Y(_2022_)
);

AOI21X1 _13684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2016_),
    .B(_2021_),
    .C(_2702_),
    .Y(_2023_)
);

OAI21X1 _13685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1835_),
    .B(\datapath.alu.b [20]),
    .C(_2015_),
    .Y(_2024_)
);

AOI21X1 _13686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1878_),
    .B(_1989_),
    .C(_2024_),
    .Y(_2025_)
);

AOI21X1 _13687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2114_),
    .B(_1817_),
    .C(_1987_),
    .Y(_2026_)
);

NOR2X1 _13688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [20]),
    .B(_1835_),
    .Y(_2027_)
);

AOI21X1 _13689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2027_),
    .B(_2016_),
    .C(_2798_),
    .Y(_2029_)
);

OAI21X1 _13690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2026_),
    .B(_1889_),
    .C(_2029_),
    .Y(_2030_)
);

NAND2X1 _13691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf4 ),
    .B(_1835_),
    .Y(_2031_)
);

OAI21X1 _13692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf3 ),
    .B(\datapath.alu.a [21]),
    .C(_2031_),
    .Y(_2032_)
);

NAND2X1 _13693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf4),
    .B(_2032_),
    .Y(_2033_)
);

NAND2X1 _13694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf1 ),
    .B(_1959_),
    .Y(_2034_)
);

NAND2X1 _13695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2033_),
    .B(_2034_),
    .Y(_2035_)
);

MUX2X1 _13696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1880_),
    .B(_2035_),
    .S(\datapath.alu.b_2_bF$buf7 ),
    .Y(_2036_)
);

MUX2X1 _13697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2036_),
    .B(_1716_),
    .S(_2497__bF$buf3),
    .Y(_2037_)
);

AND2X2 _13698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2037_),
    .B(_2480__bF$buf0),
    .Y(_2038_)
);

NAND2X1 _13699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_4_bF$buf3 ),
    .B(_3022_),
    .Y(_2040_)
);

NAND2X1 _13700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1735_),
    .B(_2040_),
    .Y(_2041_)
);

OAI21X1 _13701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2692_),
    .B(_2548_),
    .C(_2694_),
    .Y(_2042_)
);

OAI21X1 _13702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1813_),
    .B(_2688__bF$buf2),
    .C(_2680__bF$buf0),
    .Y(_2043_)
);

AOI21X1 _13703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [21]),
    .B(_2042_),
    .C(_2043_),
    .Y(_2044_)
);

INVX1 _13704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1826_),
    .Y(_2045_)
);

OAI21X1 _13705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2707_),
    .B(\datapath.alu.a [21]),
    .C(_2708__bF$buf2),
    .Y(_2046_)
);

AOI21X1 _13706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [21]),
    .B(_2046_),
    .C(_2045_),
    .Y(_2047_)
);

OAI21X1 _13707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1824_),
    .B(_2044_),
    .C(_2047_),
    .Y(_2048_)
);

INVX1 _13708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2048_),
    .Y(_2049_)
);

OAI21X1 _13709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2038_),
    .B(_2041_),
    .C(_2049_),
    .Y(_2051_)
);

AOI21X1 _13710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf5),
    .B(_2997_),
    .C(_2051_),
    .Y(_2052_)
);

OAI21X1 _13711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2030_),
    .B(_2025_),
    .C(_2052_),
    .Y(_2053_)
);

AOI21X1 _13712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2022_),
    .B(_2023_),
    .C(_2053_),
    .Y(_2054_)
);

INVX2 _13713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2054_),
    .Y(\datapath.alu.c [21])
);

AND2X2 _13714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1760_),
    .B(_1770_),
    .Y(_2055_)
);

NAND2X1 _13715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2015_),
    .B(_1968_),
    .Y(_2056_)
);

OAI21X1 _13716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1824_),
    .B(_1867_),
    .C(_1802_),
    .Y(_2057_)
);

INVX1 _13717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2057_),
    .Y(_2058_)
);

OAI21X1 _13718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1980_),
    .B(_2056_),
    .C(_2058_),
    .Y(_2059_)
);

NAND2X1 _13719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2055_),
    .B(_2059_),
    .Y(_2061_)
);

OR2X2 _13720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2059_),
    .B(_2055_),
    .Y(_2062_)
);

NAND3X1 _13721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2703__bF$buf3),
    .B(_2061_),
    .C(_2062_),
    .Y(_2063_)
);

AOI21X1 _13722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2027_),
    .B(_2016_),
    .C(_2552_),
    .Y(_2064_)
);

OAI21X1 _13723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2026_),
    .B(_1889_),
    .C(_2064_),
    .Y(_2065_)
);

NAND2X1 _13724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1781_),
    .B(_2065_),
    .Y(_2066_)
);

INVX1 _13725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1889_),
    .Y(_2067_)
);

INVX1 _13726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2064_),
    .Y(_2068_)
);

AOI21X1 _13727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2067_),
    .B(_1989_),
    .C(_2068_),
    .Y(_2069_)
);

AOI21X1 _13728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2055_),
    .B(_2069_),
    .C(_2798_),
    .Y(_2070_)
);

OR2X2 _13729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3041_),
    .B(_3043_),
    .Y(_2072_)
);

OAI21X1 _13730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2707_),
    .B(\datapath.alu.a [22]),
    .C(_2708__bF$buf1),
    .Y(_2073_)
);

OAI21X1 _13731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [22]),
    .B(\datapath.alu.b [22]),
    .C(_3113_),
    .Y(_2074_)
);

INVX1 _13732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1770_),
    .Y(_2075_)
);

AOI22X1 _13733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2075_),
    .B(_2865__bF$buf2),
    .C(_3114_),
    .D(_2055_),
    .Y(_2076_)
);

NAND3X1 _13734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2074_),
    .B(_2076_),
    .C(_1826_),
    .Y(_2077_)
);

AOI21X1 _13735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [22]),
    .B(_2073_),
    .C(_2077_),
    .Y(_2078_)
);

OAI21X1 _13736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1738_),
    .B(_2694_),
    .C(_2078_),
    .Y(_2079_)
);

AOI21X1 _13737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf4),
    .B(_2072_),
    .C(_2079_),
    .Y(_2080_)
);

MUX2X1 _13738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551_),
    .B(_1738_),
    .S(\datapath.alu.b_0_bF$buf2 ),
    .Y(_2081_)
);

NAND2X1 _13739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf3),
    .B(_2081_),
    .Y(_2083_)
);

OAI21X1 _13740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2003_),
    .B(_2489__bF$buf2),
    .C(_2083_),
    .Y(_2084_)
);

MUX2X1 _13741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2084_),
    .B(_1925_),
    .S(_2495__bF$buf4),
    .Y(_2085_)
);

NOR2X1 _13742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf6 ),
    .B(_2085_),
    .Y(_2086_)
);

OAI21X1 _13743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1743_),
    .B(_2497__bF$buf2),
    .C(_2480__bF$buf3),
    .Y(_2087_)
);

NAND2X1 _13744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_4_bF$buf2 ),
    .B(_3060_),
    .Y(_2088_)
);

OAI21X1 _13745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2086_),
    .B(_2087_),
    .C(_2088_),
    .Y(_2089_)
);

OAI21X1 _13746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2089_),
    .B(_2700_),
    .C(_2080_),
    .Y(_2090_)
);

AOI21X1 _13747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2066_),
    .B(_2070_),
    .C(_2090_),
    .Y(_2091_)
);

NAND2X1 _13748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2091_),
    .B(_2063_),
    .Y(\datapath.alu.c [22])
);

OAI21X1 _13749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1738_),
    .B(_1749_),
    .C(_2061_),
    .Y(_2093_)
);

XNOR2X1 _13750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2093_),
    .B(_1727_),
    .Y(_2094_)
);

AND2X2 _13751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1717_),
    .B(_1684_),
    .Y(_2095_)
);

NOR2X1 _13752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [22]),
    .B(_1738_),
    .Y(_2096_)
);

AOI21X1 _13753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1781_),
    .B(_2065_),
    .C(_2096_),
    .Y(_2097_)
);

AND2X2 _13754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2097_),
    .B(_2095_),
    .Y(_2098_)
);

OAI21X1 _13755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2097_),
    .B(_2095_),
    .C(_2799__bF$buf2),
    .Y(_2099_)
);

INVX1 _13756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3090_),
    .Y(_2100_)
);

NAND2X1 _13757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf6 ),
    .B(_1960_),
    .Y(_2101_)
);

MUX2X1 _13758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1738_),
    .B(_1695_),
    .S(\datapath.alu.b_0_bF$buf1 ),
    .Y(_2102_)
);

NAND2X1 _13759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf1),
    .B(_2102_),
    .Y(_2104_)
);

OAI21X1 _13760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2032_),
    .B(_2489__bF$buf0),
    .C(_2104_),
    .Y(_2105_)
);

NAND2X1 _13761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495__bF$buf3),
    .B(_2105_),
    .Y(_2106_)
);

NAND2X1 _13762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2101_),
    .B(_2106_),
    .Y(_2107_)
);

NAND2X1 _13763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf5 ),
    .B(_1780_),
    .Y(_2108_)
);

OAI21X1 _13764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2107_),
    .B(\datapath.alu.b_3_bF$buf4 ),
    .C(_2108_),
    .Y(_2109_)
);

OAI21X1 _13765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2700_),
    .B(_2109_),
    .C(_2100_),
    .Y(_2110_)
);

NAND2X1 _13766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf1),
    .B(_3109_),
    .Y(_2111_)
);

AOI21X1 _13767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1695_),
    .B(_2706__bF$buf2),
    .C(_2802_),
    .Y(_2112_)
);

OAI22X1 _13768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1727_),
    .B(_2688__bF$buf1),
    .C(_2692_),
    .D(_1684_),
    .Y(_2113_)
);

OAI21X1 _13769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [23]),
    .B(\datapath.alu.b [23]),
    .C(_3113_),
    .Y(_2115_)
);

OAI21X1 _13770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1785_),
    .B(_2480__bF$buf2),
    .C(_2115_),
    .Y(_2116_)
);

NOR2X1 _13771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2113_),
    .B(_2116_),
    .Y(_2117_)
);

OAI21X1 _13772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1706_),
    .B(_2112_),
    .C(_2117_),
    .Y(_2118_)
);

AOI21X1 _13773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [23]),
    .B(_2869__bF$buf1),
    .C(_2118_),
    .Y(_2119_)
);

OAI21X1 _13774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2111_),
    .B(_1894_),
    .C(_2119_),
    .Y(_2120_)
);

AOI21X1 _13775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf1),
    .B(_2110_),
    .C(_2120_),
    .Y(_2121_)
);

OAI21X1 _13776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2098_),
    .B(_2099_),
    .C(_2121_),
    .Y(_2122_)
);

AOI21X1 _13777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2703__bF$buf2),
    .B(_2094_),
    .C(_2122_),
    .Y(_2123_)
);

INVX2 _13778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2123_),
    .Y(\datapath.alu.c [23])
);

NOR2X1 _13779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_2439_),
    .Y(_2125_)
);

NAND2X1 _13780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2095_),
    .B(_2055_),
    .Y(_2126_)
);

NOR2X1 _13781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2126_),
    .B(_2056_),
    .Y(_2127_)
);

NAND2X1 _13782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2127_),
    .B(_1979_),
    .Y(_2128_)
);

OAI21X1 _13783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [23]),
    .B(\datapath.alu.b [23]),
    .C(_2075_),
    .Y(_2129_)
);

AND2X2 _13784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2129_),
    .B(_1684_),
    .Y(_2130_)
);

OAI21X1 _13785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2126_),
    .B(_2058_),
    .C(_2130_),
    .Y(_2131_)
);

AOI21X1 _13786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2127_),
    .B(_1972_),
    .C(_2131_),
    .Y(_2132_)
);

OAI21X1 _13787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1866_),
    .B(_2128_),
    .C(_2132_),
    .Y(_2133_)
);

NAND2X1 _13788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2125_),
    .B(_2133_),
    .Y(_2134_)
);

INVX2 _13789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2125_),
    .Y(_2136_)
);

INVX1 _13790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2127_),
    .Y(_2137_)
);

NOR2X1 _13791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1976_),
    .B(_2137_),
    .Y(_2138_)
);

INVX1 _13792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2131_),
    .Y(_2139_)
);

OAI21X1 _13793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2137_),
    .B(_2019_),
    .C(_2139_),
    .Y(_2140_)
);

AOI21X1 _13794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2138_),
    .B(_1807_),
    .C(_2140_),
    .Y(_2141_)
);

AOI21X1 _13795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2136_),
    .B(_2141_),
    .C(_2702_),
    .Y(_2142_)
);

NAND2X1 _13796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2134_),
    .B(_2142_),
    .Y(_2143_)
);

NOR2X1 _13797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [23]),
    .B(_1695_),
    .Y(_2144_)
);

AOI21X1 _13798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2096_),
    .B(_1727_),
    .C(_2144_),
    .Y(_2145_)
);

OAI21X1 _13799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2064_),
    .B(_1792_),
    .C(_2145_),
    .Y(_2147_)
);

AOI21X1 _13800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1899_),
    .B(_1987_),
    .C(_2147_),
    .Y(_2148_)
);

OAI21X1 _13801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1823_),
    .B(_2124_),
    .C(_2148_),
    .Y(_2149_)
);

AOI21X1 _13802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2136_),
    .B(_2149_),
    .C(_2798_),
    .Y(_2150_)
);

OAI21X1 _13803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2136_),
    .B(_2149_),
    .C(_2150_),
    .Y(_2151_)
);

NOR2X1 _13804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2676_),
    .B(_3132_),
    .Y(_2152_)
);

MUX2X1 _13805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1695_),
    .B(_2810_),
    .S(\datapath.alu.b_0_bF$buf0 ),
    .Y(_2153_)
);

MUX2X1 _13806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2153_),
    .B(_2081_),
    .S(_2489__bF$buf7),
    .Y(_2154_)
);

NAND2X1 _13807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf5 ),
    .B(_2004_),
    .Y(_2155_)
);

OAI21X1 _13808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf4 ),
    .B(_2154_),
    .C(_2155_),
    .Y(_2156_)
);

NAND3X1 _13809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf3 ),
    .B(_1841_),
    .C(_1837_),
    .Y(_2158_)
);

OAI21X1 _13810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2156_),
    .B(\datapath.alu.b_3_bF$buf2 ),
    .C(_2158_),
    .Y(_2159_)
);

NOR2X1 _13811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884_),
    .B(_2159_),
    .Y(_2160_)
);

INVX1 _13812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .Y(_2161_)
);

AOI21X1 _13813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [24]),
    .B(_2865__bF$buf1),
    .C(_2869__bF$buf0),
    .Y(_2162_)
);

AOI21X1 _13814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2438_),
    .B(_3114_),
    .C(_3113_),
    .Y(_2163_)
);

OAI21X1 _13815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2162_),
    .B(_2810_),
    .C(_2163_),
    .Y(_2164_)
);

AOI21X1 _13816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2810_),
    .B(_2706__bF$buf1),
    .C(_2802_),
    .Y(_2165_)
);

OAI21X1 _13817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2561_),
    .B(_2165_),
    .C(_1826_),
    .Y(_2166_)
);

AOI21X1 _13818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2161_),
    .B(_2164_),
    .C(_2166_),
    .Y(_2167_)
);

OAI21X1 _13819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3160_),
    .B(_1894_),
    .C(_2167_),
    .Y(_2169_)
);

OR2X2 _13820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2160_),
    .B(_2169_),
    .Y(_2170_)
);

AOI21X1 _13821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf0),
    .B(_2152_),
    .C(_2170_),
    .Y(_2171_)
);

NAND3X1 _13822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2171_),
    .B(_2151_),
    .C(_2143_),
    .Y(\datapath.alu.c [24])
);

AOI21X1 _13823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2125_),
    .B(_2133_),
    .C(_2439_),
    .Y(_2172_)
);

OR2X2 _13824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2172_),
    .B(_2436_),
    .Y(_2173_)
);

AOI21X1 _13825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2436_),
    .B(_2172_),
    .C(_2702_),
    .Y(_2174_)
);

INVX1 _13826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2436_),
    .Y(_2175_)
);

OAI21X1 _13827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2810_),
    .B(\datapath.alu.b [24]),
    .C(_2175_),
    .Y(_2176_)
);

AOI21X1 _13828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2136_),
    .B(_2149_),
    .C(_2176_),
    .Y(_2177_)
);

NAND2X1 _13829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1899_),
    .B(_1987_),
    .Y(_2179_)
);

OR2X2 _13830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2064_),
    .B(_1792_),
    .Y(_2180_)
);

NAND3X1 _13831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2179_),
    .B(_2145_),
    .C(_2180_),
    .Y(_2181_)
);

AOI21X1 _13832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2583_),
    .B(_1817_),
    .C(_2181_),
    .Y(_2182_)
);

NOR2X1 _13833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [24]),
    .B(_2810_),
    .Y(_2183_)
);

AOI21X1 _13834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2436_),
    .B(_2183_),
    .C(_2798_),
    .Y(_2184_)
);

OAI21X1 _13835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2182_),
    .B(_2440_),
    .C(_2184_),
    .Y(_2185_)
);

AOI22X1 _13836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560_),
    .B(_2706__bF$buf0),
    .C(_2802_),
    .D(\datapath.alu.b [25]),
    .Y(_2186_)
);

OAI21X1 _13837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2433_),
    .B(_2694_),
    .C(_2186_),
    .Y(_2187_)
);

OAI22X1 _13838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2436_),
    .B(_2688__bF$buf0),
    .C(_2692_),
    .D(_2432_),
    .Y(_2188_)
);

INVX2 _13839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2435_),
    .Y(_2190_)
);

OAI21X1 _13840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2190_),
    .B(_2680__bF$buf3),
    .C(_1826_),
    .Y(_2191_)
);

OR2X2 _13841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2191_),
    .B(_2188_),
    .Y(_2192_)
);

NOR2X1 _13842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2187_),
    .B(_2192_),
    .Y(_2193_)
);

OAI21X1 _13843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3183_),
    .B(_1894_),
    .C(_2193_),
    .Y(_2194_)
);

NAND2X1 _13844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf10 ),
    .B(_2810_),
    .Y(_2195_)
);

OAI21X1 _13845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf9 ),
    .B(\datapath.alu.a [25]),
    .C(_2195_),
    .Y(_2196_)
);

NAND2X1 _13846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf6),
    .B(_2196_),
    .Y(_2197_)
);

OAI21X1 _13847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf5),
    .B(_2102_),
    .C(_2197_),
    .Y(_2198_)
);

NOR2X1 _13848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf3 ),
    .B(_2198_),
    .Y(_2199_)
);

OAI21X1 _13849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2035_),
    .B(_2495__bF$buf2),
    .C(_2497__bF$buf0),
    .Y(_2201_)
);

OAI22X1 _13850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2201_),
    .B(_2199_),
    .C(_2497__bF$buf6),
    .D(_1881_),
    .Y(_2202_)
);

OAI21X1 _13851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2700_),
    .B(_2202_),
    .C(_3177_),
    .Y(_2203_)
);

AOI21X1 _13852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf5),
    .B(_2203_),
    .C(_2194_),
    .Y(_2204_)
);

OAI21X1 _13853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2177_),
    .B(_2185_),
    .C(_2204_),
    .Y(_2205_)
);

AOI21X1 _13854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2174_),
    .B(_2173_),
    .C(_2205_),
    .Y(_2206_)
);

INVX2 _13855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2206_),
    .Y(\datapath.alu.c [25])
);

INVX2 _13856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2430_),
    .Y(_2207_)
);

NOR2X1 _13857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2436_),
    .B(_2136_),
    .Y(_2208_)
);

INVX1 _13858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2208_),
    .Y(_2209_)
);

OAI21X1 _13859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2190_),
    .B(_2438_),
    .C(_2432_),
    .Y(_2211_)
);

INVX1 _13860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2211_),
    .Y(_2212_)
);

OAI21X1 _13861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2141_),
    .B(_2209_),
    .C(_2212_),
    .Y(_2213_)
);

AND2X2 _13862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2213_),
    .B(_2207_),
    .Y(_2214_)
);

OAI21X1 _13863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2213_),
    .B(_2207_),
    .C(_2703__bF$buf1),
    .Y(_2215_)
);

INVX1 _13864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2432_),
    .Y(_2216_)
);

OAI21X1 _13865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2190_),
    .B(_2216_),
    .C(_2183_),
    .Y(_2217_)
);

OAI21X1 _13866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2433_),
    .B(\datapath.alu.b [25]),
    .C(_2217_),
    .Y(_2218_)
);

INVX1 _13867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2218_),
    .Y(_2219_)
);

OAI21X1 _13868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2182_),
    .B(_2440_),
    .C(_2219_),
    .Y(_2220_)
);

OR2X2 _13869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2220_),
    .B(_2430_),
    .Y(_2222_)
);

AOI21X1 _13870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2430_),
    .B(_2220_),
    .C(_2798_),
    .Y(_2223_)
);

NAND2X1 _13871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf4),
    .B(_3222_),
    .Y(_2224_)
);

NAND2X1 _13872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf0 ),
    .B(_2153_),
    .Y(_2225_)
);

NAND2X1 _13873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf8 ),
    .B(_2433_),
    .Y(_2226_)
);

OAI21X1 _13874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf7 ),
    .B(\datapath.alu.a [26]),
    .C(_2226_),
    .Y(_2227_)
);

OAI21X1 _13875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2227_),
    .B(\datapath.alu.b_1_bF$buf6 ),
    .C(_2225_),
    .Y(_2228_)
);

MUX2X1 _13876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2228_),
    .B(_2084_),
    .S(_2495__bF$buf1),
    .Y(_2229_)
);

NOR2X1 _13877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf1 ),
    .B(_2229_),
    .Y(_2230_)
);

NOR2X1 _13878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf5),
    .B(_1926_),
    .Y(_2231_)
);

OAI21X1 _13879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2231_),
    .B(_2230_),
    .C(_2701_),
    .Y(_2233_)
);

AOI21X1 _13880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3234_),
    .B(_3240_),
    .C(_1894_),
    .Y(_2234_)
);

OAI21X1 _13881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2707_),
    .B(\datapath.alu.a [26]),
    .C(_2708__bF$buf0),
    .Y(_2235_)
);

AOI22X1 _13882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [26]),
    .B(_2869__bF$buf3),
    .C(_2235_),
    .D(\datapath.alu.b [26]),
    .Y(_2236_)
);

INVX1 _13883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2424_),
    .Y(_2237_)
);

AOI22X1 _13884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2237_),
    .B(_2865__bF$buf0),
    .C(_2207_),
    .D(_3114_),
    .Y(_2238_)
);

AOI21X1 _13885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2413_),
    .B(_3113_),
    .C(_2045_),
    .Y(_2239_)
);

NAND3X1 _13886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2236_),
    .B(_2238_),
    .C(_2239_),
    .Y(_2240_)
);

NOR2X1 _13887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2234_),
    .B(_2240_),
    .Y(_2241_)
);

NAND3X1 _13888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2224_),
    .B(_2233_),
    .C(_2241_),
    .Y(_2242_)
);

AOI21X1 _13889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2223_),
    .B(_2222_),
    .C(_2242_),
    .Y(_2244_)
);

OAI21X1 _13890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2214_),
    .B(_2215_),
    .C(_2244_),
    .Y(\datapath.alu.c [26])
);

OAI21X1 _13891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2214_),
    .B(_2237_),
    .C(_2381_),
    .Y(_2245_)
);

INVX2 _13892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2381_),
    .Y(_2246_)
);

NAND2X1 _13893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2207_),
    .B(_2213_),
    .Y(_2247_)
);

NAND3X1 _13894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2246_),
    .B(_2424_),
    .C(_2247_),
    .Y(_2248_)
);

AOI21X1 _13895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2248_),
    .B(_2245_),
    .C(_2702_),
    .Y(_2249_)
);

NOR2X1 _13896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [26]),
    .B(_2392_),
    .Y(_2250_)
);

AOI21X1 _13897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2430_),
    .B(_2220_),
    .C(_2250_),
    .Y(_2251_)
);

AND2X2 _13898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2251_),
    .B(_2246_),
    .Y(_2252_)
);

OAI21X1 _13899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2251_),
    .B(_2246_),
    .C(_2799__bF$buf1),
    .Y(_2254_)
);

NOR2X1 _13900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf4),
    .B(_1961_),
    .Y(_2255_)
);

NAND2X1 _13901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf6 ),
    .B(_2392_),
    .Y(_2256_)
);

OAI21X1 _13902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf5 ),
    .B(\datapath.alu.a [27]),
    .C(_2256_),
    .Y(_2257_)
);

MUX2X1 _13903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2257_),
    .B(_2196_),
    .S(_2489__bF$buf4),
    .Y(_2258_)
);

MUX2X1 _13904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2258_),
    .B(_2105_),
    .S(_2495__bF$buf0),
    .Y(_2259_)
);

NOR2X1 _13905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf0 ),
    .B(_2259_),
    .Y(_2260_)
);

OAI21X1 _13906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2260_),
    .B(_2255_),
    .C(_2701_),
    .Y(_2261_)
);

NAND2X1 _13907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1893_),
    .B(_1618_),
    .Y(_2262_)
);

AOI21X1 _13908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [27]),
    .B(_2865__bF$buf3),
    .C(_2869__bF$buf2),
    .Y(_2263_)
);

AOI21X1 _13909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2339_),
    .B(_3114_),
    .C(_3113_),
    .Y(_2265_)
);

OAI21X1 _13910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2263_),
    .B(_2349_),
    .C(_2265_),
    .Y(_2266_)
);

AOI21X1 _13911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2349_),
    .B(_2706__bF$buf3),
    .C(_2802_),
    .Y(_2267_)
);

OAI21X1 _13912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2360_),
    .B(_2267_),
    .C(_1826_),
    .Y(_2268_)
);

AOI21X1 _13913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2371_),
    .B(_2266_),
    .C(_2268_),
    .Y(_2269_)
);

NAND3X1 _13914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2261_),
    .B(_2269_),
    .C(_2262_),
    .Y(_2270_)
);

AOI21X1 _13915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf3),
    .B(_1610_),
    .C(_2270_),
    .Y(_2271_)
);

OAI21X1 _13916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2252_),
    .B(_2254_),
    .C(_2271_),
    .Y(_2272_)
);

OR2X2 _13917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2249_),
    .B(_2272_),
    .Y(\datapath.alu.c [27])
);

NOR2X1 _13918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2381_),
    .B(_2430_),
    .Y(_2273_)
);

INVX1 _13919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2273_),
    .Y(_2275_)
);

NOR2X1 _13920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2275_),
    .B(_2209_),
    .Y(_2276_)
);

OAI21X1 _13921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2381_),
    .B(_2424_),
    .C(_2339_),
    .Y(_2277_)
);

AOI21X1 _13922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2211_),
    .B(_2273_),
    .C(_2277_),
    .Y(_2278_)
);

INVX1 _13923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2278_),
    .Y(_2279_)
);

AOI21X1 _13924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2276_),
    .B(_2133_),
    .C(_2279_),
    .Y(_2280_)
);

AOI21X1 _13925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2307_),
    .B(_2280_),
    .C(_2702_),
    .Y(_2281_)
);

OAI21X1 _13926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2307_),
    .B(_2280_),
    .C(_2281_),
    .Y(_2282_)
);

INVX1 _13927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2441_),
    .Y(_2283_)
);

INVX1 _13928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2431_),
    .Y(_2284_)
);

INVX1 _13929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2250_),
    .Y(_2286_)
);

OAI21X1 _13930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2286_),
    .B(_2567_),
    .C(_2565_),
    .Y(_2287_)
);

AOI21X1 _13931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2284_),
    .B(_2218_),
    .C(_2287_),
    .Y(_2288_)
);

OAI21X1 _13932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2182_),
    .B(_2283_),
    .C(_2288_),
    .Y(_2289_)
);

AOI21X1 _13933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2307_),
    .B(_2289_),
    .C(_2798_),
    .Y(_2290_)
);

OAI21X1 _13934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2307_),
    .B(_2289_),
    .C(_2290_),
    .Y(_2291_)
);

OR2X2 _13935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1655_),
    .B(_1656_),
    .Y(_2292_)
);

OAI21X1 _13936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2707_),
    .B(\datapath.alu.a [28]),
    .C(_2708__bF$buf3),
    .Y(_2293_)
);

INVX1 _13937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2307_),
    .Y(_2294_)
);

AOI22X1 _13938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [28]),
    .B(_2869__bF$buf1),
    .C(_2294_),
    .D(_3114_),
    .Y(_2295_)
);

INVX1 _13939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2296_),
    .Y(_2297_)
);

AOI22X1 _13940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2865__bF$buf2),
    .B(_2297_),
    .C(_2285_),
    .D(_3113_),
    .Y(_2298_)
);

NAND3X1 _13941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2295_),
    .B(_2298_),
    .C(_1826_),
    .Y(_2299_)
);

AOI21X1 _13942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [28]),
    .B(_2293_),
    .C(_2299_),
    .Y(_2300_)
);

MUX2X1 _13943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2349_),
    .B(_2264_),
    .S(\datapath.alu.b_0_bF$buf4 ),
    .Y(_2301_)
);

NAND2X1 _13944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf3),
    .B(_2301_),
    .Y(_2302_)
);

OAI21X1 _13945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2227_),
    .B(_2489__bF$buf2),
    .C(_2302_),
    .Y(_2303_)
);

NAND2X1 _13946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495__bF$buf6),
    .B(_2303_),
    .Y(_2304_)
);

OAI21X1 _13947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495__bF$buf5),
    .B(_2154_),
    .C(_2304_),
    .Y(_2305_)
);

OAI21X1 _13948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2008_),
    .B(_2497__bF$buf3),
    .C(_2480__bF$buf2),
    .Y(_2306_)
);

AOI21X1 _13949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf2),
    .B(_2305_),
    .C(_2306_),
    .Y(_2308_)
);

NOR2X1 _13950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2701_),
    .B(_1671_),
    .Y(_2309_)
);

OAI21X1 _13951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2308_),
    .B(_2309_),
    .C(_2300_),
    .Y(_2310_)
);

AOI21X1 _13952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf1),
    .B(_2292_),
    .C(_2310_),
    .Y(_2311_)
);

NAND3X1 _13953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2291_),
    .B(_2311_),
    .C(_2282_),
    .Y(\datapath.alu.c [28])
);

NAND2X1 _13954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2200_),
    .B(_2243_),
    .Y(_2312_)
);

INVX1 _13955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2276_),
    .Y(_2313_)
);

OAI21X1 _13956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2141_),
    .B(_2313_),
    .C(_2278_),
    .Y(_2314_)
);

NAND2X1 _13957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2294_),
    .B(_2314_),
    .Y(_2315_)
);

AOI21X1 _13958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2296_),
    .B(_2315_),
    .C(_2312_),
    .Y(_2316_)
);

INVX2 _13959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2312_),
    .Y(_2318_)
);

OAI21X1 _13960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2280_),
    .B(_2307_),
    .C(_2296_),
    .Y(_2319_)
);

OAI21X1 _13961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2319_),
    .B(_2318_),
    .C(_2703__bF$buf0),
    .Y(_2320_)
);

NAND2X1 _13962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2307_),
    .B(_2289_),
    .Y(_2321_)
);

NOR2X1 _13963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [28]),
    .B(_2264_),
    .Y(_2322_)
);

NOR2X1 _13964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2322_),
    .B(_2312_),
    .Y(_2323_)
);

NAND2X1 _13965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2323_),
    .B(_2321_),
    .Y(_2324_)
);

INVX1 _13966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2317_),
    .Y(_2325_)
);

INVX1 _13967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2322_),
    .Y(_2326_)
);

OAI21X1 _13968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2318_),
    .B(_2326_),
    .C(_2799__bF$buf0),
    .Y(_2327_)
);

AOI21X1 _13969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2325_),
    .B(_2289_),
    .C(_2327_),
    .Y(_2329_)
);

AOI22X1 _13970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2571_),
    .B(_2706__bF$buf2),
    .C(_2802_),
    .D(\datapath.alu.b [29]),
    .Y(_2330_)
);

OAI22X1 _13971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2312_),
    .B(_2688__bF$buf3),
    .C(_2692_),
    .D(_2200_),
    .Y(_2331_)
);

OAI22X1 _13972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2221_),
    .B(_2694_),
    .C(_2680__bF$buf2),
    .D(_2253_),
    .Y(_2332_)
);

NOR2X1 _13973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2331_),
    .B(_2332_),
    .Y(_2333_)
);

NAND3X1 _13974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1826_),
    .B(_2330_),
    .C(_2333_),
    .Y(_2334_)
);

AOI21X1 _13975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480__bF$buf0),
    .B(_1698_),
    .C(_2334_),
    .Y(_2335_)
);

OAI21X1 _13976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2221_),
    .B(\datapath.alu.b_0_bF$buf3 ),
    .C(_2730_),
    .Y(_2336_)
);

NAND2X1 _13977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf5 ),
    .B(_2257_),
    .Y(_2337_)
);

OAI21X1 _13978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_1_bF$buf4 ),
    .B(_2336_),
    .C(_2337_),
    .Y(_2338_)
);

MUX2X1 _13979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2198_),
    .B(_2338_),
    .S(\datapath.alu.b_2_bF$buf2 ),
    .Y(_2340_)
);

NAND2X1 _13980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf1),
    .B(_2340_),
    .Y(_2341_)
);

NAND2X1 _13981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf6 ),
    .B(_2036_),
    .Y(_2342_)
);

NAND2X1 _13982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2342_),
    .B(_2341_),
    .Y(_2343_)
);

NAND2X1 _13983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_4_bF$buf1 ),
    .B(_1718_),
    .Y(_2344_)
);

OAI21X1 _13984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2343_),
    .B(\datapath.alu.b_4_bF$buf0 ),
    .C(_2344_),
    .Y(_2345_)
);

OAI21X1 _13985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2345_),
    .B(_2700_),
    .C(_2335_),
    .Y(_2346_)
);

AOI21X1 _13986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2329_),
    .B(_2324_),
    .C(_2346_),
    .Y(_2347_)
);

OAI21X1 _13987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2320_),
    .B(_2316_),
    .C(_2347_),
    .Y(\datapath.alu.c [29])
);

INVX4 _13988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2178_),
    .Y(_2348_)
);

OAI21X1 _13989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2253_),
    .B(_2296_),
    .C(_2200_),
    .Y(_2350_)
);

NOR2X1 _13990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2312_),
    .B(_2307_),
    .Y(_2351_)
);

AOI21X1 _13991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2351_),
    .B(_2314_),
    .C(_2350_),
    .Y(_2352_)
);

NAND2X1 _13992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2348_),
    .B(_2352_),
    .Y(_2353_)
);

OR2X2 _13993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2352_),
    .B(_2348_),
    .Y(_2354_)
);

AOI21X1 _13994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2353_),
    .B(_2354_),
    .C(_2702_),
    .Y(_2355_)
);

OAI21X1 _13995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2318_),
    .B(_2326_),
    .C(_2570_),
    .Y(_2356_)
);

AOI21X1 _13996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2325_),
    .B(_2289_),
    .C(_2356_),
    .Y(_2357_)
);

AND2X2 _13997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2357_),
    .B(_2348_),
    .Y(_2358_)
);

OAI21X1 _13998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2357_),
    .B(_2348_),
    .C(_2799__bF$buf3),
    .Y(_2359_)
);

OAI21X1 _13999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2707_),
    .B(\datapath.alu.a [30]),
    .C(_2708__bF$buf2),
    .Y(_2361_)
);

AOI22X1 _14000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [30]),
    .B(_2869__bF$buf0),
    .C(_2348_),
    .D(_3114_),
    .Y(_2362_)
);

INVX1 _14001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2168_),
    .Y(_2363_)
);

AOI22X1 _14002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2865__bF$buf1),
    .B(_2363_),
    .C(_2157_),
    .D(_3113_),
    .Y(_2364_)
);

NAND3X1 _14003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362_),
    .B(_2364_),
    .C(_1826_),
    .Y(_2365_)
);

AOI21X1 _14004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b [30]),
    .B(_2361_),
    .C(_2365_),
    .Y(_2366_)
);

OAI21X1 _14005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1754_),
    .B(\datapath.alu.b_4_bF$buf4 ),
    .C(_2366_),
    .Y(_2367_)
);

NOR2X1 _14006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_0_bF$buf2 ),
    .B(\datapath.alu.a [30]),
    .Y(_2368_)
);

NOR2X1 _14007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [29]),
    .B(_2491_),
    .Y(_2369_)
);

OAI21X1 _14008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2369_),
    .B(_2368_),
    .C(_2489__bF$buf1),
    .Y(_2370_)
);

OAI21X1 _14009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf0),
    .B(_2301_),
    .C(_2370_),
    .Y(_2372_)
);

NAND2X1 _14010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf1 ),
    .B(_2228_),
    .Y(_2373_)
);

OAI21X1 _14011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2372_),
    .B(\datapath.alu.b_2_bF$buf0 ),
    .C(_2373_),
    .Y(_2374_)
);

NAND2X1 _14012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf5 ),
    .B(_2085_),
    .Y(_2375_)
);

OAI21X1 _14013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_3_bF$buf4 ),
    .B(_2374_),
    .C(_2375_),
    .Y(_2376_)
);

AOI22X1 _14014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376_),
    .B(_2480__bF$buf5),
    .C(_1745_),
    .D(_2884_),
    .Y(_2377_)
);

NOR2X1 _14015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2377_),
    .B(_2367_),
    .Y(_2378_)
);

OAI21X1 _14016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2358_),
    .B(_2359_),
    .C(_2378_),
    .Y(_2379_)
);

NOR2X1 _14017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2379_),
    .B(_2355_),
    .Y(_2380_)
);

INVX2 _14018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2380_),
    .Y(\datapath.alu.c [30])
);

INVX2 _14019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2574_),
    .Y(_2382_)
);

OAI21X1 _14020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2352_),
    .B(_2178_),
    .C(_2168_),
    .Y(_2383_)
);

AND2X2 _14021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2383_),
    .B(_2382_),
    .Y(_2384_)
);

OAI21X1 _14022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2383_),
    .B(_2382_),
    .C(_2703__bF$buf3),
    .Y(_2385_)
);

NAND2X1 _14023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.a [30]),
    .B(_2146_),
    .Y(_2386_)
);

OAI21X1 _14024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2357_),
    .B(_2348_),
    .C(_2386_),
    .Y(_2387_)
);

XNOR2X1 _14025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2387_),
    .B(_2382_),
    .Y(_2388_)
);

AND2X2 _14026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2915_),
    .B(_2736_),
    .Y(_2389_)
);

NAND2X1 _14027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf7),
    .B(_2389_),
    .Y(_2390_)
);

OAI21X1 _14028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489__bF$buf6),
    .B(_2336_),
    .C(_2390_),
    .Y(_2391_)
);

AOI21X1 _14029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf7 ),
    .B(_2258_),
    .C(\datapath.alu.b_3_bF$buf3 ),
    .Y(_2393_)
);

OAI21X1 _14030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.b_2_bF$buf6 ),
    .B(_2391_),
    .C(_2393_),
    .Y(_2394_)
);

OAI21X1 _14031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497__bF$buf0),
    .B(_2107_),
    .C(_2394_),
    .Y(_2395_)
);

NAND2X1 _14032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1893_),
    .B(_1783_),
    .Y(_2396_)
);

AOI21X1 _14033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1620_),
    .B(_3114_),
    .C(_3113_),
    .Y(_2397_)
);

NAND2X1 _14034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1630_),
    .B(_2865__bF$buf0),
    .Y(_2398_)
);

OAI21X1 _14035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1652_),
    .B(_2708__bF$buf1),
    .C(_2398_),
    .Y(_2399_)
);

AOI21X1 _14036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2575_),
    .B(_2706__bF$buf1),
    .C(_2399_),
    .Y(_2400_)
);

OAI21X1 _14037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1674_),
    .B(_2397_),
    .C(_2400_),
    .Y(_2401_)
);

OAI21X1 _14038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2869__bF$buf3),
    .B(_2717_),
    .C(\datapath.alu.a [31]),
    .Y(_2402_)
);

NAND2X1 _14039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686_),
    .B(_3015_),
    .Y(_2404_)
);

OAI21X1 _14040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2404_),
    .B(_1786_),
    .C(_2402_),
    .Y(_2405_)
);

NOR2X1 _14041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2405_),
    .B(_2401_),
    .Y(_2406_)
);

AND2X2 _14042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2406_),
    .B(_2396_),
    .Y(_2407_)
);

OAI21X1 _14043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884_),
    .B(_2395_),
    .C(_2407_),
    .Y(_2408_)
);

AOI21X1 _14044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2799__bF$buf2),
    .B(_2388_),
    .C(_2408_),
    .Y(_2409_)
);

OAI21X1 _14045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2384_),
    .B(_2385_),
    .C(_2409_),
    .Y(\datapath.alu.c [31])
);

NOR3X1 _14046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2249_),
    .B(_2272_),
    .C(\datapath.alu.c [29]),
    .Y(_2410_)
);

NAND3X1 _14047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2091_),
    .B(_2063_),
    .C(_2206_),
    .Y(_2411_)
);

NOR3X1 _14048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [26]),
    .B(\datapath.alu.c [28]),
    .C(_2411_),
    .Y(_2412_)
);

NOR2X1 _14049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [5]),
    .B(\datapath.alu.c [8]),
    .Y(_2414_)
);

NAND3X1 _14050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2714_),
    .B(_3073_),
    .C(_2414_),
    .Y(_2415_)
);

NOR3X1 _14051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [2]),
    .B(\datapath.alu.c [4]),
    .C(\datapath.alu.c [3]),
    .Y(_2416_)
);

NAND3X1 _14052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2807_),
    .B(_3122_),
    .C(_2416_),
    .Y(_2417_)
);

NOR2X1 _14053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2415_),
    .B(_2417_),
    .Y(_2418_)
);

NAND3X1 _14054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1855_),
    .B(_1593_),
    .C(_1682_),
    .Y(_2419_)
);

NOR2X1 _14055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [9]),
    .B(_2419_),
    .Y(_2420_)
);

NAND3X1 _14056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1722_),
    .B(_2420_),
    .C(_2418_),
    .Y(_2421_)
);

NOR2X1 _14057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [20]),
    .B(\datapath.alu.c [24]),
    .Y(_2422_)
);

NAND3X1 _14058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1935_),
    .B(_2054_),
    .C(_2422_),
    .Y(_2423_)
);

NOR2X1 _14059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2423_),
    .B(_2421_),
    .Y(_2425_)
);

NAND3X1 _14060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2410_),
    .B(_2412_),
    .C(_2425_),
    .Y(_2426_)
);

NAND3X1 _14061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1766_),
    .B(_1629_),
    .C(_1898_),
    .Y(_2427_)
);

NOR3X1 _14062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [15]),
    .B(\datapath.alu.c [19]),
    .C(_2427_),
    .Y(_2428_)
);

NAND3X1 _14063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2123_),
    .B(_2380_),
    .C(_2428_),
    .Y(_2429_)
);

NOR3X1 _14064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.alu.c [31]),
    .B(_2429_),
    .C(_2426_),
    .Y(\datapath.alu.z )
);

INVX2 _14065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [0]),
    .Y(_3247_)
);

INVX1 _14066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [21]),
    .Y(_3248_)
);

NAND2X1 _14067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [20]),
    .B(_3248_),
    .Y(_3249_)
);

INVX8 _14068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret_bF$buf3 ),
    .Y(_3250_)
);

NAND2X1 _14069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.allowcsrwrite ),
    .B(_3250__bF$buf5),
    .Y(_3251_)
);

NOR2X1 _14070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3249_),
    .B(_3251_),
    .Y(_3252_)
);

INVX1 _14071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [30]),
    .Y(_3253_)
);

INVX1 _14072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [27]),
    .Y(_3254_)
);

AND2X2 _14073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3254_),
    .B(\datapath.meminstr [29]),
    .Y(_3255_)
);

INVX1 _14074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [28]),
    .Y(_3256_)
);

NOR2X1 _14075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [31]),
    .B(_3256_),
    .Y(_3257_)
);

NAND3X1 _14076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3253_),
    .B(_3257_),
    .C(_3255_),
    .Y(_3258_)
);

INVX1 _14077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [26]),
    .Y(_3259_)
);

NOR2X1 _14078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [25]),
    .B(\datapath.meminstr [24]),
    .Y(_3260_)
);

NAND2X1 _14079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3259_),
    .B(_3260_),
    .Y(_3261_)
);

NOR2X1 _14080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3261_),
    .B(_3258_),
    .Y(_3262_)
);

INVX1 _14081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [23]),
    .Y(_3263_)
);

NAND2X1 _14082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [22]),
    .B(_3263_),
    .Y(_3264_)
);

NOR2X1 _14083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf7 ),
    .B(_3264_),
    .Y(_3265_)
);

AND2X2 _14084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3262_),
    .B(_3265_),
    .Y(_3266_)
);

NAND2X1 _14085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3252_),
    .B(_3266_),
    .Y(_3267_)
);

NOR2X1 _14086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__0_bF$buf0),
    .B(_3267__bF$buf6),
    .Y(_3268_)
);

AOI21X1 _14087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3247_),
    .B(_3267__bF$buf5),
    .C(_3268_),
    .Y(\datapath.csr._13_ [0])
);

INVX1 _14088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [1]),
    .Y(_3269_)
);

NOR2X1 _14089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf5),
    .B(_3267__bF$buf4),
    .Y(_3270_)
);

AOI21X1 _14090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3269_),
    .B(_3267__bF$buf3),
    .C(_3270_),
    .Y(\datapath.csr._13_ [1])
);

INVX1 _14091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [2]),
    .Y(_3271_)
);

NOR2X1 _14092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[2]),
    .B(_3267__bF$buf2),
    .Y(_3272_)
);

AOI21X1 _14093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3271_),
    .B(_3267__bF$buf1),
    .C(_3272_),
    .Y(\datapath.csr._13_ [2])
);

INVX2 _14094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [3]),
    .Y(_3273_)
);

NOR2X1 _14095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[3]),
    .B(_3267__bF$buf0),
    .Y(_3274_)
);

AOI21X1 _14096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3273_),
    .B(_3267__bF$buf6),
    .C(_3274_),
    .Y(\datapath.csr._13_ [3])
);

INVX2 _14097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [4]),
    .Y(_3275_)
);

NOR2X1 _14098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[4]),
    .B(_3267__bF$buf5),
    .Y(_3276_)
);

AOI21X1 _14099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3275_),
    .B(_3267__bF$buf4),
    .C(_3276_),
    .Y(\datapath.csr._13_ [4])
);

INVX2 _14100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [5]),
    .Y(_3277_)
);

NOR2X1 _14101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[5]),
    .B(_3267__bF$buf3),
    .Y(_3278_)
);

AOI21X1 _14102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3277_),
    .B(_3267__bF$buf2),
    .C(_3278_),
    .Y(\datapath.csr._13_ [5])
);

INVX2 _14103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [6]),
    .Y(_3279_)
);

NOR2X1 _14104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[6]),
    .B(_3267__bF$buf1),
    .Y(_3280_)
);

AOI21X1 _14105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3279_),
    .B(_3267__bF$buf0),
    .C(_3280_),
    .Y(\datapath.csr._13_ [6])
);

INVX1 _14106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [7]),
    .Y(_3281_)
);

NOR2X1 _14107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[7]),
    .B(_3267__bF$buf6),
    .Y(_3282_)
);

AOI21X1 _14108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3281_),
    .B(_3267__bF$buf5),
    .C(_3282_),
    .Y(\datapath.csr._13_ [7])
);

INVX1 _14109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [8]),
    .Y(_3283_)
);

NOR2X1 _14110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[8]),
    .B(_3267__bF$buf4),
    .Y(_3284_)
);

AOI21X1 _14111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3283_),
    .B(_3267__bF$buf3),
    .C(_3284_),
    .Y(\datapath.csr._13_ [8])
);

INVX1 _14112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [9]),
    .Y(_3285_)
);

NOR2X1 _14113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[9]),
    .B(_3267__bF$buf2),
    .Y(_3286_)
);

AOI21X1 _14114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3285_),
    .B(_3267__bF$buf1),
    .C(_3286_),
    .Y(\datapath.csr._13_ [9])
);

INVX2 _14115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [10]),
    .Y(_3287_)
);

NOR2X1 _14116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[10]),
    .B(_3267__bF$buf0),
    .Y(_3288_)
);

AOI21X1 _14117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3287_),
    .B(_3267__bF$buf6),
    .C(_3288_),
    .Y(\datapath.csr._13_ [10])
);

INVX1 _14118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[11]),
    .Y(_3289_)
);

INVX1 _14119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [11]),
    .Y(_3290_)
);

MUX2X1 _14120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3290_),
    .B(_3289_),
    .S(_3267__bF$buf5),
    .Y(\datapath.csr._13_ [11])
);

INVX2 _14121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [12]),
    .Y(_3291_)
);

NOR2X1 _14122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[12]),
    .B(_3267__bF$buf4),
    .Y(_3292_)
);

AOI21X1 _14123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3291_),
    .B(_3267__bF$buf3),
    .C(_3292_),
    .Y(\datapath.csr._13_ [12])
);

INVX1 _14124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [13]),
    .Y(_3293_)
);

NOR2X1 _14125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[13]),
    .B(_3267__bF$buf2),
    .Y(_3294_)
);

AOI21X1 _14126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3293_),
    .B(_3267__bF$buf1),
    .C(_3294_),
    .Y(\datapath.csr._13_ [13])
);

INVX2 _14127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [14]),
    .Y(_3295_)
);

NOR2X1 _14128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[14]),
    .B(_3267__bF$buf0),
    .Y(_3296_)
);

AOI21X1 _14129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3295_),
    .B(_3267__bF$buf6),
    .C(_3296_),
    .Y(\datapath.csr._13_ [14])
);

INVX1 _14130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [15]),
    .Y(_3297_)
);

NOR2X1 _14131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[15]),
    .B(_3267__bF$buf5),
    .Y(_3298_)
);

AOI21X1 _14132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3297_),
    .B(_3267__bF$buf4),
    .C(_3298_),
    .Y(\datapath.csr._13_ [15])
);

INVX1 _14133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [16]),
    .Y(_3299_)
);

NOR2X1 _14134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[16]),
    .B(_3267__bF$buf3),
    .Y(_3300_)
);

AOI21X1 _14135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3299_),
    .B(_3267__bF$buf2),
    .C(_3300_),
    .Y(\datapath.csr._13_ [16])
);

INVX1 _14136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [17]),
    .Y(_3301_)
);

NOR2X1 _14137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[17]),
    .B(_3267__bF$buf1),
    .Y(_3302_)
);

AOI21X1 _14138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3301_),
    .B(_3267__bF$buf0),
    .C(_3302_),
    .Y(\datapath.csr._13_ [17])
);

INVX1 _14139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [18]),
    .Y(_3303_)
);

NOR2X1 _14140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[18]),
    .B(_3267__bF$buf6),
    .Y(_3304_)
);

AOI21X1 _14141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3303_),
    .B(_3267__bF$buf5),
    .C(_3304_),
    .Y(\datapath.csr._13_ [18])
);

INVX1 _14142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [19]),
    .Y(_3305_)
);

NOR2X1 _14143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[19]),
    .B(_3267__bF$buf4),
    .Y(_3306_)
);

AOI21X1 _14144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3305_),
    .B(_3267__bF$buf3),
    .C(_3306_),
    .Y(\datapath.csr._13_ [19])
);

INVX2 _14145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [20]),
    .Y(_3307_)
);

NOR2X1 _14146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[20]),
    .B(_3267__bF$buf2),
    .Y(_3308_)
);

AOI21X1 _14147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3307_),
    .B(_3267__bF$buf1),
    .C(_3308_),
    .Y(\datapath.csr._13_ [20])
);

INVX1 _14148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [21]),
    .Y(_3309_)
);

NOR2X1 _14149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[21]),
    .B(_3267__bF$buf0),
    .Y(_3310_)
);

AOI21X1 _14150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3309_),
    .B(_3267__bF$buf6),
    .C(_3310_),
    .Y(\datapath.csr._13_ [21])
);

INVX1 _14151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [22]),
    .Y(_3311_)
);

NOR2X1 _14152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[22]),
    .B(_3267__bF$buf5),
    .Y(_3312_)
);

AOI21X1 _14153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3311_),
    .B(_3267__bF$buf4),
    .C(_3312_),
    .Y(\datapath.csr._13_ [22])
);

INVX1 _14154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [23]),
    .Y(_3313_)
);

NOR2X1 _14155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[23]),
    .B(_3267__bF$buf3),
    .Y(_3314_)
);

AOI21X1 _14156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3313_),
    .B(_3267__bF$buf2),
    .C(_3314_),
    .Y(\datapath.csr._13_ [23])
);

INVX1 _14157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [24]),
    .Y(_3315_)
);

NOR2X1 _14158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[24]),
    .B(_3267__bF$buf1),
    .Y(_3316_)
);

AOI21X1 _14159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3315_),
    .B(_3267__bF$buf0),
    .C(_3316_),
    .Y(\datapath.csr._13_ [24])
);

INVX1 _14160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [25]),
    .Y(_3317_)
);

NOR2X1 _14161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[25]),
    .B(_3267__bF$buf6),
    .Y(_3318_)
);

AOI21X1 _14162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3317_),
    .B(_3267__bF$buf5),
    .C(_3318_),
    .Y(\datapath.csr._13_ [25])
);

INVX1 _14163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [26]),
    .Y(_3319_)
);

NOR2X1 _14164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[26]),
    .B(_3267__bF$buf4),
    .Y(_3320_)
);

AOI21X1 _14165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3319_),
    .B(_3267__bF$buf3),
    .C(_3320_),
    .Y(\datapath.csr._13_ [26])
);

INVX1 _14166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [27]),
    .Y(_3321_)
);

NOR2X1 _14167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[27]),
    .B(_3267__bF$buf2),
    .Y(_3322_)
);

AOI21X1 _14168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3321_),
    .B(_3267__bF$buf1),
    .C(_3322_),
    .Y(\datapath.csr._13_ [27])
);

INVX1 _14169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [28]),
    .Y(_3323_)
);

NOR2X1 _14170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[28]),
    .B(_3267__bF$buf0),
    .Y(_3324_)
);

AOI21X1 _14171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3323_),
    .B(_3267__bF$buf6),
    .C(_3324_),
    .Y(\datapath.csr._13_ [28])
);

INVX1 _14172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [29]),
    .Y(_3325_)
);

NOR2X1 _14173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[29]),
    .B(_3267__bF$buf5),
    .Y(_3326_)
);

AOI21X1 _14174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3325_),
    .B(_3267__bF$buf4),
    .C(_3326_),
    .Y(\datapath.csr._13_ [29])
);

INVX1 _14175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [30]),
    .Y(_3327_)
);

NOR2X1 _14176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[30]),
    .B(_3267__bF$buf3),
    .Y(_3328_)
);

AOI21X1 _14177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3327_),
    .B(_3267__bF$buf2),
    .C(_3328_),
    .Y(\datapath.csr._13_ [30])
);

INVX1 _14178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [31]),
    .Y(_3329_)
);

NOR2X1 _14179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[31]),
    .B(_3267__bF$buf1),
    .Y(_3330_)
);

AOI21X1 _14180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3329_),
    .B(_3267__bF$buf0),
    .C(_3330_),
    .Y(\datapath.csr._13_ [31])
);

INVX1 _14181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [20]),
    .Y(_3331_)
);

NAND2X1 _14182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3248_),
    .B(_3331_),
    .Y(_3332_)
);

NOR2X1 _14183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3251_),
    .B(_3332_),
    .Y(_3333_)
);

NAND2X1 _14184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3333_),
    .B(_3266_),
    .Y(_3334_)
);

NAND2X1 _14185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mie ),
    .B(_3334_),
    .Y(_3335_)
);

OAI21X1 _14186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3289_),
    .B(_3334_),
    .C(_3335_),
    .Y(\datapath.csr._20_ )
);

NOR2X1 _14187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [23]),
    .B(\datapath.meminstr [22]),
    .Y(_3336_)
);

NAND3X1 _14188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [26]),
    .B(_3260_),
    .C(_3336_),
    .Y(_3337_)
);

NOR2X1 _14189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3337_),
    .B(_3258_),
    .Y(_3338_)
);

NAND2X1 _14190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3252_),
    .B(_3338_),
    .Y(_3339_)
);

INVX1 _14191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [0]),
    .Y(_3340_)
);

NAND2X1 _14192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3340_),
    .B(_3339__bF$buf6),
    .Y(_3341_)
);

OAI21X1 _14193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[2]),
    .B(_3339__bF$buf5),
    .C(_3341_),
    .Y(_3342_)
);

NAND2X1 _14194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf6 ),
    .B(\datapath.csr.csr_mepc [2]),
    .Y(_3343_)
);

OAI21X1 _14195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3342_),
    .B(\datapath.regcsrtrap_bF$buf5 ),
    .C(_3343_),
    .Y(\datapath.csr._26_ [0])
);

MUX2X1 _14196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [1]),
    .B(_0_[3]),
    .S(_3339__bF$buf4),
    .Y(_3344_)
);

NAND2X1 _14197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf4 ),
    .B(\datapath.csr.csr_mepc [3]),
    .Y(_3345_)
);

OAI21X1 _14198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3344_),
    .B(\datapath.regcsrtrap_bF$buf3 ),
    .C(_3345_),
    .Y(\datapath.csr._26_ [1])
);

MUX2X1 _14199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [2]),
    .B(_0_[4]),
    .S(_3339__bF$buf3),
    .Y(_3346_)
);

NAND2X1 _14200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf2 ),
    .B(\datapath.csr.csr_mepc [4]),
    .Y(_3347_)
);

OAI21X1 _14201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3346_),
    .B(\datapath.regcsrtrap_bF$buf1 ),
    .C(_3347_),
    .Y(\datapath.csr._26_ [2])
);

MUX2X1 _14202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [3]),
    .B(_0_[5]),
    .S(_3339__bF$buf2),
    .Y(_3348_)
);

NAND2X1 _14203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf0 ),
    .B(\datapath.csr.csr_mepc [5]),
    .Y(_3349_)
);

OAI21X1 _14204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3348_),
    .B(\datapath.regcsrtrap_bF$buf7 ),
    .C(_3349_),
    .Y(\datapath.csr._26_ [3])
);

INVX1 _14205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [4]),
    .Y(_3350_)
);

NAND2X1 _14206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3350_),
    .B(_3339__bF$buf1),
    .Y(_3351_)
);

OAI21X1 _14207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[6]),
    .B(_3339__bF$buf0),
    .C(_3351_),
    .Y(_3352_)
);

NAND2X1 _14208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf6 ),
    .B(\datapath.csr.csr_mepc [6]),
    .Y(_3353_)
);

OAI21X1 _14209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3352_),
    .B(\datapath.regcsrtrap_bF$buf5 ),
    .C(_3353_),
    .Y(\datapath.csr._26_ [4])
);

MUX2X1 _14210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [5]),
    .B(_0_[7]),
    .S(_3339__bF$buf6),
    .Y(_3354_)
);

NAND2X1 _14211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf4 ),
    .B(\datapath.csr.csr_mepc [7]),
    .Y(_3355_)
);

OAI21X1 _14212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3354_),
    .B(\datapath.regcsrtrap_bF$buf3 ),
    .C(_3355_),
    .Y(\datapath.csr._26_ [5])
);

INVX1 _14213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [6]),
    .Y(_3356_)
);

NAND2X1 _14214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3356_),
    .B(_3339__bF$buf5),
    .Y(_3357_)
);

OAI21X1 _14215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[8]),
    .B(_3339__bF$buf4),
    .C(_3357_),
    .Y(_3358_)
);

NAND2X1 _14216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf2 ),
    .B(\datapath.csr.csr_mepc [8]),
    .Y(_3359_)
);

OAI21X1 _14217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3358_),
    .B(\datapath.regcsrtrap_bF$buf1 ),
    .C(_3359_),
    .Y(\datapath.csr._26_ [6])
);

INVX1 _14218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [7]),
    .Y(_3360_)
);

NAND2X1 _14219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3360_),
    .B(_3339__bF$buf3),
    .Y(_3361_)
);

OAI21X1 _14220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[9]),
    .B(_3339__bF$buf2),
    .C(_3361_),
    .Y(_3362_)
);

NAND2X1 _14221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf0 ),
    .B(\datapath.csr.csr_mepc [9]),
    .Y(_3363_)
);

OAI21X1 _14222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3362_),
    .B(\datapath.regcsrtrap_bF$buf7 ),
    .C(_3363_),
    .Y(\datapath.csr._26_ [7])
);

MUX2X1 _14223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [8]),
    .B(_0_[10]),
    .S(_3339__bF$buf1),
    .Y(_3364_)
);

NAND2X1 _14224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf6 ),
    .B(\datapath.csr.csr_mepc [10]),
    .Y(_3365_)
);

OAI21X1 _14225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3364_),
    .B(\datapath.regcsrtrap_bF$buf5 ),
    .C(_3365_),
    .Y(\datapath.csr._26_ [8])
);

MUX2X1 _14226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [9]),
    .B(_0_[11]),
    .S(_3339__bF$buf0),
    .Y(_3366_)
);

NAND2X1 _14227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf4 ),
    .B(\datapath.csr.csr_mepc [11]),
    .Y(_3367_)
);

OAI21X1 _14228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3366_),
    .B(\datapath.regcsrtrap_bF$buf3 ),
    .C(_3367_),
    .Y(\datapath.csr._26_ [9])
);

MUX2X1 _14229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [10]),
    .B(_0_[12]),
    .S(_3339__bF$buf6),
    .Y(_3368_)
);

NAND2X1 _14230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf2 ),
    .B(\datapath.csr.csr_mepc [12]),
    .Y(_3369_)
);

OAI21X1 _14231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3368_),
    .B(\datapath.regcsrtrap_bF$buf1 ),
    .C(_3369_),
    .Y(\datapath.csr._26_ [10])
);

INVX1 _14232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [11]),
    .Y(_3370_)
);

NAND2X1 _14233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3370_),
    .B(_3339__bF$buf5),
    .Y(_3371_)
);

OAI21X1 _14234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[13]),
    .B(_3339__bF$buf4),
    .C(_3371_),
    .Y(_3372_)
);

NAND2X1 _14235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf0 ),
    .B(\datapath.csr.csr_mepc [13]),
    .Y(_3373_)
);

OAI21X1 _14236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3372_),
    .B(\datapath.regcsrtrap_bF$buf7 ),
    .C(_3373_),
    .Y(\datapath.csr._26_ [11])
);

INVX1 _14237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [12]),
    .Y(_3374_)
);

NAND2X1 _14238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3374_),
    .B(_3339__bF$buf3),
    .Y(_3375_)
);

OAI21X1 _14239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[14]),
    .B(_3339__bF$buf2),
    .C(_3375_),
    .Y(_3376_)
);

NAND2X1 _14240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf6 ),
    .B(\datapath.csr.csr_mepc [14]),
    .Y(_3377_)
);

OAI21X1 _14241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3376_),
    .B(\datapath.regcsrtrap_bF$buf5 ),
    .C(_3377_),
    .Y(\datapath.csr._26_ [12])
);

MUX2X1 _14242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [13]),
    .B(_0_[15]),
    .S(_3339__bF$buf1),
    .Y(_3378_)
);

NAND2X1 _14243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf4 ),
    .B(\datapath.csr.csr_mepc [15]),
    .Y(_3379_)
);

OAI21X1 _14244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3378_),
    .B(\datapath.regcsrtrap_bF$buf3 ),
    .C(_3379_),
    .Y(\datapath.csr._26_ [13])
);

INVX1 _14245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [14]),
    .Y(_3380_)
);

NAND2X1 _14246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3380_),
    .B(_3339__bF$buf0),
    .Y(_3381_)
);

OAI21X1 _14247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[16]),
    .B(_3339__bF$buf6),
    .C(_3381_),
    .Y(_3382_)
);

NAND2X1 _14248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf2 ),
    .B(\datapath.csr.csr_mepc [16]),
    .Y(_3383_)
);

OAI21X1 _14249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3382_),
    .B(\datapath.regcsrtrap_bF$buf1 ),
    .C(_3383_),
    .Y(\datapath.csr._26_ [14])
);

INVX1 _14250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [15]),
    .Y(_3384_)
);

NAND2X1 _14251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3384_),
    .B(_3339__bF$buf5),
    .Y(_3385_)
);

OAI21X1 _14252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[17]),
    .B(_3339__bF$buf4),
    .C(_3385_),
    .Y(_3386_)
);

NAND2X1 _14253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf0 ),
    .B(\datapath.csr.csr_mepc [17]),
    .Y(_3387_)
);

OAI21X1 _14254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3386_),
    .B(\datapath.regcsrtrap_bF$buf7 ),
    .C(_3387_),
    .Y(\datapath.csr._26_ [15])
);

INVX1 _14255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [16]),
    .Y(_3388_)
);

NAND2X1 _14256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3388_),
    .B(_3339__bF$buf3),
    .Y(_3389_)
);

OAI21X1 _14257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[18]),
    .B(_3339__bF$buf2),
    .C(_3389_),
    .Y(_3390_)
);

NAND2X1 _14258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf6 ),
    .B(\datapath.csr.csr_mepc [18]),
    .Y(_3391_)
);

OAI21X1 _14259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3390_),
    .B(\datapath.regcsrtrap_bF$buf5 ),
    .C(_3391_),
    .Y(\datapath.csr._26_ [16])
);

INVX1 _14260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [17]),
    .Y(_3392_)
);

NAND2X1 _14261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3392_),
    .B(_3339__bF$buf1),
    .Y(_3393_)
);

OAI21X1 _14262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[19]),
    .B(_3339__bF$buf0),
    .C(_3393_),
    .Y(_3394_)
);

NAND2X1 _14263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf4 ),
    .B(\datapath.csr.csr_mepc [19]),
    .Y(_3395_)
);

OAI21X1 _14264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3394_),
    .B(\datapath.regcsrtrap_bF$buf3 ),
    .C(_3395_),
    .Y(\datapath.csr._26_ [17])
);

INVX1 _14265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [18]),
    .Y(_3396_)
);

NAND2X1 _14266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3396_),
    .B(_3339__bF$buf6),
    .Y(_3397_)
);

OAI21X1 _14267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[20]),
    .B(_3339__bF$buf5),
    .C(_3397_),
    .Y(_3398_)
);

NAND2X1 _14268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf2 ),
    .B(\datapath.csr.csr_mepc [20]),
    .Y(_3399_)
);

OAI21X1 _14269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3398_),
    .B(\datapath.regcsrtrap_bF$buf1 ),
    .C(_3399_),
    .Y(\datapath.csr._26_ [18])
);

INVX1 _14270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [19]),
    .Y(_3400_)
);

NAND2X1 _14271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3400_),
    .B(_3339__bF$buf4),
    .Y(_3401_)
);

OAI21X1 _14272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[21]),
    .B(_3339__bF$buf3),
    .C(_3401_),
    .Y(_3402_)
);

NAND2X1 _14273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf0 ),
    .B(\datapath.csr.csr_mepc [21]),
    .Y(_3403_)
);

OAI21X1 _14274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3402_),
    .B(\datapath.regcsrtrap_bF$buf7 ),
    .C(_3403_),
    .Y(\datapath.csr._26_ [19])
);

INVX1 _14275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [20]),
    .Y(_3404_)
);

NAND2X1 _14276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3404_),
    .B(_3339__bF$buf2),
    .Y(_3405_)
);

OAI21X1 _14277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[22]),
    .B(_3339__bF$buf1),
    .C(_3405_),
    .Y(_3406_)
);

NAND2X1 _14278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf6 ),
    .B(\datapath.csr.csr_mepc [22]),
    .Y(_3407_)
);

OAI21X1 _14279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3406_),
    .B(\datapath.regcsrtrap_bF$buf5 ),
    .C(_3407_),
    .Y(\datapath.csr._26_ [20])
);

INVX1 _14280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [21]),
    .Y(_3408_)
);

NAND2X1 _14281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3408_),
    .B(_3339__bF$buf0),
    .Y(_3409_)
);

OAI21X1 _14282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[23]),
    .B(_3339__bF$buf6),
    .C(_3409_),
    .Y(_3410_)
);

NAND2X1 _14283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf4 ),
    .B(\datapath.csr.csr_mepc [23]),
    .Y(_3411_)
);

OAI21X1 _14284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3410_),
    .B(\datapath.regcsrtrap_bF$buf3 ),
    .C(_3411_),
    .Y(\datapath.csr._26_ [21])
);

INVX1 _14285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [22]),
    .Y(_3412_)
);

NAND2X1 _14286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3412_),
    .B(_3339__bF$buf5),
    .Y(_3413_)
);

OAI21X1 _14287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[24]),
    .B(_3339__bF$buf4),
    .C(_3413_),
    .Y(_3414_)
);

NAND2X1 _14288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf2 ),
    .B(\datapath.csr.csr_mepc [24]),
    .Y(_3415_)
);

OAI21X1 _14289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3414_),
    .B(\datapath.regcsrtrap_bF$buf1 ),
    .C(_3415_),
    .Y(\datapath.csr._26_ [22])
);

INVX1 _14290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [23]),
    .Y(_3416_)
);

NAND2X1 _14291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3416_),
    .B(_3339__bF$buf3),
    .Y(_3417_)
);

OAI21X1 _14292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[25]),
    .B(_3339__bF$buf2),
    .C(_3417_),
    .Y(_3418_)
);

NAND2X1 _14293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf0 ),
    .B(\datapath.csr.csr_mepc [25]),
    .Y(_3419_)
);

OAI21X1 _14294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3418_),
    .B(\datapath.regcsrtrap_bF$buf7 ),
    .C(_3419_),
    .Y(\datapath.csr._26_ [23])
);

INVX1 _14295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [24]),
    .Y(_3420_)
);

NAND2X1 _14296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3420_),
    .B(_3339__bF$buf1),
    .Y(_3421_)
);

OAI21X1 _14297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[26]),
    .B(_3339__bF$buf0),
    .C(_3421_),
    .Y(_3422_)
);

NAND2X1 _14298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf6 ),
    .B(\datapath.csr.csr_mepc [26]),
    .Y(_3423_)
);

OAI21X1 _14299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3422_),
    .B(\datapath.regcsrtrap_bF$buf5 ),
    .C(_3423_),
    .Y(\datapath.csr._26_ [24])
);

INVX1 _14300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [25]),
    .Y(_3424_)
);

NAND2X1 _14301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3424_),
    .B(_3339__bF$buf6),
    .Y(_3425_)
);

OAI21X1 _14302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[27]),
    .B(_3339__bF$buf5),
    .C(_3425_),
    .Y(_3426_)
);

NAND2X1 _14303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf4 ),
    .B(\datapath.csr.csr_mepc [27]),
    .Y(_3427_)
);

OAI21X1 _14304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3426_),
    .B(\datapath.regcsrtrap_bF$buf3 ),
    .C(_3427_),
    .Y(\datapath.csr._26_ [25])
);

INVX1 _14305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [26]),
    .Y(_3428_)
);

NAND2X1 _14306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3428_),
    .B(_3339__bF$buf4),
    .Y(_3429_)
);

OAI21X1 _14307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[28]),
    .B(_3339__bF$buf3),
    .C(_3429_),
    .Y(_3430_)
);

NAND2X1 _14308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf2 ),
    .B(\datapath.csr.csr_mepc [28]),
    .Y(_3431_)
);

OAI21X1 _14309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3430_),
    .B(\datapath.regcsrtrap_bF$buf1 ),
    .C(_3431_),
    .Y(\datapath.csr._26_ [26])
);

INVX1 _14310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [27]),
    .Y(_3432_)
);

NAND2X1 _14311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3432_),
    .B(_3339__bF$buf2),
    .Y(_3433_)
);

OAI21X1 _14312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[29]),
    .B(_3339__bF$buf1),
    .C(_3433_),
    .Y(_3434_)
);

NAND2X1 _14313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf0 ),
    .B(\datapath.csr.csr_mepc [29]),
    .Y(_3435_)
);

OAI21X1 _14314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3434_),
    .B(\datapath.regcsrtrap_bF$buf7 ),
    .C(_3435_),
    .Y(\datapath.csr._26_ [27])
);

INVX1 _14315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [28]),
    .Y(_3436_)
);

NAND2X1 _14316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3436_),
    .B(_3339__bF$buf0),
    .Y(_3437_)
);

OAI21X1 _14317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[30]),
    .B(_3339__bF$buf6),
    .C(_3437_),
    .Y(_3438_)
);

NAND2X1 _14318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf6 ),
    .B(\datapath.csr.csr_mepc [30]),
    .Y(_3439_)
);

OAI21X1 _14319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3438_),
    .B(\datapath.regcsrtrap_bF$buf5 ),
    .C(_3439_),
    .Y(\datapath.csr._26_ [28])
);

MUX2X1 _14320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [29]),
    .B(_0_[31]),
    .S(_3339__bF$buf5),
    .Y(_3440_)
);

NAND2X1 _14321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf4 ),
    .B(\datapath.csr.csr_mepc [31]),
    .Y(_3441_)
);

OAI21X1 _14322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3440_),
    .B(\datapath.regcsrtrap_bF$buf3 ),
    .C(_3441_),
    .Y(\datapath.csr._26_ [29])
);

NAND2X1 _14323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf2 ),
    .B(\datapath.csr.csr_mcause [0]),
    .Y(_3442_)
);

NAND2X1 _14324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [21]),
    .B(_3331_),
    .Y(_3443_)
);

NOR2X1 _14325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3251_),
    .B(_3443_),
    .Y(_3444_)
);

NAND2X1 _14326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3444_),
    .B(_3338_),
    .Y(_3445_)
);

INVX2 _14327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3445_),
    .Y(_3446_)
);

NOR2X1 _14328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [0]),
    .B(_3446_),
    .Y(_3447_)
);

INVX8 _14329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf1 ),
    .Y(_3448_)
);

OAI21X1 _14330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3445_),
    .B(_0__0_bF$buf4),
    .C(_3448__bF$buf4),
    .Y(_3449_)
);

OAI21X1 _14331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3447_),
    .B(_3449_),
    .C(_3442_),
    .Y(\datapath.csr._32_ [0])
);

NAND2X1 _14332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf0 ),
    .B(\datapath.csr.csr_mcause [1]),
    .Y(_3450_)
);

NOR2X1 _14333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [1]),
    .B(_3446_),
    .Y(_3451_)
);

OAI21X1 _14334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3445_),
    .B(_0__1_bF$buf4),
    .C(_3448__bF$buf3),
    .Y(_3452_)
);

OAI21X1 _14335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3451_),
    .B(_3452_),
    .C(_3450_),
    .Y(\datapath.csr._32_ [1])
);

NAND2X1 _14336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf7 ),
    .B(\datapath.csr.csr_mcause [2]),
    .Y(_3453_)
);

NOR2X1 _14337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [2]),
    .B(_3446_),
    .Y(_3454_)
);

OAI21X1 _14338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3445_),
    .B(_0_[2]),
    .C(_3448__bF$buf2),
    .Y(_3455_)
);

OAI21X1 _14339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3454_),
    .B(_3455_),
    .C(_3453_),
    .Y(\datapath.csr._32_ [2])
);

NAND2X1 _14340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf6 ),
    .B(\datapath.csr.csr_mcause [3]),
    .Y(_3456_)
);

NOR2X1 _14341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [3]),
    .B(_3446_),
    .Y(_3457_)
);

OAI21X1 _14342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3445_),
    .B(_0_[3]),
    .C(_3448__bF$buf1),
    .Y(_3458_)
);

OAI21X1 _14343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3457_),
    .B(_3458_),
    .C(_3456_),
    .Y(\datapath.csr._32_ [3])
);

INVX1 _14344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [4]),
    .Y(_3459_)
);

NAND3X1 _14345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [29]),
    .B(_3253_),
    .C(_3257_),
    .Y(_3460_)
);

NAND3X1 _14346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [26]),
    .B(_3254_),
    .C(_3260_),
    .Y(_3461_)
);

NOR2X1 _14347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3461_),
    .B(_3460_),
    .Y(_3462_)
);

NAND3X1 _14348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3336_),
    .B(_3444_),
    .C(_3462_),
    .Y(_3463_)
);

OAI21X1 _14349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf6),
    .B(_0_[4]),
    .C(_3448__bF$buf0),
    .Y(_3464_)
);

AOI21X1 _14350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3459_),
    .B(_3463__bF$buf5),
    .C(_3464_),
    .Y(\datapath.csr._32_ [4])
);

INVX1 _14351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [5]),
    .Y(_3465_)
);

OAI21X1 _14352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf4),
    .B(_0_[5]),
    .C(_3448__bF$buf4),
    .Y(_3466_)
);

AOI21X1 _14353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3465_),
    .B(_3463__bF$buf3),
    .C(_3466_),
    .Y(\datapath.csr._32_ [5])
);

INVX1 _14354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [6]),
    .Y(_3467_)
);

OAI21X1 _14355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf2),
    .B(_0_[6]),
    .C(_3448__bF$buf3),
    .Y(_3468_)
);

AOI21X1 _14356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3467_),
    .B(_3463__bF$buf1),
    .C(_3468_),
    .Y(\datapath.csr._32_ [6])
);

INVX1 _14357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [7]),
    .Y(_3469_)
);

OAI21X1 _14358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf0),
    .B(_0_[7]),
    .C(_3448__bF$buf2),
    .Y(_3470_)
);

AOI21X1 _14359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3469_),
    .B(_3463__bF$buf6),
    .C(_3470_),
    .Y(\datapath.csr._32_ [7])
);

INVX1 _14360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [8]),
    .Y(_3471_)
);

OAI21X1 _14361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf5),
    .B(_0_[8]),
    .C(_3448__bF$buf1),
    .Y(_3472_)
);

AOI21X1 _14362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3471_),
    .B(_3463__bF$buf4),
    .C(_3472_),
    .Y(\datapath.csr._32_ [8])
);

INVX1 _14363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [9]),
    .Y(_3473_)
);

OAI21X1 _14364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf3),
    .B(_0_[9]),
    .C(_3448__bF$buf0),
    .Y(_3474_)
);

AOI21X1 _14365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3473_),
    .B(_3463__bF$buf2),
    .C(_3474_),
    .Y(\datapath.csr._32_ [9])
);

INVX1 _14366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [10]),
    .Y(_3475_)
);

OAI21X1 _14367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf1),
    .B(_0_[10]),
    .C(_3448__bF$buf4),
    .Y(_3476_)
);

AOI21X1 _14368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3475_),
    .B(_3463__bF$buf0),
    .C(_3476_),
    .Y(\datapath.csr._32_ [10])
);

INVX1 _14369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [11]),
    .Y(_3477_)
);

OAI21X1 _14370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf6),
    .B(_0_[11]),
    .C(_3448__bF$buf3),
    .Y(_3478_)
);

AOI21X1 _14371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3477_),
    .B(_3463__bF$buf5),
    .C(_3478_),
    .Y(\datapath.csr._32_ [11])
);

INVX1 _14372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [12]),
    .Y(_3479_)
);

OAI21X1 _14373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf4),
    .B(_0_[12]),
    .C(_3448__bF$buf2),
    .Y(_3480_)
);

AOI21X1 _14374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3479_),
    .B(_3463__bF$buf3),
    .C(_3480_),
    .Y(\datapath.csr._32_ [12])
);

INVX1 _14375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [13]),
    .Y(_3481_)
);

OAI21X1 _14376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf2),
    .B(_0_[13]),
    .C(_3448__bF$buf1),
    .Y(_3482_)
);

AOI21X1 _14377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3481_),
    .B(_3463__bF$buf1),
    .C(_3482_),
    .Y(\datapath.csr._32_ [13])
);

INVX1 _14378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [14]),
    .Y(_3483_)
);

OAI21X1 _14379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf0),
    .B(_0_[14]),
    .C(_3448__bF$buf0),
    .Y(_3484_)
);

AOI21X1 _14380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3483_),
    .B(_3463__bF$buf6),
    .C(_3484_),
    .Y(\datapath.csr._32_ [14])
);

INVX1 _14381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [15]),
    .Y(_3485_)
);

OAI21X1 _14382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf5),
    .B(_0_[15]),
    .C(_3448__bF$buf4),
    .Y(_3486_)
);

AOI21X1 _14383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3485_),
    .B(_3463__bF$buf4),
    .C(_3486_),
    .Y(\datapath.csr._32_ [15])
);

INVX1 _14384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [16]),
    .Y(_3487_)
);

OAI21X1 _14385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf3),
    .B(_0_[16]),
    .C(_3448__bF$buf3),
    .Y(_3488_)
);

AOI21X1 _14386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3487_),
    .B(_3463__bF$buf2),
    .C(_3488_),
    .Y(\datapath.csr._32_ [16])
);

INVX1 _14387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [17]),
    .Y(_3489_)
);

OAI21X1 _14388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf1),
    .B(_0_[17]),
    .C(_3448__bF$buf2),
    .Y(_3490_)
);

AOI21X1 _14389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3489_),
    .B(_3463__bF$buf0),
    .C(_3490_),
    .Y(\datapath.csr._32_ [17])
);

INVX1 _14390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [18]),
    .Y(_3491_)
);

OAI21X1 _14391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf6),
    .B(_0_[18]),
    .C(_3448__bF$buf1),
    .Y(_3492_)
);

AOI21X1 _14392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3491_),
    .B(_3463__bF$buf5),
    .C(_3492_),
    .Y(\datapath.csr._32_ [18])
);

INVX1 _14393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [19]),
    .Y(_3493_)
);

OAI21X1 _14394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf4),
    .B(_0_[19]),
    .C(_3448__bF$buf0),
    .Y(_3494_)
);

AOI21X1 _14395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3493_),
    .B(_3463__bF$buf3),
    .C(_3494_),
    .Y(\datapath.csr._32_ [19])
);

INVX1 _14396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [20]),
    .Y(_3495_)
);

OAI21X1 _14397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf2),
    .B(_0_[20]),
    .C(_3448__bF$buf4),
    .Y(_3496_)
);

AOI21X1 _14398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3495_),
    .B(_3463__bF$buf1),
    .C(_3496_),
    .Y(\datapath.csr._32_ [20])
);

INVX1 _14399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [21]),
    .Y(_3497_)
);

OAI21X1 _14400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf0),
    .B(_0_[21]),
    .C(_3448__bF$buf3),
    .Y(_3498_)
);

AOI21X1 _14401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3497_),
    .B(_3463__bF$buf6),
    .C(_3498_),
    .Y(\datapath.csr._32_ [21])
);

INVX1 _14402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [22]),
    .Y(_3499_)
);

OAI21X1 _14403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf5),
    .B(_0_[22]),
    .C(_3448__bF$buf2),
    .Y(_3500_)
);

AOI21X1 _14404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3499_),
    .B(_3463__bF$buf4),
    .C(_3500_),
    .Y(\datapath.csr._32_ [22])
);

INVX1 _14405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [23]),
    .Y(_3501_)
);

OAI21X1 _14406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf3),
    .B(_0_[23]),
    .C(_3448__bF$buf1),
    .Y(_3502_)
);

AOI21X1 _14407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3501_),
    .B(_3463__bF$buf2),
    .C(_3502_),
    .Y(\datapath.csr._32_ [23])
);

INVX1 _14408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [24]),
    .Y(_3503_)
);

OAI21X1 _14409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf1),
    .B(_0_[24]),
    .C(_3448__bF$buf0),
    .Y(_3504_)
);

AOI21X1 _14410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3503_),
    .B(_3463__bF$buf0),
    .C(_3504_),
    .Y(\datapath.csr._32_ [24])
);

INVX1 _14411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [25]),
    .Y(_3505_)
);

OAI21X1 _14412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf6),
    .B(_0_[25]),
    .C(_3448__bF$buf4),
    .Y(_3506_)
);

AOI21X1 _14413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3505_),
    .B(_3463__bF$buf5),
    .C(_3506_),
    .Y(\datapath.csr._32_ [25])
);

INVX1 _14414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [26]),
    .Y(_3507_)
);

OAI21X1 _14415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf4),
    .B(_0_[26]),
    .C(_3448__bF$buf3),
    .Y(_3508_)
);

AOI21X1 _14416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3507_),
    .B(_3463__bF$buf3),
    .C(_3508_),
    .Y(\datapath.csr._32_ [26])
);

INVX1 _14417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [27]),
    .Y(_3509_)
);

OAI21X1 _14418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf2),
    .B(_0_[27]),
    .C(_3448__bF$buf2),
    .Y(_3510_)
);

AOI21X1 _14419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3509_),
    .B(_3463__bF$buf1),
    .C(_3510_),
    .Y(\datapath.csr._32_ [27])
);

INVX1 _14420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [28]),
    .Y(_3511_)
);

OAI21X1 _14421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf0),
    .B(_0_[28]),
    .C(_3448__bF$buf1),
    .Y(_3512_)
);

AOI21X1 _14422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3511_),
    .B(_3463__bF$buf6),
    .C(_3512_),
    .Y(\datapath.csr._32_ [28])
);

INVX1 _14423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [29]),
    .Y(_3513_)
);

OAI21X1 _14424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf5),
    .B(_0_[29]),
    .C(_3448__bF$buf0),
    .Y(_3514_)
);

AOI21X1 _14425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3513_),
    .B(_3463__bF$buf4),
    .C(_3514_),
    .Y(\datapath.csr._32_ [29])
);

INVX1 _14426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [30]),
    .Y(_3515_)
);

OAI21X1 _14427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463__bF$buf3),
    .B(_0_[30]),
    .C(_3448__bF$buf4),
    .Y(_3516_)
);

AOI21X1 _14428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3515_),
    .B(_3463__bF$buf2),
    .C(_3516_),
    .Y(\datapath.csr._32_ [30])
);

NAND3X1 _14429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mie ),
    .B(\datapath.csr.mip ),
    .C(\datapath.csr.mstatus [0]),
    .Y(_3517_)
);

INVX1 _14430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3517_),
    .Y(\datapath.csr.csr_irq )
);

NAND3X1 _14431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3448__bF$buf3),
    .B(\datapath.csr.mcause [31]),
    .C(_3445_),
    .Y(_3518_)
);

OAI21X1 _14432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3448__bF$buf2),
    .B(_3517_),
    .C(_3518_),
    .Y(\datapath.csr._32_ [31])
);

INVX1 _14433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3336_),
    .Y(_3519_)
);

NOR2X1 _14434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3332_),
    .B(_3519_),
    .Y(_3520_)
);

NAND3X1 _14435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.allowcsrwrite ),
    .B(_3520_),
    .C(_3262_),
    .Y(_3521_)
);

INVX2 _14436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mstatus [0]),
    .Y(_3522_)
);

NAND2X1 _14437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3522_),
    .B(_3521_),
    .Y(_3523_)
);

OAI21X1 _14438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[3]),
    .B(_3521_),
    .C(_3523_),
    .Y(_3524_)
);

OAI21X1 _14439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf4),
    .B(\datapath.csr.mstatus [1]),
    .C(_3448__bF$buf1),
    .Y(_3525_)
);

AOI21X1 _14440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf3),
    .B(_3524_),
    .C(_3525_),
    .Y(\datapath.csr._37_ [0])
);

MUX2X1 _14441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mstatus [1]),
    .B(_0_[7]),
    .S(_3521_),
    .Y(_3526_)
);

NOR2X1 _14442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret_bF$buf2 ),
    .B(\datapath.regcsrtrap_bF$buf5 ),
    .Y(_3527_)
);

AOI22X1 _14443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regcsrtrap_bF$buf4 ),
    .B(_3522_),
    .C(_3526_),
    .D(_3527_),
    .Y(\datapath.csr._37_ [1])
);

NOR2X1 _14444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3247_),
    .B(_3517_),
    .Y(_3528_)
);

NAND2X1 _14445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3271_),
    .B(_3528_),
    .Y(_3529_)
);

INVX2 _14446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3528_),
    .Y(_3530_)
);

AOI21X1 _14447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [2]),
    .B(_3530_),
    .C(\datapath.regmret_bF$buf1 ),
    .Y(_3531_)
);

AOI22X1 _14448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret_bF$buf0 ),
    .B(_3340_),
    .C(_3531_),
    .D(_3529_),
    .Y(\datapath.csr.csr_pcaddr [2])
);

XNOR2X1 _14449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529_),
    .B(_3273_),
    .Y(_3532_)
);

NAND2X1 _14450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret_bF$buf4 ),
    .B(\datapath.csr.mepc [1]),
    .Y(_3533_)
);

OAI21X1 _14451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3532_),
    .B(\datapath.regmret_bF$buf3 ),
    .C(_3533_),
    .Y(\datapath.csr.csr_pcaddr [3])
);

NOR2X1 _14452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [2]),
    .B(\datapath.csr.mvect [3]),
    .Y(_3534_)
);

OAI21X1 _14453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3530_),
    .B(_3534_),
    .C(_3275_),
    .Y(_3535_)
);

OAI21X1 _14454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [2]),
    .B(\datapath.csr.mvect [3]),
    .C(\datapath.csr.mvect [4]),
    .Y(_3536_)
);

OAI21X1 _14455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3530_),
    .B(_3536_),
    .C(_3535_),
    .Y(_3537_)
);

NAND2X1 _14456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret_bF$buf2 ),
    .B(\datapath.csr.mepc [2]),
    .Y(_3538_)
);

OAI21X1 _14457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3537_),
    .B(\datapath.regmret_bF$buf1 ),
    .C(_3538_),
    .Y(\datapath.csr.csr_pcaddr [4])
);

OAI21X1 _14458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3275_),
    .B(_3534_),
    .C(_3528_),
    .Y(_3539_)
);

XNOR2X1 _14459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3539_),
    .B(_3277_),
    .Y(_3540_)
);

NAND2X1 _14460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret_bF$buf0 ),
    .B(\datapath.csr.mepc [3]),
    .Y(_3541_)
);

OAI21X1 _14461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3540_),
    .B(\datapath.regmret_bF$buf4 ),
    .C(_3541_),
    .Y(\datapath.csr.csr_pcaddr [5])
);

OAI21X1 _14462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3534_),
    .B(_3275_),
    .C(_3277_),
    .Y(_3542_)
);

AOI21X1 _14463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3528_),
    .B(_3542_),
    .C(\datapath.csr.mvect [6]),
    .Y(_3543_)
);

NAND2X1 _14464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3528_),
    .B(_3542_),
    .Y(_3544_)
);

OAI21X1 _14465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3544_),
    .B(_3279_),
    .C(_3250__bF$buf2),
    .Y(_3545_)
);

OAI22X1 _14466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf1),
    .B(_3350_),
    .C(_3545_),
    .D(_3543_),
    .Y(\datapath.csr.csr_pcaddr [6])
);

OAI21X1 _14467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3544_),
    .B(_3279_),
    .C(_3281_),
    .Y(_3546_)
);

NAND2X1 _14468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [6]),
    .B(\datapath.csr.mvect [7]),
    .Y(_3547_)
);

OAI21X1 _14469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3544_),
    .B(_3547_),
    .C(_3546_),
    .Y(_3548_)
);

NAND2X1 _14470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret_bF$buf3 ),
    .B(\datapath.csr.mepc [5]),
    .Y(_3549_)
);

OAI21X1 _14471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3548_),
    .B(\datapath.regmret_bF$buf2 ),
    .C(_3549_),
    .Y(\datapath.csr.csr_pcaddr [7])
);

AOI21X1 _14472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3277_),
    .B(_3536_),
    .C(_3547_),
    .Y(_3550_)
);

AND2X2 _14473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3550_),
    .B(_3528_),
    .Y(_3551_)
);

NAND2X1 _14474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [8]),
    .B(_3551_),
    .Y(_3552_)
);

INVX1 _14475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3552_),
    .Y(_3553_)
);

OAI21X1 _14476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3551_),
    .B(\datapath.csr.mvect [8]),
    .C(_3250__bF$buf0),
    .Y(_3554_)
);

OAI22X1 _14477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf5),
    .B(_3356_),
    .C(_3553_),
    .D(_3554_),
    .Y(\datapath.csr.csr_pcaddr [8])
);

NAND2X1 _14478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3528_),
    .B(_3550_),
    .Y(_3555_)
);

OAI21X1 _14479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3555_),
    .B(_3283_),
    .C(_3285_),
    .Y(_3556_)
);

NAND2X1 _14480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [8]),
    .B(\datapath.csr.mvect [9]),
    .Y(_3557_)
);

OR2X2 _14481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3555_),
    .B(_3557_),
    .Y(_3558_)
);

NAND3X1 _14482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf4),
    .B(_3556_),
    .C(_3558_),
    .Y(_3559_)
);

OAI21X1 _14483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf3),
    .B(_3360_),
    .C(_3559_),
    .Y(\datapath.csr.csr_pcaddr [9])
);

XNOR2X1 _14484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3558_),
    .B(_3287_),
    .Y(_3560_)
);

NAND2X1 _14485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret_bF$buf1 ),
    .B(\datapath.csr.mepc [8]),
    .Y(_3561_)
);

OAI21X1 _14486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3560_),
    .B(\datapath.regmret_bF$buf0 ),
    .C(_3561_),
    .Y(\datapath.csr.csr_pcaddr [10])
);

OAI21X1 _14487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3558_),
    .B(_3287_),
    .C(_3290_),
    .Y(_3562_)
);

NAND2X1 _14488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [10]),
    .B(\datapath.csr.mvect [11]),
    .Y(_3563_)
);

OR2X2 _14489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3557_),
    .B(_3563_),
    .Y(_3564_)
);

OAI21X1 _14490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3555_),
    .B(_3564_),
    .C(_3562_),
    .Y(_3565_)
);

NAND2X1 _14491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret_bF$buf4 ),
    .B(\datapath.csr.mepc [9]),
    .Y(_3566_)
);

OAI21X1 _14492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3565_),
    .B(\datapath.regmret_bF$buf3 ),
    .C(_3566_),
    .Y(\datapath.csr.csr_pcaddr [11])
);

NOR2X1 _14493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3557_),
    .B(_3563_),
    .Y(_3567_)
);

NAND3X1 _14494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3528_),
    .B(_3567_),
    .C(_3550_),
    .Y(_3568_)
);

XNOR2X1 _14495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3568_),
    .B(_3291_),
    .Y(_3569_)
);

NAND2X1 _14496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret_bF$buf2 ),
    .B(\datapath.csr.mepc [10]),
    .Y(_3570_)
);

OAI21X1 _14497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3569_),
    .B(\datapath.regmret_bF$buf1 ),
    .C(_3570_),
    .Y(\datapath.csr.csr_pcaddr [12])
);

OAI21X1 _14498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3568_),
    .B(_3291_),
    .C(_3293_),
    .Y(_3571_)
);

INVX1 _14499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3571_),
    .Y(_3572_)
);

NAND2X1 _14500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [12]),
    .B(\datapath.csr.mvect [13]),
    .Y(_3573_)
);

OAI21X1 _14501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3568_),
    .B(_3573_),
    .C(_3250__bF$buf2),
    .Y(_3574_)
);

OAI22X1 _14502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf1),
    .B(_3370_),
    .C(_3572_),
    .D(_3574_),
    .Y(\datapath.csr.csr_pcaddr [13])
);

OAI21X1 _14503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3568_),
    .B(_3573_),
    .C(_3295_),
    .Y(_3575_)
);

INVX1 _14504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3575_),
    .Y(_3576_)
);

OR2X2 _14505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3568_),
    .B(_3573_),
    .Y(_3577_)
);

OAI21X1 _14506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3577_),
    .B(_3295_),
    .C(_3250__bF$buf0),
    .Y(_3578_)
);

OAI22X1 _14507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf5),
    .B(_3374_),
    .C(_3578_),
    .D(_3576_),
    .Y(\datapath.csr.csr_pcaddr [14])
);

NAND2X1 _14508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret_bF$buf0 ),
    .B(\datapath.csr.mepc [13]),
    .Y(_3579_)
);

OAI21X1 _14509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3577_),
    .B(_3295_),
    .C(_3297_),
    .Y(_3580_)
);

INVX1 _14510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3580_),
    .Y(_3581_)
);

NAND2X1 _14511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [14]),
    .B(\datapath.csr.mvect [15]),
    .Y(_3582_)
);

OR2X2 _14512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3573_),
    .B(_3582_),
    .Y(_3583_)
);

OAI21X1 _14513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3568_),
    .B(_3583_),
    .C(_3250__bF$buf4),
    .Y(_3584_)
);

OAI21X1 _14514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3581_),
    .B(_3584_),
    .C(_3579_),
    .Y(\datapath.csr.csr_pcaddr [15])
);

NOR2X1 _14515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3573_),
    .B(_3582_),
    .Y(_3585_)
);

NAND3X1 _14516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3567_),
    .B(_3585_),
    .C(_3550_),
    .Y(_3586_)
);

NOR2X1 _14517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3530_),
    .B(_3586_),
    .Y(_3587_)
);

NOR2X1 _14518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [16]),
    .B(_3587_),
    .Y(_3588_)
);

NOR2X1 _14519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3583_),
    .B(_3568_),
    .Y(_3589_)
);

INVX2 _14520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3589_),
    .Y(_3590_)
);

OAI21X1 _14521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3590_),
    .B(_3299_),
    .C(_3250__bF$buf3),
    .Y(_3591_)
);

OAI22X1 _14522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf2),
    .B(_3380_),
    .C(_3591_),
    .D(_3588_),
    .Y(\datapath.csr.csr_pcaddr [16])
);

AOI21X1 _14523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [16]),
    .B(_3587_),
    .C(\datapath.csr.mvect [17]),
    .Y(_3592_)
);

NAND2X1 _14524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [16]),
    .B(\datapath.csr.mvect [17]),
    .Y(_3593_)
);

OAI21X1 _14525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3590_),
    .B(_3593_),
    .C(_3250__bF$buf1),
    .Y(_3594_)
);

OAI22X1 _14526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf0),
    .B(_3384_),
    .C(_3594_),
    .D(_3592_),
    .Y(\datapath.csr.csr_pcaddr [17])
);

AND2X2 _14527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [16]),
    .B(\datapath.csr.mvect [17]),
    .Y(_3595_)
);

AOI21X1 _14528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3595_),
    .B(_3589_),
    .C(\datapath.csr.mvect [18]),
    .Y(_3596_)
);

NAND2X1 _14529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [18]),
    .B(_3595_),
    .Y(_3597_)
);

OAI21X1 _14530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3590_),
    .B(_3597_),
    .C(_3250__bF$buf5),
    .Y(_3598_)
);

OAI22X1 _14531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf4),
    .B(_3388_),
    .C(_3598_),
    .D(_3596_),
    .Y(\datapath.csr.csr_pcaddr [18])
);

INVX1 _14532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3597_),
    .Y(_3599_)
);

AOI21X1 _14533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3599_),
    .B(_3587_),
    .C(\datapath.csr.mvect [19]),
    .Y(_3600_)
);

AND2X2 _14534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [18]),
    .B(\datapath.csr.mvect [19]),
    .Y(_3601_)
);

NAND2X1 _14535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3595_),
    .B(_3601_),
    .Y(_3602_)
);

OAI21X1 _14536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3590_),
    .B(_3602_),
    .C(_3250__bF$buf3),
    .Y(_3603_)
);

OAI22X1 _14537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf2),
    .B(_3392_),
    .C(_3603_),
    .D(_3600_),
    .Y(\datapath.csr.csr_pcaddr [19])
);

NAND3X1 _14538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3595_),
    .B(_3601_),
    .C(_3589_),
    .Y(_3604_)
);

AND2X2 _14539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3604_),
    .B(_3307_),
    .Y(_3605_)
);

OAI21X1 _14540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3604_),
    .B(_3307_),
    .C(_3250__bF$buf1),
    .Y(_3606_)
);

OAI22X1 _14541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf0),
    .B(_3396_),
    .C(_3605_),
    .D(_3606_),
    .Y(\datapath.csr.csr_pcaddr [20])
);

NOR2X1 _14542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3307_),
    .B(_3602_),
    .Y(_3607_)
);

AOI21X1 _14543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3607_),
    .B(_3587_),
    .C(\datapath.csr.mvect [21]),
    .Y(_3608_)
);

AND2X2 _14544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [20]),
    .B(\datapath.csr.mvect [21]),
    .Y(_3609_)
);

NAND3X1 _14545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3595_),
    .B(_3601_),
    .C(_3609_),
    .Y(_3610_)
);

OAI21X1 _14546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3590_),
    .B(_3610_),
    .C(_3250__bF$buf5),
    .Y(_3611_)
);

OAI22X1 _14547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf4),
    .B(_3400_),
    .C(_3611_),
    .D(_3608_),
    .Y(\datapath.csr.csr_pcaddr [21])
);

NAND2X1 _14548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [18]),
    .B(\datapath.csr.mvect [19]),
    .Y(_3612_)
);

NAND2X1 _14549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [20]),
    .B(\datapath.csr.mvect [21]),
    .Y(_3613_)
);

NOR3X1 _14550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3593_),
    .B(_3612_),
    .C(_3613_),
    .Y(_3614_)
);

NAND3X1 _14551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3567_),
    .B(_3585_),
    .C(_3614_),
    .Y(_3615_)
);

NOR2X1 _14552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3555_),
    .B(_3615_),
    .Y(_3616_)
);

AOI21X1 _14553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [22]),
    .B(_3616_),
    .C(\datapath.regmret_bF$buf4 ),
    .Y(_3617_)
);

OAI21X1 _14554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [22]),
    .B(_3616_),
    .C(_3617_),
    .Y(_3618_)
);

OAI21X1 _14555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf3),
    .B(_3404_),
    .C(_3618_),
    .Y(\datapath.csr.csr_pcaddr [22])
);

NAND2X1 _14556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [22]),
    .B(_3616_),
    .Y(_3619_)
);

OR2X2 _14557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3619_),
    .B(\datapath.csr.mvect [23]),
    .Y(_3620_)
);

AOI21X1 _14558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [23]),
    .B(_3619_),
    .C(\datapath.regmret_bF$buf3 ),
    .Y(_3621_)
);

AOI22X1 _14559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret_bF$buf2 ),
    .B(_3408_),
    .C(_3620_),
    .D(_3621_),
    .Y(\datapath.csr.csr_pcaddr [23])
);

NAND2X1 _14560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [22]),
    .B(\datapath.csr.mvect [23]),
    .Y(_3622_)
);

NOR3X1 _14561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3555_),
    .B(_3622_),
    .C(_3615_),
    .Y(_3623_)
);

NOR2X1 _14562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [24]),
    .B(_3623_),
    .Y(_3624_)
);

INVX1 _14563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3623_),
    .Y(_3625_)
);

OAI21X1 _14564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3625_),
    .B(_3315_),
    .C(_3250__bF$buf2),
    .Y(_3626_)
);

OAI22X1 _14565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf1),
    .B(_3412_),
    .C(_3626_),
    .D(_3624_),
    .Y(\datapath.csr.csr_pcaddr [24])
);

AOI21X1 _14566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [24]),
    .B(_3623_),
    .C(\datapath.csr.mvect [25]),
    .Y(_3627_)
);

NAND2X1 _14567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [24]),
    .B(\datapath.csr.mvect [25]),
    .Y(_3628_)
);

OAI21X1 _14568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3625_),
    .B(_3628_),
    .C(_3250__bF$buf0),
    .Y(_3629_)
);

OAI22X1 _14569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf5),
    .B(_3416_),
    .C(_3629_),
    .D(_3627_),
    .Y(\datapath.csr.csr_pcaddr [25])
);

INVX1 _14570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3628_),
    .Y(_3630_)
);

AOI21X1 _14571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3630_),
    .B(_3623_),
    .C(\datapath.csr.mvect [26]),
    .Y(_3631_)
);

NAND3X1 _14572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [26]),
    .B(_3630_),
    .C(_3623_),
    .Y(_3632_)
);

NAND2X1 _14573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf4),
    .B(_3632_),
    .Y(_3633_)
);

OAI22X1 _14574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf3),
    .B(_3420_),
    .C(_3633_),
    .D(_3631_),
    .Y(\datapath.csr.csr_pcaddr [26])
);

NAND3X1 _14575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf2),
    .B(_3321_),
    .C(_3632_),
    .Y(_3634_)
);

NAND2X1 _14576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [26]),
    .B(\datapath.csr.mvect [27]),
    .Y(_3635_)
);

NOR2X1 _14577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3628_),
    .B(_3635_),
    .Y(_3636_)
);

AND2X2 _14578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3636_),
    .B(_3250__bF$buf1),
    .Y(_3637_)
);

AOI22X1 _14579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret_bF$buf1 ),
    .B(_3424_),
    .C(_3623_),
    .D(_3637_),
    .Y(_3638_)
);

AND2X2 _14580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3634_),
    .B(_3638_),
    .Y(\datapath.csr.csr_pcaddr [27])
);

NOR3X1 _14581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3622_),
    .B(_3628_),
    .C(_3635_),
    .Y(_3639_)
);

INVX1 _14582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3639_),
    .Y(_3640_)
);

NOR3X1 _14583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3555_),
    .B(_3640_),
    .C(_3615_),
    .Y(_3641_)
);

NOR2X1 _14584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [28]),
    .B(_3641_),
    .Y(_3642_)
);

NOR3X1 _14585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3564_),
    .B(_3583_),
    .C(_3610_),
    .Y(_3643_)
);

NAND3X1 _14586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3551_),
    .B(_3639_),
    .C(_3643_),
    .Y(_3644_)
);

OAI21X1 _14587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3644_),
    .B(_3323_),
    .C(_3250__bF$buf0),
    .Y(_3645_)
);

OAI22X1 _14588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf5),
    .B(_3428_),
    .C(_3645_),
    .D(_3642_),
    .Y(\datapath.csr.csr_pcaddr [28])
);

NAND2X1 _14589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [28]),
    .B(_3641_),
    .Y(_3646_)
);

OR2X2 _14590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646_),
    .B(\datapath.csr.mvect [29]),
    .Y(_3647_)
);

AOI21X1 _14591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [29]),
    .B(_3646_),
    .C(\datapath.regmret_bF$buf0 ),
    .Y(_3648_)
);

AOI22X1 _14592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret_bF$buf4 ),
    .B(_3432_),
    .C(_3647_),
    .D(_3648_),
    .Y(\datapath.csr.csr_pcaddr [29])
);

NAND2X1 _14593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [28]),
    .B(\datapath.csr.mvect [29]),
    .Y(_3649_)
);

NOR3X1 _14594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3247_),
    .B(_3649_),
    .C(_3517_),
    .Y(_3650_)
);

NAND3X1 _14595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3550_),
    .B(_3639_),
    .C(_3650_),
    .Y(_3651_)
);

OAI21X1 _14596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3651_),
    .B(_3615_),
    .C(\datapath.csr.mvect [30]),
    .Y(_3652_)
);

INVX1 _14597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3652_),
    .Y(_3653_)
);

NOR2X1 _14598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3615_),
    .B(_3651_),
    .Y(_3654_)
);

AND2X2 _14599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3654_),
    .B(_3327_),
    .Y(_3655_)
);

OAI21X1 _14600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3655_),
    .B(_3653_),
    .C(_3250__bF$buf4),
    .Y(_3656_)
);

OAI21X1 _14601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3250__bF$buf3),
    .B(_3436_),
    .C(_3656_),
    .Y(\datapath.csr.csr_pcaddr [30])
);

INVX1 _14602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3649_),
    .Y(_3657_)
);

NAND2X1 _14603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [30]),
    .B(_3657_),
    .Y(_3658_)
);

INVX1 _14604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3658_),
    .Y(_3659_)
);

AOI21X1 _14605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3659_),
    .B(_3641_),
    .C(_3329_),
    .Y(_3660_)
);

NOR3X1 _14606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [31]),
    .B(_3658_),
    .C(_3644_),
    .Y(_3661_)
);

OAI21X1 _14607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3661_),
    .B(_3660_),
    .C(_3250__bF$buf2),
    .Y(_3662_)
);

NAND2X1 _14608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regmret_bF$buf3 ),
    .B(\datapath.csr.mepc [29]),
    .Y(_3663_)
);

NAND2X1 _14609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3663_),
    .B(_3662_),
    .Y(\datapath.csr.csr_pcaddr [31])
);

NOR2X1 _14610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [31]),
    .B(\datapath.idinstr [30]),
    .Y(_3664_)
);

NAND3X1 _14611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [29]),
    .B(\datapath.idinstr [28]),
    .C(_3664_),
    .Y(_3665_)
);

INVX1 _14612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [27]),
    .Y(_3666_)
);

NOR2X1 _14613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [25]),
    .B(\datapath.idinstr_24_bF$buf4 ),
    .Y(_3667_)
);

NAND3X1 _14614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3666_),
    .B(\datapath.idinstr [26]),
    .C(_3667_),
    .Y(_3668_)
);

NOR2X1 _14615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3665_),
    .B(_3668_),
    .Y(_3669_)
);

NOR2X1 _14616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_23_bF$buf6 ),
    .B(\datapath.idinstr_22_bF$buf42 ),
    .Y(_3670_)
);

INVX1 _14617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3670_),
    .Y(_3671_)
);

INVX1 _14618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf54 ),
    .Y(_3672_)
);

NAND2X1 _14619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf43 ),
    .B(_3672_),
    .Y(_3673_)
);

NOR2X1 _14620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3673_),
    .B(_3671_),
    .Y(_3674_)
);

NAND2X1 _14621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3674_),
    .B(_3669_),
    .Y(_3675_)
);

INVX4 _14622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3675__bF$buf4),
    .Y(_3676_)
);

NAND2X1 _14623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [0]),
    .B(_3676_),
    .Y(_3677_)
);

NOR2X1 _14624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [27]),
    .B(\datapath.idinstr [26]),
    .Y(_3678_)
);

NAND2X1 _14625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3667_),
    .B(_3678_),
    .Y(_3679_)
);

NOR2X1 _14626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3679_),
    .B(_3665_),
    .Y(_3680_)
);

OR2X2 _14627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3672_),
    .B(\datapath.idinstr_21_bF$buf42 ),
    .Y(_3681_)
);

INVX1 _14628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_23_bF$buf5 ),
    .Y(_3682_)
);

NAND2X1 _14629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf41 ),
    .B(_3682_),
    .Y(_3683_)
);

NOR2X1 _14630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3683_),
    .B(_3681_),
    .Y(_3684_)
);

AND2X2 _14631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3680_),
    .B(_3684_),
    .Y(_3685_)
);

INVX1 _14632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf4),
    .Y(_3686_)
);

OAI21X1 _14633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3247_),
    .B(_3686_),
    .C(_3677_),
    .Y(\datapath.csr.csr_data [0])
);

NAND2X1 _14634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [1]),
    .B(_3676_),
    .Y(_3687_)
);

OAI21X1 _14635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3269_),
    .B(_3686_),
    .C(_3687_),
    .Y(\datapath.csr.csr_data [1])
);

INVX1 _14636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [2]),
    .Y(_3688_)
);

NOR2X1 _14637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3671_),
    .B(_3681_),
    .Y(_3689_)
);

AND2X2 _14638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3669_),
    .B(_3689_),
    .Y(_3690_)
);

AOI22X1 _14639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf3),
    .B(\datapath.csr.mvect [2]),
    .C(\datapath.csr.mepc [0]),
    .D(_3690__bF$buf4),
    .Y(_3691_)
);

OAI21X1 _14640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3688_),
    .B(_3675__bF$buf3),
    .C(_3691_),
    .Y(\datapath.csr.csr_data [2])
);

NOR2X1 _14641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf41 ),
    .B(\datapath.idinstr_20_bF$buf53 ),
    .Y(_3692_)
);

AND2X2 _14642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3680_),
    .B(_3670_),
    .Y(_3693_)
);

NAND2X1 _14643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3692_),
    .B(_3693_),
    .Y(_3694_)
);

NAND2X1 _14644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [3]),
    .B(_3676_),
    .Y(_3695_)
);

AOI22X1 _14645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf2),
    .B(\datapath.csr.mvect [3]),
    .C(\datapath.csr.mepc [1]),
    .D(_3690__bF$buf3),
    .Y(_3696_)
);

AND2X2 _14646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3695_),
    .B(_3696_),
    .Y(_3697_)
);

OAI21X1 _14647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3522_),
    .B(_3694_),
    .C(_3697_),
    .Y(\datapath.csr.csr_data [3])
);

AOI22X1 _14648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf1),
    .B(\datapath.csr.mvect [4]),
    .C(\datapath.csr.mepc [2]),
    .D(_3690__bF$buf2),
    .Y(_3698_)
);

OAI21X1 _14649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3459_),
    .B(_3675__bF$buf2),
    .C(_3698_),
    .Y(\datapath.csr.csr_data [4])
);

AOI22X1 _14650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf0),
    .B(\datapath.csr.mvect [5]),
    .C(\datapath.csr.mepc [3]),
    .D(_3690__bF$buf1),
    .Y(_3699_)
);

OAI21X1 _14651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3465_),
    .B(_3675__bF$buf1),
    .C(_3699_),
    .Y(\datapath.csr.csr_data [5])
);

AOI22X1 _14652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf4),
    .B(\datapath.csr.mvect [6]),
    .C(\datapath.csr.mepc [4]),
    .D(_3690__bF$buf0),
    .Y(_3700_)
);

OAI21X1 _14653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3467_),
    .B(_3675__bF$buf0),
    .C(_3700_),
    .Y(\datapath.csr.csr_data [6])
);

INVX1 _14654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3694_),
    .Y(_3701_)
);

NAND2X1 _14655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mstatus [1]),
    .B(_3701_),
    .Y(_3702_)
);

NAND2X1 _14656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [7]),
    .B(_3676_),
    .Y(_3703_)
);

AOI22X1 _14657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf3),
    .B(\datapath.csr.mvect [7]),
    .C(\datapath.csr.mepc [5]),
    .D(_3690__bF$buf4),
    .Y(_3704_)
);

NAND3X1 _14658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3703_),
    .B(_3704_),
    .C(_3702_),
    .Y(\datapath.csr.csr_data [7])
);

AOI22X1 _14659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [6]),
    .B(_3690__bF$buf3),
    .C(_3676_),
    .D(\datapath.csr.mcause [8]),
    .Y(_3705_)
);

NAND2X1 _14660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [8]),
    .B(_3685__bF$buf2),
    .Y(_3706_)
);

INVX1 _14661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3681_),
    .Y(_3707_)
);

NAND2X1 _14662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3707_),
    .B(_3693_),
    .Y(_3708_)
);

NAND3X1 _14663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3706_),
    .B(_3708_),
    .C(_3705_),
    .Y(\datapath.csr.csr_data [8])
);

AOI22X1 _14664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf1),
    .B(\datapath.csr.mvect [9]),
    .C(\datapath.csr.mepc [7]),
    .D(_3690__bF$buf2),
    .Y(_3709_)
);

OAI21X1 _14665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3473_),
    .B(_3675__bF$buf4),
    .C(_3709_),
    .Y(\datapath.csr.csr_data [9])
);

AOI22X1 _14666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf0),
    .B(\datapath.csr.mvect [10]),
    .C(\datapath.csr.mepc [8]),
    .D(_3690__bF$buf1),
    .Y(_3710_)
);

OAI21X1 _14667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3475_),
    .B(_3675__bF$buf3),
    .C(_3710_),
    .Y(\datapath.csr.csr_data [10])
);

AOI21X1 _14668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [9]),
    .B(_3690__bF$buf0),
    .C(_3701_),
    .Y(_3711_)
);

INVX1 _14669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mip ),
    .Y(_3712_)
);

NOR2X1 _14670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3712_),
    .B(_3668_),
    .Y(_3713_)
);

INVX1 _14671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mie ),
    .Y(_3714_)
);

NOR2X1 _14672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3714_),
    .B(_3679_),
    .Y(_3715_)
);

NAND3X1 _14673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3682_),
    .B(\datapath.idinstr_22_bF$buf40 ),
    .C(_3692_),
    .Y(_3716_)
);

NOR2X1 _14674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3665_),
    .B(_3716_),
    .Y(_3717_)
);

OAI21X1 _14675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3713_),
    .B(_3715_),
    .C(_3717_),
    .Y(_3718_)
);

AOI22X1 _14676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [11]),
    .B(_3685__bF$buf4),
    .C(_3676_),
    .D(\datapath.csr.mcause [11]),
    .Y(_3719_)
);

NAND3X1 _14677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3718_),
    .B(_3719_),
    .C(_3711_),
    .Y(\datapath.csr.csr_data [11])
);

NAND2X1 _14678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [12]),
    .B(_3685__bF$buf3),
    .Y(_3720_)
);

AOI22X1 _14679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [10]),
    .B(_3690__bF$buf4),
    .C(_3676_),
    .D(\datapath.csr.mcause [12]),
    .Y(_3721_)
);

NAND3X1 _14680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3694_),
    .B(_3720_),
    .C(_3721_),
    .Y(\datapath.csr.csr_data [12])
);

AOI22X1 _14681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf2),
    .B(\datapath.csr.mvect [13]),
    .C(\datapath.csr.mepc [11]),
    .D(_3690__bF$buf3),
    .Y(_3722_)
);

OAI21X1 _14682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3481_),
    .B(_3675__bF$buf2),
    .C(_3722_),
    .Y(\datapath.csr.csr_data [13])
);

AOI22X1 _14683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf1),
    .B(\datapath.csr.mvect [14]),
    .C(\datapath.csr.mepc [12]),
    .D(_3690__bF$buf2),
    .Y(_3723_)
);

OAI21X1 _14684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3483_),
    .B(_3675__bF$buf1),
    .C(_3723_),
    .Y(\datapath.csr.csr_data [14])
);

AOI22X1 _14685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf0),
    .B(\datapath.csr.mvect [15]),
    .C(\datapath.csr.mepc [13]),
    .D(_3690__bF$buf1),
    .Y(_3724_)
);

OAI21X1 _14686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3485_),
    .B(_3675__bF$buf0),
    .C(_3724_),
    .Y(\datapath.csr.csr_data [15])
);

AOI22X1 _14687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf4),
    .B(\datapath.csr.mvect [16]),
    .C(\datapath.csr.mepc [14]),
    .D(_3690__bF$buf0),
    .Y(_3725_)
);

OAI21X1 _14688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3487_),
    .B(_3675__bF$buf4),
    .C(_3725_),
    .Y(\datapath.csr.csr_data [16])
);

AOI22X1 _14689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf3),
    .B(\datapath.csr.mvect [17]),
    .C(\datapath.csr.mepc [15]),
    .D(_3690__bF$buf4),
    .Y(_3726_)
);

OAI21X1 _14690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3489_),
    .B(_3675__bF$buf3),
    .C(_3726_),
    .Y(\datapath.csr.csr_data [17])
);

AOI22X1 _14691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf2),
    .B(\datapath.csr.mvect [18]),
    .C(\datapath.csr.mepc [16]),
    .D(_3690__bF$buf3),
    .Y(_3727_)
);

OAI21X1 _14692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3491_),
    .B(_3675__bF$buf2),
    .C(_3727_),
    .Y(\datapath.csr.csr_data [18])
);

AOI22X1 _14693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf1),
    .B(\datapath.csr.mvect [19]),
    .C(\datapath.csr.mepc [17]),
    .D(_3690__bF$buf2),
    .Y(_3728_)
);

OAI21X1 _14694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3493_),
    .B(_3675__bF$buf1),
    .C(_3728_),
    .Y(\datapath.csr.csr_data [19])
);

AOI22X1 _14695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf0),
    .B(\datapath.csr.mvect [20]),
    .C(\datapath.csr.mepc [18]),
    .D(_3690__bF$buf1),
    .Y(_3729_)
);

OAI21X1 _14696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3495_),
    .B(_3675__bF$buf0),
    .C(_3729_),
    .Y(\datapath.csr.csr_data [20])
);

AOI22X1 _14697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf4),
    .B(\datapath.csr.mvect [21]),
    .C(\datapath.csr.mepc [19]),
    .D(_3690__bF$buf0),
    .Y(_3730_)
);

OAI21X1 _14698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3497_),
    .B(_3675__bF$buf4),
    .C(_3730_),
    .Y(\datapath.csr.csr_data [21])
);

AOI22X1 _14699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf3),
    .B(\datapath.csr.mvect [22]),
    .C(\datapath.csr.mepc [20]),
    .D(_3690__bF$buf4),
    .Y(_3731_)
);

OAI21X1 _14700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3499_),
    .B(_3675__bF$buf3),
    .C(_3731_),
    .Y(\datapath.csr.csr_data [22])
);

AOI22X1 _14701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf2),
    .B(\datapath.csr.mvect [23]),
    .C(\datapath.csr.mepc [21]),
    .D(_3690__bF$buf3),
    .Y(_3732_)
);

OAI21X1 _14702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3501_),
    .B(_3675__bF$buf2),
    .C(_3732_),
    .Y(\datapath.csr.csr_data [23])
);

AOI22X1 _14703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf1),
    .B(\datapath.csr.mvect [24]),
    .C(\datapath.csr.mepc [22]),
    .D(_3690__bF$buf2),
    .Y(_3733_)
);

OAI21X1 _14704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3503_),
    .B(_3675__bF$buf1),
    .C(_3733_),
    .Y(\datapath.csr.csr_data [24])
);

AOI22X1 _14705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf0),
    .B(\datapath.csr.mvect [25]),
    .C(\datapath.csr.mepc [23]),
    .D(_3690__bF$buf1),
    .Y(_3734_)
);

OAI21X1 _14706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3505_),
    .B(_3675__bF$buf0),
    .C(_3734_),
    .Y(\datapath.csr.csr_data [25])
);

AOI22X1 _14707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf4),
    .B(\datapath.csr.mvect [26]),
    .C(\datapath.csr.mepc [24]),
    .D(_3690__bF$buf0),
    .Y(_3735_)
);

OAI21X1 _14708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3507_),
    .B(_3675__bF$buf4),
    .C(_3735_),
    .Y(\datapath.csr.csr_data [26])
);

AOI22X1 _14709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf3),
    .B(\datapath.csr.mvect [27]),
    .C(\datapath.csr.mepc [25]),
    .D(_3690__bF$buf4),
    .Y(_3736_)
);

OAI21X1 _14710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3509_),
    .B(_3675__bF$buf3),
    .C(_3736_),
    .Y(\datapath.csr.csr_data [27])
);

AOI22X1 _14711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf2),
    .B(\datapath.csr.mvect [28]),
    .C(\datapath.csr.mepc [26]),
    .D(_3690__bF$buf3),
    .Y(_3737_)
);

OAI21X1 _14712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3511_),
    .B(_3675__bF$buf2),
    .C(_3737_),
    .Y(\datapath.csr.csr_data [28])
);

AOI22X1 _14713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf1),
    .B(\datapath.csr.mvect [29]),
    .C(\datapath.csr.mepc [27]),
    .D(_3690__bF$buf2),
    .Y(_3242_)
);

OAI21X1 _14714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3513_),
    .B(_3675__bF$buf1),
    .C(_3242_),
    .Y(\datapath.csr.csr_data [29])
);

NAND2X1 _14715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mvect [30]),
    .B(_3685__bF$buf0),
    .Y(_3243_)
);

AOI22X1 _14716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mepc [28]),
    .B(_3690__bF$buf1),
    .C(_3676_),
    .D(\datapath.csr.mcause [30]),
    .Y(_3244_)
);

NAND3X1 _14717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3708_),
    .B(_3243_),
    .C(_3244_),
    .Y(\datapath.csr.csr_data [30])
);

INVX1 _14718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.mcause [31]),
    .Y(_3245_)
);

AOI22X1 _14719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685__bF$buf4),
    .B(\datapath.csr.mvect [31]),
    .C(\datapath.csr.mepc [29]),
    .D(_3690__bF$buf0),
    .Y(_3246_)
);

OAI21X1 _14720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3245_),
    .B(_3675__bF$buf0),
    .C(_3246_),
    .Y(\datapath.csr.csr_data [31])
);

DFFPOSX1 _14721_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf1),
    .D(\datapath.csr._37_ [0]),
    .Q(\datapath.csr.mstatus [0])
);

DFFPOSX1 _14722_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf0),
    .D(\datapath.csr._37_ [1]),
    .Q(\datapath.csr.mstatus [1])
);

DFFPOSX1 _14723_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf153),
    .D(\datapath.csr._32_ [0]),
    .Q(\datapath.csr.mcause [0])
);

DFFPOSX1 _14724_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf152),
    .D(\datapath.csr._32_ [1]),
    .Q(\datapath.csr.mcause [1])
);

DFFPOSX1 _14725_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf151),
    .D(\datapath.csr._32_ [2]),
    .Q(\datapath.csr.mcause [2])
);

DFFPOSX1 _14726_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf150),
    .D(\datapath.csr._32_ [3]),
    .Q(\datapath.csr.mcause [3])
);

DFFPOSX1 _14727_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf149),
    .D(\datapath.csr._32_ [4]),
    .Q(\datapath.csr.mcause [4])
);

DFFPOSX1 _14728_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf148),
    .D(\datapath.csr._32_ [5]),
    .Q(\datapath.csr.mcause [5])
);

DFFPOSX1 _14729_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf147),
    .D(\datapath.csr._32_ [6]),
    .Q(\datapath.csr.mcause [6])
);

DFFPOSX1 _14730_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf146),
    .D(\datapath.csr._32_ [7]),
    .Q(\datapath.csr.mcause [7])
);

DFFPOSX1 _14731_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf145),
    .D(\datapath.csr._32_ [8]),
    .Q(\datapath.csr.mcause [8])
);

DFFPOSX1 _14732_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf144),
    .D(\datapath.csr._32_ [9]),
    .Q(\datapath.csr.mcause [9])
);

DFFPOSX1 _14733_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf143),
    .D(\datapath.csr._32_ [10]),
    .Q(\datapath.csr.mcause [10])
);

DFFPOSX1 _14734_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf142),
    .D(\datapath.csr._32_ [11]),
    .Q(\datapath.csr.mcause [11])
);

DFFPOSX1 _14735_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf141),
    .D(\datapath.csr._32_ [12]),
    .Q(\datapath.csr.mcause [12])
);

DFFPOSX1 _14736_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf140),
    .D(\datapath.csr._32_ [13]),
    .Q(\datapath.csr.mcause [13])
);

DFFPOSX1 _14737_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf139),
    .D(\datapath.csr._32_ [14]),
    .Q(\datapath.csr.mcause [14])
);

DFFPOSX1 _14738_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf138),
    .D(\datapath.csr._32_ [15]),
    .Q(\datapath.csr.mcause [15])
);

DFFPOSX1 _14739_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf137),
    .D(\datapath.csr._32_ [16]),
    .Q(\datapath.csr.mcause [16])
);

DFFPOSX1 _14740_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf136),
    .D(\datapath.csr._32_ [17]),
    .Q(\datapath.csr.mcause [17])
);

DFFPOSX1 _14741_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf135),
    .D(\datapath.csr._32_ [18]),
    .Q(\datapath.csr.mcause [18])
);

DFFPOSX1 _14742_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf134),
    .D(\datapath.csr._32_ [19]),
    .Q(\datapath.csr.mcause [19])
);

DFFPOSX1 _14743_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf133),
    .D(\datapath.csr._32_ [20]),
    .Q(\datapath.csr.mcause [20])
);

DFFPOSX1 _14744_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf132),
    .D(\datapath.csr._32_ [21]),
    .Q(\datapath.csr.mcause [21])
);

DFFPOSX1 _14745_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf131),
    .D(\datapath.csr._32_ [22]),
    .Q(\datapath.csr.mcause [22])
);

DFFPOSX1 _14746_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf130),
    .D(\datapath.csr._32_ [23]),
    .Q(\datapath.csr.mcause [23])
);

DFFPOSX1 _14747_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf129),
    .D(\datapath.csr._32_ [24]),
    .Q(\datapath.csr.mcause [24])
);

DFFPOSX1 _14748_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf128),
    .D(\datapath.csr._32_ [25]),
    .Q(\datapath.csr.mcause [25])
);

DFFPOSX1 _14749_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf127),
    .D(\datapath.csr._32_ [26]),
    .Q(\datapath.csr.mcause [26])
);

DFFPOSX1 _14750_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf126),
    .D(\datapath.csr._32_ [27]),
    .Q(\datapath.csr.mcause [27])
);

DFFPOSX1 _14751_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf125),
    .D(\datapath.csr._32_ [28]),
    .Q(\datapath.csr.mcause [28])
);

DFFPOSX1 _14752_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf124),
    .D(\datapath.csr._32_ [29]),
    .Q(\datapath.csr.mcause [29])
);

DFFPOSX1 _14753_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf123),
    .D(\datapath.csr._32_ [30]),
    .Q(\datapath.csr.mcause [30])
);

DFFPOSX1 _14754_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf122),
    .D(\datapath.csr._32_ [31]),
    .Q(\datapath.csr.mcause [31])
);

DFFPOSX1 _14755_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf121),
    .D(\datapath.csr._26_ [0]),
    .Q(\datapath.csr.mepc [0])
);

DFFPOSX1 _14756_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf120),
    .D(\datapath.csr._26_ [1]),
    .Q(\datapath.csr.mepc [1])
);

DFFPOSX1 _14757_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf119),
    .D(\datapath.csr._26_ [2]),
    .Q(\datapath.csr.mepc [2])
);

DFFPOSX1 _14758_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf118),
    .D(\datapath.csr._26_ [3]),
    .Q(\datapath.csr.mepc [3])
);

DFFPOSX1 _14759_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf117),
    .D(\datapath.csr._26_ [4]),
    .Q(\datapath.csr.mepc [4])
);

DFFPOSX1 _14760_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf116),
    .D(\datapath.csr._26_ [5]),
    .Q(\datapath.csr.mepc [5])
);

DFFPOSX1 _14761_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf115),
    .D(\datapath.csr._26_ [6]),
    .Q(\datapath.csr.mepc [6])
);

DFFPOSX1 _14762_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf114),
    .D(\datapath.csr._26_ [7]),
    .Q(\datapath.csr.mepc [7])
);

DFFPOSX1 _14763_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf113),
    .D(\datapath.csr._26_ [8]),
    .Q(\datapath.csr.mepc [8])
);

DFFPOSX1 _14764_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf112),
    .D(\datapath.csr._26_ [9]),
    .Q(\datapath.csr.mepc [9])
);

DFFPOSX1 _14765_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf111),
    .D(\datapath.csr._26_ [10]),
    .Q(\datapath.csr.mepc [10])
);

DFFPOSX1 _14766_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf110),
    .D(\datapath.csr._26_ [11]),
    .Q(\datapath.csr.mepc [11])
);

DFFPOSX1 _14767_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf109),
    .D(\datapath.csr._26_ [12]),
    .Q(\datapath.csr.mepc [12])
);

DFFPOSX1 _14768_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf108),
    .D(\datapath.csr._26_ [13]),
    .Q(\datapath.csr.mepc [13])
);

DFFPOSX1 _14769_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf107),
    .D(\datapath.csr._26_ [14]),
    .Q(\datapath.csr.mepc [14])
);

DFFPOSX1 _14770_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf106),
    .D(\datapath.csr._26_ [15]),
    .Q(\datapath.csr.mepc [15])
);

DFFPOSX1 _14771_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf105),
    .D(\datapath.csr._26_ [16]),
    .Q(\datapath.csr.mepc [16])
);

DFFPOSX1 _14772_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf104),
    .D(\datapath.csr._26_ [17]),
    .Q(\datapath.csr.mepc [17])
);

DFFPOSX1 _14773_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf103),
    .D(\datapath.csr._26_ [18]),
    .Q(\datapath.csr.mepc [18])
);

DFFPOSX1 _14774_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf102),
    .D(\datapath.csr._26_ [19]),
    .Q(\datapath.csr.mepc [19])
);

DFFPOSX1 _14775_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf101),
    .D(\datapath.csr._26_ [20]),
    .Q(\datapath.csr.mepc [20])
);

DFFPOSX1 _14776_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf100),
    .D(\datapath.csr._26_ [21]),
    .Q(\datapath.csr.mepc [21])
);

DFFPOSX1 _14777_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf99),
    .D(\datapath.csr._26_ [22]),
    .Q(\datapath.csr.mepc [22])
);

DFFPOSX1 _14778_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf98),
    .D(\datapath.csr._26_ [23]),
    .Q(\datapath.csr.mepc [23])
);

DFFPOSX1 _14779_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf97),
    .D(\datapath.csr._26_ [24]),
    .Q(\datapath.csr.mepc [24])
);

DFFPOSX1 _14780_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf96),
    .D(\datapath.csr._26_ [25]),
    .Q(\datapath.csr.mepc [25])
);

DFFPOSX1 _14781_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf95),
    .D(\datapath.csr._26_ [26]),
    .Q(\datapath.csr.mepc [26])
);

DFFPOSX1 _14782_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf94),
    .D(\datapath.csr._26_ [27]),
    .Q(\datapath.csr.mepc [27])
);

DFFPOSX1 _14783_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf93),
    .D(\datapath.csr._26_ [28]),
    .Q(\datapath.csr.mepc [28])
);

DFFPOSX1 _14784_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf92),
    .D(\datapath.csr._26_ [29]),
    .Q(\datapath.csr.mepc [29])
);

DFFPOSX1 _14785_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf91),
    .D(IRQ),
    .Q(\datapath.csr.meta_irq )
);

DFFPOSX1 _14786_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf90),
    .D(\datapath.csr.meta_irq ),
    .Q(\datapath.csr.mip )
);

DFFPOSX1 _14787_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf89),
    .D(\datapath.csr._20_ ),
    .Q(\datapath.csr.mie )
);

DFFPOSX1 _14788_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf88),
    .D(\datapath.csr._13_ [0]),
    .Q(\datapath.csr.mvect [0])
);

DFFPOSX1 _14789_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf87),
    .D(\datapath.csr._13_ [1]),
    .Q(\datapath.csr.mvect [1])
);

DFFPOSX1 _14790_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf86),
    .D(\datapath.csr._13_ [2]),
    .Q(\datapath.csr.mvect [2])
);

DFFPOSX1 _14791_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf85),
    .D(\datapath.csr._13_ [3]),
    .Q(\datapath.csr.mvect [3])
);

DFFPOSX1 _14792_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf84),
    .D(\datapath.csr._13_ [4]),
    .Q(\datapath.csr.mvect [4])
);

DFFPOSX1 _14793_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf83),
    .D(\datapath.csr._13_ [5]),
    .Q(\datapath.csr.mvect [5])
);

DFFPOSX1 _14794_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf82),
    .D(\datapath.csr._13_ [6]),
    .Q(\datapath.csr.mvect [6])
);

DFFPOSX1 _14795_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf81),
    .D(\datapath.csr._13_ [7]),
    .Q(\datapath.csr.mvect [7])
);

DFFPOSX1 _14796_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf80),
    .D(\datapath.csr._13_ [8]),
    .Q(\datapath.csr.mvect [8])
);

DFFPOSX1 _14797_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf79),
    .D(\datapath.csr._13_ [9]),
    .Q(\datapath.csr.mvect [9])
);

DFFPOSX1 _14798_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf78),
    .D(\datapath.csr._13_ [10]),
    .Q(\datapath.csr.mvect [10])
);

DFFPOSX1 _14799_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf77),
    .D(\datapath.csr._13_ [11]),
    .Q(\datapath.csr.mvect [11])
);

DFFPOSX1 _14800_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf76),
    .D(\datapath.csr._13_ [12]),
    .Q(\datapath.csr.mvect [12])
);

DFFPOSX1 _14801_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf75),
    .D(\datapath.csr._13_ [13]),
    .Q(\datapath.csr.mvect [13])
);

DFFPOSX1 _14802_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf74),
    .D(\datapath.csr._13_ [14]),
    .Q(\datapath.csr.mvect [14])
);

DFFPOSX1 _14803_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf73),
    .D(\datapath.csr._13_ [15]),
    .Q(\datapath.csr.mvect [15])
);

DFFPOSX1 _14804_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf72),
    .D(\datapath.csr._13_ [16]),
    .Q(\datapath.csr.mvect [16])
);

DFFPOSX1 _14805_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf71),
    .D(\datapath.csr._13_ [17]),
    .Q(\datapath.csr.mvect [17])
);

DFFPOSX1 _14806_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf70),
    .D(\datapath.csr._13_ [18]),
    .Q(\datapath.csr.mvect [18])
);

DFFPOSX1 _14807_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf69),
    .D(\datapath.csr._13_ [19]),
    .Q(\datapath.csr.mvect [19])
);

DFFPOSX1 _14808_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf68),
    .D(\datapath.csr._13_ [20]),
    .Q(\datapath.csr.mvect [20])
);

DFFPOSX1 _14809_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf67),
    .D(\datapath.csr._13_ [21]),
    .Q(\datapath.csr.mvect [21])
);

DFFPOSX1 _14810_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf66),
    .D(\datapath.csr._13_ [22]),
    .Q(\datapath.csr.mvect [22])
);

DFFPOSX1 _14811_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf65),
    .D(\datapath.csr._13_ [23]),
    .Q(\datapath.csr.mvect [23])
);

DFFPOSX1 _14812_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf64),
    .D(\datapath.csr._13_ [24]),
    .Q(\datapath.csr.mvect [24])
);

DFFPOSX1 _14813_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf63),
    .D(\datapath.csr._13_ [25]),
    .Q(\datapath.csr.mvect [25])
);

DFFPOSX1 _14814_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf62),
    .D(\datapath.csr._13_ [26]),
    .Q(\datapath.csr.mvect [26])
);

DFFPOSX1 _14815_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf61),
    .D(\datapath.csr._13_ [27]),
    .Q(\datapath.csr.mvect [27])
);

DFFPOSX1 _14816_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf60),
    .D(\datapath.csr._13_ [28]),
    .Q(\datapath.csr.mvect [28])
);

DFFPOSX1 _14817_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf59),
    .D(\datapath.csr._13_ [29]),
    .Q(\datapath.csr.mvect [29])
);

DFFPOSX1 _14818_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf58),
    .D(\datapath.csr._13_ [30]),
    .Q(\datapath.csr.mvect [30])
);

DFFPOSX1 _14819_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf57),
    .D(\datapath.csr._13_ [31]),
    .Q(\datapath.csr.mvect [31])
);

INVX2 _14820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.imm_sel [2]),
    .Y(_3774_)
);

INVX2 _14821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.imm_sel [1]),
    .Y(_3775_)
);

NAND2X1 _14822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.imm_sel [0]),
    .B(_3775_),
    .Y(_3776_)
);

OAI21X1 _14823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3776_),
    .B(_3774_),
    .C(\datapath.idinstr [31]),
    .Y(_3777_)
);

INVX1 _14824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3777_),
    .Y(\datapath.immediatedecoder._12_ )
);

INVX1 _14825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [25]),
    .Y(_3778_)
);

NAND3X1 _14826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.imm_sel [1]),
    .B(\controlunit.imm_sel [0]),
    .C(_3774_),
    .Y(_3779_)
);

OAI21X1 _14827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3776_),
    .B(_3774_),
    .C(_3779_),
    .Y(_3780_)
);

NOR2X1 _14828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3778_),
    .B(_3780_),
    .Y(\datapath.imm [5])
);

INVX1 _14829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [26]),
    .Y(_3781_)
);

NOR2X1 _14830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .B(_3780_),
    .Y(\datapath.imm [6])
);

INVX1 _14831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [27]),
    .Y(_3782_)
);

NOR2X1 _14832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3782_),
    .B(_3780_),
    .Y(\datapath.imm [7])
);

INVX1 _14833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [28]),
    .Y(_3783_)
);

NOR2X1 _14834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3783_),
    .B(_3780_),
    .Y(\datapath.imm [8])
);

INVX1 _14835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [29]),
    .Y(_3784_)
);

NOR2X1 _14836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3784_),
    .B(_3780_),
    .Y(\datapath.imm [9])
);

INVX1 _14837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [30]),
    .Y(_3785_)
);

NOR2X1 _14838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3785_),
    .B(_3780_),
    .Y(\datapath.imm [10])
);

INVX1 _14839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf52 ),
    .Y(_3786_)
);

NOR2X1 _14840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.imm_sel [1]),
    .B(\controlunit.imm_sel [0]),
    .Y(_3787_)
);

AOI21X1 _14841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.imm_sel [1]),
    .B(\controlunit.imm_sel [0]),
    .C(\controlunit.imm_sel [2]),
    .Y(_3788_)
);

OAI21X1 _14842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3788_),
    .B(_3787_),
    .C(\datapath.idinstr [31]),
    .Y(_3789_)
);

OAI21X1 _14843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.imm_sel [0]),
    .B(\controlunit.imm_sel [2]),
    .C(\controlunit.imm_sel [1]),
    .Y(_3790_)
);

OAI21X1 _14844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3786_),
    .B(_3790_),
    .C(_3789_),
    .Y(\datapath.imm [20])
);

INVX1 _14845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf40 ),
    .Y(_3791_)
);

OAI21X1 _14846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3791_),
    .B(_3790_),
    .C(_3789_),
    .Y(\datapath.imm [21])
);

INVX1 _14847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf39 ),
    .Y(_3792_)
);

OAI21X1 _14848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3792_),
    .B(_3790_),
    .C(_3789_),
    .Y(\datapath.imm [22])
);

INVX1 _14849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_23_bF$buf4 ),
    .Y(_3793_)
);

OAI21X1 _14850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3793_),
    .B(_3790_),
    .C(_3789_),
    .Y(\datapath.imm [23])
);

INVX1 _14851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_24_bF$buf3 ),
    .Y(_3794_)
);

OAI21X1 _14852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3794_),
    .B(_3790_),
    .C(_3789_),
    .Y(\datapath.imm [24])
);

OAI21X1 _14853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3778_),
    .B(_3790_),
    .C(_3789_),
    .Y(\datapath.imm [25])
);

OAI21X1 _14854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .B(_3790_),
    .C(_3789_),
    .Y(\datapath.imm [26])
);

OAI21X1 _14855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3782_),
    .B(_3790_),
    .C(_3789_),
    .Y(\datapath.imm [27])
);

OAI21X1 _14856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3783_),
    .B(_3790_),
    .C(_3789_),
    .Y(\datapath.imm [28])
);

OAI21X1 _14857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3784_),
    .B(_3790_),
    .C(_3789_),
    .Y(\datapath.imm [29])
);

OAI21X1 _14858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3785_),
    .B(_3790_),
    .C(_3789_),
    .Y(\datapath.imm [30])
);

INVX2 _14859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.imm_sel [0]),
    .Y(_3738_)
);

NAND2X1 _14860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3775_),
    .B(_3738_),
    .Y(_3739_)
);

OAI21X1 _14861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3739_),
    .B(_3774_),
    .C(_3779_),
    .Y(_3740_)
);

INVX4 _14862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3788_),
    .Y(_3741_)
);

OAI21X1 _14863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.imm_sel [1]),
    .B(\controlunit.imm_sel [0]),
    .C(\controlunit.imm_sel [2]),
    .Y(_3742_)
);

NAND3X1 _14864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [12]),
    .B(_3742_),
    .C(_3741_),
    .Y(_3743_)
);

OAI21X1 _14865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3740_),
    .B(_3777_),
    .C(_3743_),
    .Y(\datapath.imm [12])
);

NAND3X1 _14866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [13]),
    .B(_3742_),
    .C(_3741_),
    .Y(_3744_)
);

OAI21X1 _14867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3740_),
    .B(_3777_),
    .C(_3744_),
    .Y(\datapath.imm [13])
);

NAND3X1 _14868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [14]),
    .B(_3742_),
    .C(_3741_),
    .Y(_3745_)
);

OAI21X1 _14869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3740_),
    .B(_3777_),
    .C(_3745_),
    .Y(\datapath.imm [14])
);

NAND3X1 _14870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf52 ),
    .B(_3742_),
    .C(_3741_),
    .Y(_3746_)
);

OAI21X1 _14871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3740_),
    .B(_3777_),
    .C(_3746_),
    .Y(\datapath.imm [15])
);

NAND3X1 _14872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_bF$buf44 ),
    .B(_3742_),
    .C(_3741_),
    .Y(_3747_)
);

OAI21X1 _14873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3740_),
    .B(_3777_),
    .C(_3747_),
    .Y(\datapath.imm [16])
);

NAND3X1 _14874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf40 ),
    .B(_3742_),
    .C(_3741_),
    .Y(_3748_)
);

OAI21X1 _14875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3740_),
    .B(_3777_),
    .C(_3748_),
    .Y(\datapath.imm [17])
);

NAND3X1 _14876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_18_bF$buf6 ),
    .B(_3742_),
    .C(_3741_),
    .Y(_3749_)
);

OAI21X1 _14877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3740_),
    .B(_3777_),
    .C(_3749_),
    .Y(\datapath.imm [18])
);

NAND3X1 _14878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_19_bF$buf4 ),
    .B(_3742_),
    .C(_3741_),
    .Y(_3750_)
);

OAI21X1 _14879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3740_),
    .B(_3777_),
    .C(_3750_),
    .Y(\datapath.imm [19])
);

NAND2X1 _14880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.imm_sel [1]),
    .B(_3774_),
    .Y(_3751_)
);

NAND2X1 _14881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.imm_sel [2]),
    .B(_3775_),
    .Y(_3752_)
);

NAND3X1 _14882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [31]),
    .B(_3751_),
    .C(_3752_),
    .Y(_3753_)
);

NAND3X1 _14883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.imm_sel [2]),
    .B(\datapath.idinstr_20_bF$buf51 ),
    .C(_3787_),
    .Y(_3754_)
);

NOR2X1 _14884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.imm_sel [2]),
    .B(_3775_),
    .Y(_3755_)
);

NAND3X1 _14885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3738_),
    .B(\datapath.idinstr [7]),
    .C(_3755_),
    .Y(_3756_)
);

NAND3X1 _14886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3753_),
    .B(_3754_),
    .C(_3756_),
    .Y(\datapath.immediatedecoder._09_ )
);

OAI21X1 _14887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3738_),
    .B(\controlunit.imm_sel [2]),
    .C(_3775_),
    .Y(_3757_)
);

NAND3X1 _14888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [8]),
    .B(_3779_),
    .C(_3757_),
    .Y(_3758_)
);

NAND2X1 _14889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf39 ),
    .B(_3787_),
    .Y(_3759_)
);

NOR2X1 _14890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.imm_sel [1]),
    .B(_3738_),
    .Y(_3760_)
);

NAND3X1 _14891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.imm_sel [2]),
    .B(\datapath.idinstr_16_bF$buf43 ),
    .C(_3760_),
    .Y(_3761_)
);

NAND3X1 _14892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3759_),
    .B(_3761_),
    .C(_3758_),
    .Y(\datapath.imm [1])
);

NAND3X1 _14893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [9]),
    .B(_3779_),
    .C(_3757_),
    .Y(_3762_)
);

NAND2X1 _14894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf38 ),
    .B(_3787_),
    .Y(_3763_)
);

NAND3X1 _14895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.imm_sel [2]),
    .B(\datapath.idinstr_17_bF$buf39 ),
    .C(_3760_),
    .Y(_3764_)
);

NAND3X1 _14896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3763_),
    .B(_3764_),
    .C(_3762_),
    .Y(\datapath.imm [2])
);

NAND3X1 _14897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [10]),
    .B(_3779_),
    .C(_3757_),
    .Y(_3765_)
);

NAND2X1 _14898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_23_bF$buf3 ),
    .B(_3787_),
    .Y(_3766_)
);

NAND3X1 _14899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.imm_sel [2]),
    .B(\datapath.idinstr_18_bF$buf5 ),
    .C(_3760_),
    .Y(_3767_)
);

NAND3X1 _14900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3766_),
    .B(_3767_),
    .C(_3765_),
    .Y(\datapath.imm [3])
);

NAND3X1 _14901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [11]),
    .B(_3779_),
    .C(_3757_),
    .Y(_3768_)
);

NAND2X1 _14902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_24_bF$buf2 ),
    .B(_3787_),
    .Y(_3769_)
);

NAND3X1 _14903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.imm_sel [2]),
    .B(\datapath.idinstr_19_bF$buf3 ),
    .C(_3760_),
    .Y(_3770_)
);

NAND3X1 _14904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3769_),
    .B(_3770_),
    .C(_3768_),
    .Y(\datapath.imm [4])
);

NAND2X1 _14905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3751_),
    .B(_3752_),
    .Y(_3771_)
);

MUX2X1 _14906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf51 ),
    .B(\datapath.idinstr [7]),
    .S(\controlunit.imm_sel [2]),
    .Y(_3772_)
);

OAI21X1 _14907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3738_),
    .B(\controlunit.imm_sel [1]),
    .C(\datapath.idinstr_20_bF$buf50 ),
    .Y(_3773_)
);

OAI22X1 _14908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3776_),
    .B(_3772_),
    .C(_3771_),
    .D(_3773_),
    .Y(\datapath.immediatedecoder._06_ )
);

INVX1 _14909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [12]),
    .Y(_3795_)
);

NAND2X1 _14910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [13]),
    .B(_3795_),
    .Y(_3796_)
);

INVX1 _14911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [13]),
    .Y(_3797_)
);

NAND2X1 _14912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [12]),
    .B(_3797_),
    .Y(_3798_)
);

NAND3X1 _14913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [0]),
    .B(_3796__bF$buf4),
    .C(_3798__bF$buf4),
    .Y(_3799_)
);

NOR2X1 _14914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [12]),
    .B(_3797_),
    .Y(_3800_)
);

NAND2X1 _14915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [0]),
    .B(_3800__bF$buf7),
    .Y(_3801_)
);

NOR2X1 _14916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [13]),
    .B(_3795_),
    .Y(_3802_)
);

INVX2 _14917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [0]),
    .Y(_3803_)
);

NAND2X1 _14918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[0]),
    .B(_0__1_bF$buf3),
    .Y(_3804_)
);

OAI21X1 _14919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3803_),
    .B(_0__1_bF$buf2),
    .C(_3804_),
    .Y(_3805_)
);

NAND2X1 _14920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf6),
    .B(_3805_),
    .Y(_3806_)
);

NAND3X1 _14921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3801_),
    .B(_3799_),
    .C(_3806_),
    .Y(_1_[0])
);

NAND3X1 _14922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [1]),
    .B(_3796__bF$buf3),
    .C(_3798__bF$buf3),
    .Y(_3807_)
);

NAND2X1 _14923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [1]),
    .B(_3800__bF$buf6),
    .Y(_3808_)
);

INVX2 _14924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [1]),
    .Y(_3809_)
);

NAND2X1 _14925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf1),
    .B(DMEM_DATA_L[1]),
    .Y(_3810_)
);

OAI21X1 _14926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3809_),
    .B(_0__1_bF$buf0),
    .C(_3810_),
    .Y(_3811_)
);

NAND2X1 _14927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf5),
    .B(_3811_),
    .Y(_3812_)
);

NAND3X1 _14928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3808_),
    .B(_3807_),
    .C(_3812_),
    .Y(_1_[1])
);

NAND3X1 _14929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [2]),
    .B(_3796__bF$buf2),
    .C(_3798__bF$buf2),
    .Y(_3813_)
);

NAND2X1 _14930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [2]),
    .B(_3800__bF$buf5),
    .Y(_3814_)
);

INVX2 _14931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [2]),
    .Y(_3815_)
);

NAND2X1 _14932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf9),
    .B(DMEM_DATA_L[2]),
    .Y(_3816_)
);

OAI21X1 _14933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3815_),
    .B(_0__1_bF$buf8),
    .C(_3816_),
    .Y(_3817_)
);

NAND2X1 _14934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf4),
    .B(_3817_),
    .Y(_3818_)
);

NAND3X1 _14935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3814_),
    .B(_3813_),
    .C(_3818_),
    .Y(_1_[2])
);

NAND3X1 _14936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [3]),
    .B(_3796__bF$buf1),
    .C(_3798__bF$buf1),
    .Y(_3819_)
);

NAND2X1 _14937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [3]),
    .B(_3800__bF$buf4),
    .Y(_3820_)
);

INVX2 _14938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [3]),
    .Y(_3821_)
);

NAND2X1 _14939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf7),
    .B(DMEM_DATA_L[3]),
    .Y(_3822_)
);

OAI21X1 _14940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3821_),
    .B(_0__1_bF$buf6),
    .C(_3822_),
    .Y(_3823_)
);

NAND2X1 _14941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf3),
    .B(_3823_),
    .Y(_3824_)
);

NAND3X1 _14942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3820_),
    .B(_3819_),
    .C(_3824_),
    .Y(_1_[3])
);

NAND3X1 _14943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [4]),
    .B(_3796__bF$buf0),
    .C(_3798__bF$buf0),
    .Y(_3825_)
);

NAND2X1 _14944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [4]),
    .B(_3800__bF$buf3),
    .Y(_3826_)
);

INVX2 _14945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [4]),
    .Y(_3827_)
);

NAND2X1 _14946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf5),
    .B(DMEM_DATA_L[4]),
    .Y(_3828_)
);

OAI21X1 _14947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3827_),
    .B(_0__1_bF$buf4),
    .C(_3828_),
    .Y(_3829_)
);

NAND2X1 _14948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf2),
    .B(_3829_),
    .Y(_3830_)
);

NAND3X1 _14949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3826_),
    .B(_3825_),
    .C(_3830_),
    .Y(_1_[4])
);

NAND3X1 _14950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [5]),
    .B(_3796__bF$buf4),
    .C(_3798__bF$buf4),
    .Y(_3831_)
);

NAND2X1 _14951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [5]),
    .B(_3800__bF$buf2),
    .Y(_3832_)
);

INVX2 _14952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [5]),
    .Y(_3833_)
);

NAND2X1 _14953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf3),
    .B(DMEM_DATA_L[5]),
    .Y(_3834_)
);

OAI21X1 _14954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3833_),
    .B(_0__1_bF$buf2),
    .C(_3834_),
    .Y(_3835_)
);

NAND2X1 _14955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf1),
    .B(_3835_),
    .Y(_3836_)
);

NAND3X1 _14956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3832_),
    .B(_3831_),
    .C(_3836_),
    .Y(_1_[5])
);

NAND3X1 _14957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [6]),
    .B(_3796__bF$buf3),
    .C(_3798__bF$buf3),
    .Y(_3837_)
);

NAND2X1 _14958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [6]),
    .B(_3800__bF$buf1),
    .Y(_3838_)
);

INVX2 _14959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [6]),
    .Y(_3839_)
);

NAND2X1 _14960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf1),
    .B(DMEM_DATA_L[6]),
    .Y(_3840_)
);

OAI21X1 _14961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3839_),
    .B(_0__1_bF$buf0),
    .C(_3840_),
    .Y(_3841_)
);

NAND2X1 _14962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf0),
    .B(_3841_),
    .Y(_3842_)
);

NAND3X1 _14963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3838_),
    .B(_3837_),
    .C(_3842_),
    .Y(_1_[6])
);

NAND3X1 _14964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [7]),
    .B(_3796__bF$buf2),
    .C(_3798__bF$buf2),
    .Y(_3843_)
);

NAND2X1 _14965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [7]),
    .B(_3800__bF$buf0),
    .Y(_3844_)
);

INVX2 _14966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [7]),
    .Y(_3845_)
);

NAND2X1 _14967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf9),
    .B(DMEM_DATA_L[7]),
    .Y(_3846_)
);

OAI21X1 _14968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3845_),
    .B(_0__1_bF$buf8),
    .C(_3846_),
    .Y(_3847_)
);

NAND2X1 _14969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf6),
    .B(_3847_),
    .Y(_3848_)
);

NAND3X1 _14970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3844_),
    .B(_3843_),
    .C(_3848_),
    .Y(_1_[7])
);

INVX1 _14971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [8]),
    .Y(_3849_)
);

NAND2X1 _14972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3796__bF$buf1),
    .B(_3798__bF$buf1),
    .Y(_3850_)
);

INVX1 _14973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [8]),
    .Y(_3851_)
);

NAND2X1 _14974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf7),
    .B(DMEM_DATA_L[8]),
    .Y(_3852_)
);

OAI21X1 _14975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3851_),
    .B(_0__1_bF$buf6),
    .C(_3852_),
    .Y(_3853_)
);

AOI22X1 _14976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [8]),
    .B(_3800__bF$buf7),
    .C(_3853_),
    .D(_3802__bF$buf5),
    .Y(_3854_)
);

OAI21X1 _14977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3849_),
    .B(_3850_),
    .C(_3854_),
    .Y(_1_[8])
);

INVX1 _14978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [9]),
    .Y(_3855_)
);

INVX1 _14979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [9]),
    .Y(_3856_)
);

NAND2X1 _14980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf5),
    .B(DMEM_DATA_L[9]),
    .Y(_3857_)
);

OAI21X1 _14981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3856_),
    .B(_0__1_bF$buf4),
    .C(_3857_),
    .Y(_3858_)
);

AOI22X1 _14982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [9]),
    .B(_3800__bF$buf6),
    .C(_3858_),
    .D(_3802__bF$buf4),
    .Y(_3859_)
);

OAI21X1 _14983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3855_),
    .B(_3850_),
    .C(_3859_),
    .Y(_1_[9])
);

INVX1 _14984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [10]),
    .Y(_3860_)
);

INVX1 _14985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [10]),
    .Y(_3861_)
);

NAND2X1 _14986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf3),
    .B(DMEM_DATA_L[10]),
    .Y(_3862_)
);

OAI21X1 _14987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3861_),
    .B(_0__1_bF$buf2),
    .C(_3862_),
    .Y(_3863_)
);

AOI22X1 _14988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [10]),
    .B(_3800__bF$buf5),
    .C(_3863_),
    .D(_3802__bF$buf3),
    .Y(_3864_)
);

OAI21X1 _14989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3860_),
    .B(_3850_),
    .C(_3864_),
    .Y(_1_[10])
);

INVX1 _14990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [11]),
    .Y(_3865_)
);

INVX1 _14991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [11]),
    .Y(_3866_)
);

NAND2X1 _14992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf1),
    .B(DMEM_DATA_L[11]),
    .Y(_3867_)
);

OAI21X1 _14993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3866_),
    .B(_0__1_bF$buf0),
    .C(_3867_),
    .Y(_3868_)
);

AOI22X1 _14994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [11]),
    .B(_3800__bF$buf4),
    .C(_3868_),
    .D(_3802__bF$buf2),
    .Y(_3869_)
);

OAI21X1 _14995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3865_),
    .B(_3850_),
    .C(_3869_),
    .Y(_1_[11])
);

INVX1 _14996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [12]),
    .Y(_3870_)
);

INVX1 _14997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [12]),
    .Y(_3871_)
);

NAND2X1 _14998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf9),
    .B(DMEM_DATA_L[12]),
    .Y(_3872_)
);

OAI21X1 _14999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3871_),
    .B(_0__1_bF$buf8),
    .C(_3872_),
    .Y(_3873_)
);

AOI22X1 _15000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [12]),
    .B(_3800__bF$buf3),
    .C(_3873_),
    .D(_3802__bF$buf1),
    .Y(_3874_)
);

OAI21X1 _15001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3870_),
    .B(_3850_),
    .C(_3874_),
    .Y(_1_[12])
);

INVX1 _15002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [13]),
    .Y(_3875_)
);

INVX1 _15003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [13]),
    .Y(_3876_)
);

NAND2X1 _15004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf7),
    .B(DMEM_DATA_L[13]),
    .Y(_3877_)
);

OAI21X1 _15005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3876_),
    .B(_0__1_bF$buf6),
    .C(_3877_),
    .Y(_3878_)
);

AOI22X1 _15006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [13]),
    .B(_3800__bF$buf2),
    .C(_3878_),
    .D(_3802__bF$buf0),
    .Y(_3879_)
);

OAI21X1 _15007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3875_),
    .B(_3850_),
    .C(_3879_),
    .Y(_1_[13])
);

INVX1 _15008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [14]),
    .Y(_3880_)
);

INVX1 _15009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [14]),
    .Y(_3881_)
);

NAND2X1 _15010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf5),
    .B(DMEM_DATA_L[14]),
    .Y(_3882_)
);

OAI21X1 _15011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3881_),
    .B(_0__1_bF$buf4),
    .C(_3882_),
    .Y(_3883_)
);

AOI22X1 _15012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [14]),
    .B(_3800__bF$buf1),
    .C(_3883_),
    .D(_3802__bF$buf6),
    .Y(_3884_)
);

OAI21X1 _15013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3880_),
    .B(_3850_),
    .C(_3884_),
    .Y(_1_[14])
);

INVX1 _15014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [15]),
    .Y(_3885_)
);

INVX1 _15015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [15]),
    .Y(_3886_)
);

NAND2X1 _15016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf3),
    .B(DMEM_DATA_L[15]),
    .Y(_3887_)
);

OAI21X1 _15017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3886_),
    .B(_0__1_bF$buf2),
    .C(_3887_),
    .Y(_3888_)
);

AOI22X1 _15018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [15]),
    .B(_3800__bF$buf0),
    .C(_3888_),
    .D(_3802__bF$buf5),
    .Y(_3889_)
);

OAI21X1 _15019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3885_),
    .B(_3850_),
    .C(_3889_),
    .Y(_1_[15])
);

INVX1 _15020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[16]),
    .Y(_3890_)
);

NAND2X1 _15021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [0]),
    .B(_0__1_bF$buf1),
    .Y(_3891_)
);

OAI21X1 _15022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3890_),
    .B(_0__1_bF$buf0),
    .C(_3891_),
    .Y(_3892_)
);

NAND2X1 _15023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf4),
    .B(_3892_),
    .Y(_3893_)
);

NAND3X1 _15024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [16]),
    .B(_3796__bF$buf0),
    .C(_3798__bF$buf0),
    .Y(_3894_)
);

NAND2X1 _15025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [16]),
    .B(_3800__bF$buf7),
    .Y(_3895_)
);

NAND3X1 _15026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3895_),
    .B(_3894_),
    .C(_3893_),
    .Y(_1_[16])
);

INVX1 _15027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[17]),
    .Y(_3896_)
);

NAND2X1 _15028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf9),
    .B(\datapath.memoryinterface.data_store [1]),
    .Y(_3897_)
);

OAI21X1 _15029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3896_),
    .B(_0__1_bF$buf8),
    .C(_3897_),
    .Y(_3898_)
);

NAND2X1 _15030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf3),
    .B(_3898_),
    .Y(_3899_)
);

NAND3X1 _15031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [17]),
    .B(_3796__bF$buf4),
    .C(_3798__bF$buf4),
    .Y(_3900_)
);

NAND2X1 _15032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [17]),
    .B(_3800__bF$buf6),
    .Y(_3901_)
);

NAND3X1 _15033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3901_),
    .B(_3900_),
    .C(_3899_),
    .Y(_1_[17])
);

INVX1 _15034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[18]),
    .Y(_3902_)
);

NAND2X1 _15035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf7),
    .B(\datapath.memoryinterface.data_store [2]),
    .Y(_3903_)
);

OAI21X1 _15036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3902_),
    .B(_0__1_bF$buf6),
    .C(_3903_),
    .Y(_3904_)
);

NAND2X1 _15037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf2),
    .B(_3904_),
    .Y(_3905_)
);

NAND3X1 _15038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [18]),
    .B(_3796__bF$buf3),
    .C(_3798__bF$buf3),
    .Y(_3906_)
);

NAND2X1 _15039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [18]),
    .B(_3800__bF$buf5),
    .Y(_3907_)
);

NAND3X1 _15040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3907_),
    .B(_3906_),
    .C(_3905_),
    .Y(_1_[18])
);

INVX1 _15041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[19]),
    .Y(_3908_)
);

NAND2X1 _15042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf5),
    .B(\datapath.memoryinterface.data_store [3]),
    .Y(_3909_)
);

OAI21X1 _15043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3908_),
    .B(_0__1_bF$buf4),
    .C(_3909_),
    .Y(_3910_)
);

NAND2X1 _15044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf1),
    .B(_3910_),
    .Y(_3911_)
);

NAND3X1 _15045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [19]),
    .B(_3796__bF$buf2),
    .C(_3798__bF$buf2),
    .Y(_3912_)
);

NAND2X1 _15046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [19]),
    .B(_3800__bF$buf4),
    .Y(_3913_)
);

NAND3X1 _15047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3913_),
    .B(_3912_),
    .C(_3911_),
    .Y(_1_[19])
);

INVX1 _15048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[20]),
    .Y(_3914_)
);

NAND2X1 _15049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf3),
    .B(\datapath.memoryinterface.data_store [4]),
    .Y(_3915_)
);

OAI21X1 _15050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3914_),
    .B(_0__1_bF$buf2),
    .C(_3915_),
    .Y(_3916_)
);

NAND2X1 _15051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf0),
    .B(_3916_),
    .Y(_3917_)
);

NAND3X1 _15052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [20]),
    .B(_3796__bF$buf1),
    .C(_3798__bF$buf1),
    .Y(_3918_)
);

NAND2X1 _15053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [20]),
    .B(_3800__bF$buf3),
    .Y(_3919_)
);

NAND3X1 _15054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3919_),
    .B(_3918_),
    .C(_3917_),
    .Y(_1_[20])
);

INVX1 _15055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[21]),
    .Y(_3920_)
);

NAND2X1 _15056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf1),
    .B(\datapath.memoryinterface.data_store [5]),
    .Y(_3921_)
);

OAI21X1 _15057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3920_),
    .B(_0__1_bF$buf0),
    .C(_3921_),
    .Y(_3922_)
);

NAND2X1 _15058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf6),
    .B(_3922_),
    .Y(_3923_)
);

NAND3X1 _15059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [21]),
    .B(_3796__bF$buf0),
    .C(_3798__bF$buf0),
    .Y(_3924_)
);

NAND2X1 _15060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [21]),
    .B(_3800__bF$buf2),
    .Y(_3925_)
);

NAND3X1 _15061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3925_),
    .B(_3924_),
    .C(_3923_),
    .Y(_1_[21])
);

INVX1 _15062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[22]),
    .Y(_3926_)
);

NAND2X1 _15063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf9),
    .B(\datapath.memoryinterface.data_store [6]),
    .Y(_3927_)
);

OAI21X1 _15064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3926_),
    .B(_0__1_bF$buf8),
    .C(_3927_),
    .Y(_3928_)
);

NAND2X1 _15065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf5),
    .B(_3928_),
    .Y(_3929_)
);

NAND3X1 _15066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [22]),
    .B(_3796__bF$buf4),
    .C(_3798__bF$buf4),
    .Y(_3930_)
);

NAND2X1 _15067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [22]),
    .B(_3800__bF$buf1),
    .Y(_3931_)
);

NAND3X1 _15068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3931_),
    .B(_3930_),
    .C(_3929_),
    .Y(_1_[22])
);

INVX1 _15069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[23]),
    .Y(_3932_)
);

NAND2X1 _15070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf7),
    .B(\datapath.memoryinterface.data_store [7]),
    .Y(_3933_)
);

OAI21X1 _15071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3932_),
    .B(_0__1_bF$buf6),
    .C(_3933_),
    .Y(_3934_)
);

NAND2X1 _15072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf4),
    .B(_3934_),
    .Y(_3935_)
);

NAND3X1 _15073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [23]),
    .B(_3796__bF$buf3),
    .C(_3798__bF$buf3),
    .Y(_3936_)
);

NAND2X1 _15074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [23]),
    .B(_3800__bF$buf0),
    .Y(_3937_)
);

NAND3X1 _15075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3937_),
    .B(_3936_),
    .C(_3935_),
    .Y(_1_[23])
);

INVX1 _15076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[24]),
    .Y(_3938_)
);

NAND2X1 _15077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf5),
    .B(\datapath.memoryinterface.data_store [8]),
    .Y(_3939_)
);

OAI21X1 _15078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3938_),
    .B(_0__1_bF$buf4),
    .C(_3939_),
    .Y(_3940_)
);

NAND2X1 _15079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf3),
    .B(_3940_),
    .Y(_3941_)
);

NAND3X1 _15080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [24]),
    .B(_3796__bF$buf2),
    .C(_3798__bF$buf2),
    .Y(_3942_)
);

NAND2X1 _15081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [24]),
    .B(_3800__bF$buf7),
    .Y(_3943_)
);

NAND3X1 _15082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3943_),
    .B(_3942_),
    .C(_3941_),
    .Y(_1_[24])
);

INVX1 _15083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[25]),
    .Y(_3944_)
);

NAND2X1 _15084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf3),
    .B(\datapath.memoryinterface.data_store [9]),
    .Y(_3945_)
);

OAI21X1 _15085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3944_),
    .B(_0__1_bF$buf2),
    .C(_3945_),
    .Y(_3946_)
);

NAND2X1 _15086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf2),
    .B(_3946_),
    .Y(_3947_)
);

NAND3X1 _15087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [25]),
    .B(_3796__bF$buf1),
    .C(_3798__bF$buf1),
    .Y(_3948_)
);

NAND2X1 _15088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [25]),
    .B(_3800__bF$buf6),
    .Y(_3949_)
);

NAND3X1 _15089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3949_),
    .B(_3948_),
    .C(_3947_),
    .Y(_1_[25])
);

INVX1 _15090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[26]),
    .Y(_3950_)
);

NAND2X1 _15091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf1),
    .B(\datapath.memoryinterface.data_store [10]),
    .Y(_3951_)
);

OAI21X1 _15092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3950_),
    .B(_0__1_bF$buf0),
    .C(_3951_),
    .Y(_3952_)
);

NAND2X1 _15093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf1),
    .B(_3952_),
    .Y(_3953_)
);

NAND3X1 _15094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [26]),
    .B(_3796__bF$buf0),
    .C(_3798__bF$buf0),
    .Y(_3954_)
);

NAND2X1 _15095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [26]),
    .B(_3800__bF$buf5),
    .Y(_3955_)
);

NAND3X1 _15096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3955_),
    .B(_3954_),
    .C(_3953_),
    .Y(_1_[26])
);

INVX1 _15097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[27]),
    .Y(_3956_)
);

NAND2X1 _15098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf9),
    .B(\datapath.memoryinterface.data_store [11]),
    .Y(_3957_)
);

OAI21X1 _15099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3956_),
    .B(_0__1_bF$buf8),
    .C(_3957_),
    .Y(_3958_)
);

NAND2X1 _15100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf0),
    .B(_3958_),
    .Y(_3959_)
);

NAND3X1 _15101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [27]),
    .B(_3796__bF$buf4),
    .C(_3798__bF$buf4),
    .Y(_3960_)
);

NAND2X1 _15102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [27]),
    .B(_3800__bF$buf4),
    .Y(_3961_)
);

NAND3X1 _15103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3961_),
    .B(_3960_),
    .C(_3959_),
    .Y(_1_[27])
);

INVX1 _15104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[28]),
    .Y(_3962_)
);

NAND2X1 _15105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf7),
    .B(\datapath.memoryinterface.data_store [12]),
    .Y(_3963_)
);

OAI21X1 _15106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3962_),
    .B(_0__1_bF$buf6),
    .C(_3963_),
    .Y(_3964_)
);

NAND2X1 _15107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf6),
    .B(_3964_),
    .Y(_3965_)
);

NAND3X1 _15108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [28]),
    .B(_3796__bF$buf3),
    .C(_3798__bF$buf3),
    .Y(_3966_)
);

NAND2X1 _15109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [28]),
    .B(_3800__bF$buf3),
    .Y(_3967_)
);

NAND3X1 _15110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3967_),
    .B(_3966_),
    .C(_3965_),
    .Y(_1_[28])
);

INVX1 _15111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[29]),
    .Y(_3968_)
);

NAND2X1 _15112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf5),
    .B(\datapath.memoryinterface.data_store [13]),
    .Y(_3969_)
);

OAI21X1 _15113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3968_),
    .B(_0__1_bF$buf4),
    .C(_3969_),
    .Y(_3970_)
);

NAND2X1 _15114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf5),
    .B(_3970_),
    .Y(_3971_)
);

NAND3X1 _15115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [29]),
    .B(_3796__bF$buf2),
    .C(_3798__bF$buf2),
    .Y(_3972_)
);

NAND2X1 _15116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [29]),
    .B(_3800__bF$buf2),
    .Y(_3973_)
);

NAND3X1 _15117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3973_),
    .B(_3972_),
    .C(_3971_),
    .Y(_1_[29])
);

INVX1 _15118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[30]),
    .Y(_3974_)
);

NAND2X1 _15119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf3),
    .B(\datapath.memoryinterface.data_store [14]),
    .Y(_3975_)
);

OAI21X1 _15120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3974_),
    .B(_0__1_bF$buf2),
    .C(_3975_),
    .Y(_3976_)
);

NAND2X1 _15121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf4),
    .B(_3976_),
    .Y(_3977_)
);

NAND3X1 _15122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [30]),
    .B(_3796__bF$buf1),
    .C(_3798__bF$buf1),
    .Y(_3978_)
);

NAND2X1 _15123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [30]),
    .B(_3800__bF$buf1),
    .Y(_3979_)
);

NAND3X1 _15124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3979_),
    .B(_3978_),
    .C(_3977_),
    .Y(_1_[30])
);

INVX1 _15125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[31]),
    .Y(_3980_)
);

NAND2X1 _15126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf1),
    .B(\datapath.memoryinterface.data_store [15]),
    .Y(_3981_)
);

OAI21X1 _15127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3980_),
    .B(_0__1_bF$buf0),
    .C(_3981_),
    .Y(_3982_)
);

NAND2X1 _15128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf3),
    .B(_3982_),
    .Y(_3983_)
);

NAND3X1 _15129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_store.storebyte [31]),
    .B(_3796__bF$buf0),
    .C(_3798__bF$buf0),
    .Y(_3984_)
);

NAND2X1 _15130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [31]),
    .B(_3800__bF$buf0),
    .Y(_3985_)
);

NAND3X1 _15131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3985_),
    .B(_3984_),
    .C(_3983_),
    .Y(_1_[31])
);

NOR2X1 _15132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf9),
    .B(_0__0_bF$buf3),
    .Y(_3986_)
);

INVX4 _15133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3986_),
    .Y(_3987_)
);

OAI21X1 _15134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf8),
    .B(_0__0_bF$buf2),
    .C(DMEM_DATA_L[0]),
    .Y(_3988_)
);

OAI21X1 _15135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3987_),
    .B(_3803_),
    .C(_3988_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [0])
);

OAI21X1 _15136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf7),
    .B(_0__0_bF$buf1),
    .C(DMEM_DATA_L[1]),
    .Y(_3989_)
);

OAI21X1 _15137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3987_),
    .B(_3809_),
    .C(_3989_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [1])
);

OAI21X1 _15138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf6),
    .B(_0__0_bF$buf0),
    .C(DMEM_DATA_L[2]),
    .Y(_3990_)
);

OAI21X1 _15139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3987_),
    .B(_3815_),
    .C(_3990_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [2])
);

OAI21X1 _15140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf5),
    .B(_0__0_bF$buf4),
    .C(DMEM_DATA_L[3]),
    .Y(_3991_)
);

OAI21X1 _15141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3987_),
    .B(_3821_),
    .C(_3991_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [3])
);

OAI21X1 _15142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf4),
    .B(_0__0_bF$buf3),
    .C(DMEM_DATA_L[4]),
    .Y(_3992_)
);

OAI21X1 _15143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3987_),
    .B(_3827_),
    .C(_3992_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [4])
);

OAI21X1 _15144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf3),
    .B(_0__0_bF$buf2),
    .C(DMEM_DATA_L[5]),
    .Y(_3993_)
);

OAI21X1 _15145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3987_),
    .B(_3833_),
    .C(_3993_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [5])
);

OAI21X1 _15146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf2),
    .B(_0__0_bF$buf1),
    .C(DMEM_DATA_L[6]),
    .Y(_3994_)
);

OAI21X1 _15147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3987_),
    .B(_3839_),
    .C(_3994_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [6])
);

OAI21X1 _15148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf1),
    .B(_0__0_bF$buf0),
    .C(DMEM_DATA_L[7]),
    .Y(_3995_)
);

OAI21X1 _15149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3987_),
    .B(_3845_),
    .C(_3995_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [7])
);

INVX1 _15150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[8]),
    .Y(_3996_)
);

INVX1 _15151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__0_bF$buf4),
    .Y(_3997_)
);

NOR2X1 _15152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf0),
    .B(_3997_),
    .Y(_3998_)
);

MUX2X1 _15153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3803_),
    .B(_3996_),
    .S(_3998_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [8])
);

INVX1 _15154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[9]),
    .Y(_3999_)
);

MUX2X1 _15155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3809_),
    .B(_3999_),
    .S(_3998_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [9])
);

INVX1 _15156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[10]),
    .Y(_4000_)
);

MUX2X1 _15157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3815_),
    .B(_4000_),
    .S(_3998_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [10])
);

INVX1 _15158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[11]),
    .Y(_4001_)
);

MUX2X1 _15159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3821_),
    .B(_4001_),
    .S(_3998_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [11])
);

INVX1 _15160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[12]),
    .Y(_4002_)
);

MUX2X1 _15161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3827_),
    .B(_4002_),
    .S(_3998_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [12])
);

INVX1 _15162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[13]),
    .Y(_4003_)
);

MUX2X1 _15163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3833_),
    .B(_4003_),
    .S(_3998_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [13])
);

INVX1 _15164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[14]),
    .Y(_4004_)
);

MUX2X1 _15165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3839_),
    .B(_4004_),
    .S(_3998_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [14])
);

INVX1 _15166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[15]),
    .Y(_4005_)
);

MUX2X1 _15167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3845_),
    .B(_4005_),
    .S(_3998_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [15])
);

INVX1 _15168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf9),
    .Y(_4006_)
);

NOR2X1 _15169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__0_bF$buf3),
    .B(_4006_),
    .Y(_4007_)
);

OAI22X1 _15170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__0_bF$buf2),
    .B(_3891_),
    .C(_4007_),
    .D(_3890_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [16])
);

OAI22X1 _15171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__0_bF$buf1),
    .B(_3897_),
    .C(_4007_),
    .D(_3896_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [17])
);

OAI22X1 _15172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__0_bF$buf0),
    .B(_3903_),
    .C(_4007_),
    .D(_3902_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [18])
);

OAI22X1 _15173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__0_bF$buf4),
    .B(_3909_),
    .C(_4007_),
    .D(_3908_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [19])
);

OAI22X1 _15174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__0_bF$buf3),
    .B(_3915_),
    .C(_4007_),
    .D(_3914_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [20])
);

OAI22X1 _15175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__0_bF$buf2),
    .B(_3921_),
    .C(_4007_),
    .D(_3920_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [21])
);

OAI22X1 _15176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__0_bF$buf1),
    .B(_3927_),
    .C(_4007_),
    .D(_3926_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [22])
);

OAI22X1 _15177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__0_bF$buf0),
    .B(_3933_),
    .C(_4007_),
    .D(_3932_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [23])
);

NOR2X1 _15178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4006_),
    .B(_3997_),
    .Y(_4008_)
);

NAND2X1 _15179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [0]),
    .B(_4008__bF$buf3),
    .Y(_4009_)
);

OAI21X1 _15180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3938_),
    .B(_4008__bF$buf2),
    .C(_4009_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [24])
);

NAND2X1 _15181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [1]),
    .B(_4008__bF$buf1),
    .Y(_4010_)
);

OAI21X1 _15182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3944_),
    .B(_4008__bF$buf0),
    .C(_4010_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [25])
);

NAND2X1 _15183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [2]),
    .B(_4008__bF$buf3),
    .Y(_4011_)
);

OAI21X1 _15184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3950_),
    .B(_4008__bF$buf2),
    .C(_4011_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [26])
);

NAND2X1 _15185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [3]),
    .B(_4008__bF$buf1),
    .Y(_4012_)
);

OAI21X1 _15186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3956_),
    .B(_4008__bF$buf0),
    .C(_4012_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [27])
);

NAND2X1 _15187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [4]),
    .B(_4008__bF$buf3),
    .Y(_4013_)
);

OAI21X1 _15188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3962_),
    .B(_4008__bF$buf2),
    .C(_4013_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [28])
);

NAND2X1 _15189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [5]),
    .B(_4008__bF$buf1),
    .Y(_4014_)
);

OAI21X1 _15190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3968_),
    .B(_4008__bF$buf0),
    .C(_4014_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [29])
);

NAND2X1 _15191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [6]),
    .B(_4008__bF$buf3),
    .Y(_4015_)
);

OAI21X1 _15192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3974_),
    .B(_4008__bF$buf2),
    .C(_4015_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [30])
);

NAND2X1 _15193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.data_store [7]),
    .B(_4008__bF$buf1),
    .Y(_4016_)
);

OAI21X1 _15194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3980_),
    .B(_4008__bF$buf0),
    .C(_4016_),
    .Y(\datapath.memoryinterface.byte_size_store.storebyte [31])
);

INVX1 _15195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_load.byteval [0]),
    .Y(_4017_)
);

INVX1 _15196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[0]),
    .Y(_4018_)
);

NAND2X1 _15197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf8),
    .B(DMEM_DATA_L[16]),
    .Y(_4019_)
);

OAI21X1 _15198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4018_),
    .B(_0__1_bF$buf7),
    .C(_4019_),
    .Y(_4020_)
);

AOI22X1 _15199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[0]),
    .B(_3800__bF$buf7),
    .C(_4020_),
    .D(_3802__bF$buf2),
    .Y(_4021_)
);

OAI21X1 _15200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4017_),
    .B(_3850_),
    .C(_4021_),
    .Y(\datapath.memdataload [0])
);

INVX1 _15201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_load.byteval [1]),
    .Y(_4022_)
);

INVX1 _15202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[1]),
    .Y(_4023_)
);

NAND2X1 _15203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf6),
    .B(DMEM_DATA_L[17]),
    .Y(_4024_)
);

OAI21X1 _15204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4023_),
    .B(_0__1_bF$buf5),
    .C(_4024_),
    .Y(_4025_)
);

AOI22X1 _15205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[1]),
    .B(_3800__bF$buf6),
    .C(_4025_),
    .D(_3802__bF$buf1),
    .Y(_4026_)
);

OAI21X1 _15206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4022_),
    .B(_3850_),
    .C(_4026_),
    .Y(\datapath.memdataload [1])
);

INVX1 _15207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_load.byteval [2]),
    .Y(_4027_)
);

INVX1 _15208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[2]),
    .Y(_4028_)
);

NAND2X1 _15209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf4),
    .B(DMEM_DATA_L[18]),
    .Y(_4029_)
);

OAI21X1 _15210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4028_),
    .B(_0__1_bF$buf3),
    .C(_4029_),
    .Y(_4030_)
);

AOI22X1 _15211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[2]),
    .B(_3800__bF$buf5),
    .C(_4030_),
    .D(_3802__bF$buf0),
    .Y(_4031_)
);

OAI21X1 _15212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4027_),
    .B(_3850_),
    .C(_4031_),
    .Y(\datapath.memdataload [2])
);

INVX1 _15213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_load.byteval [3]),
    .Y(_4032_)
);

INVX1 _15214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[3]),
    .Y(_4033_)
);

NAND2X1 _15215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf2),
    .B(DMEM_DATA_L[19]),
    .Y(_4034_)
);

OAI21X1 _15216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4033_),
    .B(_0__1_bF$buf1),
    .C(_4034_),
    .Y(_4035_)
);

AOI22X1 _15217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[3]),
    .B(_3800__bF$buf4),
    .C(_4035_),
    .D(_3802__bF$buf6),
    .Y(_4036_)
);

OAI21X1 _15218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4032_),
    .B(_3850_),
    .C(_4036_),
    .Y(\datapath.memdataload [3])
);

INVX1 _15219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_load.byteval [4]),
    .Y(_4037_)
);

INVX1 _15220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[4]),
    .Y(_4038_)
);

NAND2X1 _15221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf0),
    .B(DMEM_DATA_L[20]),
    .Y(_4039_)
);

OAI21X1 _15222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4038_),
    .B(_0__1_bF$buf9),
    .C(_4039_),
    .Y(_4040_)
);

AOI22X1 _15223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[4]),
    .B(_3800__bF$buf3),
    .C(_4040_),
    .D(_3802__bF$buf5),
    .Y(_4041_)
);

OAI21X1 _15224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4037_),
    .B(_3850_),
    .C(_4041_),
    .Y(\datapath.memdataload [4])
);

INVX1 _15225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_load.byteval [5]),
    .Y(_4042_)
);

INVX1 _15226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[5]),
    .Y(_4043_)
);

NAND2X1 _15227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf8),
    .B(DMEM_DATA_L[21]),
    .Y(_4044_)
);

OAI21X1 _15228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4043_),
    .B(_0__1_bF$buf7),
    .C(_4044_),
    .Y(_4045_)
);

AOI22X1 _15229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[5]),
    .B(_3800__bF$buf2),
    .C(_4045_),
    .D(_3802__bF$buf4),
    .Y(_4046_)
);

OAI21X1 _15230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4042_),
    .B(_3850_),
    .C(_4046_),
    .Y(\datapath.memdataload [5])
);

INVX1 _15231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_load.byteval [6]),
    .Y(_4047_)
);

INVX1 _15232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[6]),
    .Y(_4048_)
);

NAND2X1 _15233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf6),
    .B(DMEM_DATA_L[22]),
    .Y(_4049_)
);

OAI21X1 _15234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4048_),
    .B(_0__1_bF$buf5),
    .C(_4049_),
    .Y(_4050_)
);

AOI22X1 _15235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[6]),
    .B(_3800__bF$buf1),
    .C(_4050_),
    .D(_3802__bF$buf3),
    .Y(_4051_)
);

OAI21X1 _15236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4047_),
    .B(_3850_),
    .C(_4051_),
    .Y(\datapath.memdataload [6])
);

NAND3X1 _15237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_load.byteval [7]),
    .B(_3796__bF$buf4),
    .C(_3798__bF$buf4),
    .Y(_4052_)
);

NAND2X1 _15238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[7]),
    .B(_3800__bF$buf0),
    .Y(_4053_)
);

INVX1 _15239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[7]),
    .Y(_4054_)
);

NAND2X1 _15240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf4),
    .B(DMEM_DATA_L[23]),
    .Y(_4055_)
);

OAI21X1 _15241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4054_),
    .B(_0__1_bF$buf3),
    .C(_4055_),
    .Y(_4056_)
);

NAND2X1 _15242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf2),
    .B(_4056_),
    .Y(_4057_)
);

NAND3X1 _15243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4053_),
    .B(_4052_),
    .C(_4057_),
    .Y(\datapath.memdataload [7])
);

INVX1 _15244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memoryinterface.byte_size_load.byteval [7]),
    .Y(_4058_)
);

NOR2X1 _15245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [14]),
    .B(_4058_),
    .Y(_4059_)
);

NAND3X1 _15246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3796__bF$buf3),
    .B(_3798__bF$buf3),
    .C(_4059_),
    .Y(_4060_)
);

NAND2X1 _15247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[8]),
    .B(_3800__bF$buf7),
    .Y(_4061_)
);

NAND2X1 _15248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf2),
    .B(DMEM_DATA_L[24]),
    .Y(_4062_)
);

OAI21X1 _15249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3996_),
    .B(_0__1_bF$buf1),
    .C(_4062_),
    .Y(_4063_)
);

NAND2X1 _15250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf1),
    .B(_4063_),
    .Y(_4064_)
);

NAND3X1 _15251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4061_),
    .B(_4064_),
    .C(_4060__bF$buf3),
    .Y(\datapath.memdataload [8])
);

NAND2X1 _15252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[9]),
    .B(_3800__bF$buf6),
    .Y(_4065_)
);

NAND2X1 _15253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf0),
    .B(DMEM_DATA_L[25]),
    .Y(_4066_)
);

OAI21X1 _15254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3999_),
    .B(_0__1_bF$buf9),
    .C(_4066_),
    .Y(_4067_)
);

NAND2X1 _15255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf0),
    .B(_4067_),
    .Y(_4068_)
);

NAND3X1 _15256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4065_),
    .B(_4068_),
    .C(_4060__bF$buf2),
    .Y(\datapath.memdataload [9])
);

NAND2X1 _15257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[10]),
    .B(_3800__bF$buf5),
    .Y(_4069_)
);

NAND2X1 _15258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf8),
    .B(DMEM_DATA_L[26]),
    .Y(_4070_)
);

OAI21X1 _15259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4000_),
    .B(_0__1_bF$buf7),
    .C(_4070_),
    .Y(_4071_)
);

NAND2X1 _15260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf6),
    .B(_4071_),
    .Y(_4072_)
);

NAND3X1 _15261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4069_),
    .B(_4072_),
    .C(_4060__bF$buf1),
    .Y(\datapath.memdataload [10])
);

NAND2X1 _15262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[11]),
    .B(_3800__bF$buf4),
    .Y(_4073_)
);

NAND2X1 _15263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf6),
    .B(DMEM_DATA_L[27]),
    .Y(_4074_)
);

OAI21X1 _15264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4001_),
    .B(_0__1_bF$buf5),
    .C(_4074_),
    .Y(_4075_)
);

NAND2X1 _15265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf5),
    .B(_4075_),
    .Y(_4076_)
);

NAND3X1 _15266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4073_),
    .B(_4076_),
    .C(_4060__bF$buf0),
    .Y(\datapath.memdataload [11])
);

NAND2X1 _15267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[12]),
    .B(_3800__bF$buf3),
    .Y(_4077_)
);

NAND2X1 _15268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf4),
    .B(DMEM_DATA_L[28]),
    .Y(_4078_)
);

OAI21X1 _15269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4002_),
    .B(_0__1_bF$buf3),
    .C(_4078_),
    .Y(_4079_)
);

NAND2X1 _15270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf4),
    .B(_4079_),
    .Y(_4080_)
);

NAND3X1 _15271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4077_),
    .B(_4080_),
    .C(_4060__bF$buf3),
    .Y(\datapath.memdataload [12])
);

NAND2X1 _15272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[13]),
    .B(_3800__bF$buf2),
    .Y(_4081_)
);

NAND2X1 _15273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf2),
    .B(DMEM_DATA_L[29]),
    .Y(_4082_)
);

OAI21X1 _15274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4003_),
    .B(_0__1_bF$buf1),
    .C(_4082_),
    .Y(_4083_)
);

NAND2X1 _15275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf3),
    .B(_4083_),
    .Y(_4084_)
);

NAND3X1 _15276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4081_),
    .B(_4084_),
    .C(_4060__bF$buf2),
    .Y(\datapath.memdataload [13])
);

NAND2X1 _15277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[14]),
    .B(_3800__bF$buf1),
    .Y(_4085_)
);

NAND2X1 _15278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf0),
    .B(DMEM_DATA_L[30]),
    .Y(_4086_)
);

OAI21X1 _15279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4004_),
    .B(_0__1_bF$buf9),
    .C(_4086_),
    .Y(_4087_)
);

NAND2X1 _15280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf2),
    .B(_4087_),
    .Y(_4088_)
);

NAND3X1 _15281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4085_),
    .B(_4088_),
    .C(_4060__bF$buf1),
    .Y(\datapath.memdataload [14])
);

NAND2X1 _15282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf8),
    .B(DMEM_DATA_L[31]),
    .Y(_4089_)
);

OAI21X1 _15283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4005_),
    .B(_0__1_bF$buf7),
    .C(_4089_),
    .Y(_4090_)
);

NAND2X1 _15284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802__bF$buf1),
    .B(_4090_),
    .Y(_4091_)
);

NAND2X1 _15285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[15]),
    .B(_3800__bF$buf0),
    .Y(_4092_)
);

NAND3X1 _15286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4092_),
    .B(_4091_),
    .C(_4060__bF$buf0),
    .Y(\datapath.memdataload [15])
);

NAND2X1 _15287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[16]),
    .B(_3800__bF$buf7),
    .Y(_4093_)
);

INVX1 _15288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [14]),
    .Y(_4094_)
);

NAND3X1 _15289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4094_),
    .B(_3802__bF$buf0),
    .C(_4090_),
    .Y(_4095_)
);

NAND3X1 _15290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060__bF$buf3),
    .B(_4093_),
    .C(_4095_),
    .Y(\datapath.memdataload [16])
);

NAND2X1 _15291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[17]),
    .B(_3800__bF$buf6),
    .Y(_4096_)
);

NAND3X1 _15292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060__bF$buf2),
    .B(_4096_),
    .C(_4095_),
    .Y(\datapath.memdataload [17])
);

NAND2X1 _15293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[18]),
    .B(_3800__bF$buf5),
    .Y(_4097_)
);

NAND3X1 _15294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060__bF$buf1),
    .B(_4097_),
    .C(_4095_),
    .Y(\datapath.memdataload [18])
);

NAND2X1 _15295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[19]),
    .B(_3800__bF$buf4),
    .Y(_4098_)
);

NAND3X1 _15296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060__bF$buf0),
    .B(_4098_),
    .C(_4095_),
    .Y(\datapath.memdataload [19])
);

NAND2X1 _15297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[20]),
    .B(_3800__bF$buf3),
    .Y(_4099_)
);

NAND3X1 _15298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060__bF$buf3),
    .B(_4099_),
    .C(_4095_),
    .Y(\datapath.memdataload [20])
);

NAND2X1 _15299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[21]),
    .B(_3800__bF$buf2),
    .Y(_4100_)
);

NAND3X1 _15300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060__bF$buf2),
    .B(_4100_),
    .C(_4095_),
    .Y(\datapath.memdataload [21])
);

NAND2X1 _15301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[22]),
    .B(_3800__bF$buf1),
    .Y(_4101_)
);

NAND3X1 _15302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060__bF$buf1),
    .B(_4101_),
    .C(_4095_),
    .Y(\datapath.memdataload [22])
);

NAND2X1 _15303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[23]),
    .B(_3800__bF$buf0),
    .Y(_4102_)
);

NAND3X1 _15304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060__bF$buf0),
    .B(_4102_),
    .C(_4095_),
    .Y(\datapath.memdataload [23])
);

NAND2X1 _15305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[24]),
    .B(_3800__bF$buf7),
    .Y(_4103_)
);

NAND3X1 _15306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060__bF$buf3),
    .B(_4103_),
    .C(_4095_),
    .Y(\datapath.memdataload [24])
);

NAND2X1 _15307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[25]),
    .B(_3800__bF$buf6),
    .Y(_4104_)
);

NAND3X1 _15308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060__bF$buf2),
    .B(_4104_),
    .C(_4095_),
    .Y(\datapath.memdataload [25])
);

NAND2X1 _15309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[26]),
    .B(_3800__bF$buf5),
    .Y(_4105_)
);

NAND3X1 _15310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060__bF$buf1),
    .B(_4105_),
    .C(_4095_),
    .Y(\datapath.memdataload [26])
);

NAND2X1 _15311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[27]),
    .B(_3800__bF$buf4),
    .Y(_4106_)
);

NAND3X1 _15312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060__bF$buf0),
    .B(_4106_),
    .C(_4095_),
    .Y(\datapath.memdataload [27])
);

NAND2X1 _15313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[28]),
    .B(_3800__bF$buf3),
    .Y(_4107_)
);

NAND3X1 _15314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060__bF$buf3),
    .B(_4107_),
    .C(_4095_),
    .Y(\datapath.memdataload [28])
);

NAND2X1 _15315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[29]),
    .B(_3800__bF$buf2),
    .Y(_4108_)
);

NAND3X1 _15316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060__bF$buf2),
    .B(_4108_),
    .C(_4095_),
    .Y(\datapath.memdataload [29])
);

NAND2X1 _15317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[30]),
    .B(_3800__bF$buf1),
    .Y(_4109_)
);

NAND3X1 _15318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060__bF$buf1),
    .B(_4109_),
    .C(_4095_),
    .Y(\datapath.memdataload [30])
);

NAND2X1 _15319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[31]),
    .B(_3800__bF$buf0),
    .Y(_4110_)
);

NAND3X1 _15320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060__bF$buf0),
    .B(_4110_),
    .C(_4095_),
    .Y(\datapath.memdataload [31])
);

AOI22X1 _15321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4007_),
    .B(DMEM_DATA_L[16]),
    .C(DMEM_DATA_L[24]),
    .D(_4008__bF$buf3),
    .Y(_4111_)
);

AOI22X1 _15322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[0]),
    .B(_3986_),
    .C(_3998_),
    .D(DMEM_DATA_L[8]),
    .Y(_4112_)
);

NAND2X1 _15323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4112_),
    .B(_4111_),
    .Y(\datapath.memoryinterface.byte_size_load.byteval [0])
);

AOI22X1 _15324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4007_),
    .B(DMEM_DATA_L[17]),
    .C(DMEM_DATA_L[25]),
    .D(_4008__bF$buf2),
    .Y(_4113_)
);

AOI22X1 _15325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[1]),
    .B(_3986_),
    .C(_3998_),
    .D(DMEM_DATA_L[9]),
    .Y(_4114_)
);

NAND2X1 _15326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4114_),
    .B(_4113_),
    .Y(\datapath.memoryinterface.byte_size_load.byteval [1])
);

AOI22X1 _15327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4007_),
    .B(DMEM_DATA_L[18]),
    .C(DMEM_DATA_L[26]),
    .D(_4008__bF$buf1),
    .Y(_4115_)
);

AOI22X1 _15328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[2]),
    .B(_3986_),
    .C(_3998_),
    .D(DMEM_DATA_L[10]),
    .Y(_4116_)
);

NAND2X1 _15329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116_),
    .B(_4115_),
    .Y(\datapath.memoryinterface.byte_size_load.byteval [2])
);

AOI22X1 _15330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4007_),
    .B(DMEM_DATA_L[19]),
    .C(DMEM_DATA_L[27]),
    .D(_4008__bF$buf0),
    .Y(_4117_)
);

AOI22X1 _15331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[3]),
    .B(_3986_),
    .C(_3998_),
    .D(DMEM_DATA_L[11]),
    .Y(_4118_)
);

NAND2X1 _15332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4118_),
    .B(_4117_),
    .Y(\datapath.memoryinterface.byte_size_load.byteval [3])
);

AOI22X1 _15333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4007_),
    .B(DMEM_DATA_L[20]),
    .C(DMEM_DATA_L[28]),
    .D(_4008__bF$buf3),
    .Y(_4119_)
);

AOI22X1 _15334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[4]),
    .B(_3986_),
    .C(_3998_),
    .D(DMEM_DATA_L[12]),
    .Y(_4120_)
);

NAND2X1 _15335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4120_),
    .B(_4119_),
    .Y(\datapath.memoryinterface.byte_size_load.byteval [4])
);

AOI22X1 _15336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4007_),
    .B(DMEM_DATA_L[21]),
    .C(DMEM_DATA_L[29]),
    .D(_4008__bF$buf2),
    .Y(_4121_)
);

AOI22X1 _15337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[5]),
    .B(_3986_),
    .C(_3998_),
    .D(DMEM_DATA_L[13]),
    .Y(_4122_)
);

NAND2X1 _15338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4122_),
    .B(_4121_),
    .Y(\datapath.memoryinterface.byte_size_load.byteval [5])
);

AOI22X1 _15339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4007_),
    .B(DMEM_DATA_L[22]),
    .C(DMEM_DATA_L[30]),
    .D(_4008__bF$buf1),
    .Y(_4123_)
);

AOI22X1 _15340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[6]),
    .B(_3986_),
    .C(_3998_),
    .D(DMEM_DATA_L[14]),
    .Y(_4124_)
);

NAND2X1 _15341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4124_),
    .B(_4123_),
    .Y(\datapath.memoryinterface.byte_size_load.byteval [6])
);

AOI22X1 _15342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[7]),
    .B(_3986_),
    .C(_4007_),
    .D(DMEM_DATA_L[23]),
    .Y(_4125_)
);

NAND2X1 _15343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[15]),
    .B(_3998_),
    .Y(_4126_)
);

NAND2X1 _15344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(DMEM_DATA_L[31]),
    .B(_4008__bF$buf0),
    .Y(_4127_)
);

NAND3X1 _15345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4126_),
    .B(_4127_),
    .C(_4125_),
    .Y(\datapath.memoryinterface.byte_size_load.byteval [7])
);

INVX1 _15346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc_mux [0]),
    .Y(_4128_)
);

NAND2X1 _15347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [0]),
    .B(\datapath.pcstall_bF$buf7 ),
    .Y(_4129_)
);

OAI21X1 _15348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4128_),
    .B(\datapath.pcstall_bF$buf6 ),
    .C(_4129_),
    .Y(\datapath.programcounter._1_ [0])
);

INVX1 _15349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc_mux [1]),
    .Y(_4130_)
);

NAND2X1 _15350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf5 ),
    .B(\datapath.programcounter.pc [1]),
    .Y(_4131_)
);

OAI21X1 _15351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4130_),
    .B(\datapath.pcstall_bF$buf4 ),
    .C(_4131_),
    .Y(\datapath.programcounter._1_ [1])
);

INVX2 _15352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [2]),
    .Y(\datapath.nextpc [2])
);

NOR2X1 _15353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf3 ),
    .B(\datapath.programcounter.pc_mux [2]),
    .Y(_4132_)
);

AOI21X1 _15354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf2 ),
    .B(\datapath.nextpc [2]),
    .C(_4132_),
    .Y(\datapath.programcounter._1_ [2])
);

INVX1 _15355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [3]),
    .Y(_4133_)
);

NOR2X1 _15356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf1 ),
    .B(\datapath.programcounter.pc_mux [3]),
    .Y(_4134_)
);

AOI21X1 _15357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf0 ),
    .B(_4133_),
    .C(_4134_),
    .Y(\datapath.programcounter._1_ [3])
);

INVX1 _15358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [4]),
    .Y(_4135_)
);

NOR2X1 _15359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf7 ),
    .B(\datapath.programcounter.pc_mux [4]),
    .Y(_4136_)
);

AOI21X1 _15360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf6 ),
    .B(_4135_),
    .C(_4136_),
    .Y(\datapath.programcounter._1_ [4])
);

INVX1 _15361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [5]),
    .Y(_4137_)
);

NOR2X1 _15362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf5 ),
    .B(\datapath.programcounter.pc_mux [5]),
    .Y(_4138_)
);

AOI21X1 _15363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf4 ),
    .B(_4137_),
    .C(_4138_),
    .Y(\datapath.programcounter._1_ [5])
);

INVX1 _15364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [6]),
    .Y(_4139_)
);

NOR2X1 _15365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf3 ),
    .B(\datapath.programcounter.pc_mux [6]),
    .Y(_4140_)
);

AOI21X1 _15366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf2 ),
    .B(_4139_),
    .C(_4140_),
    .Y(\datapath.programcounter._1_ [6])
);

INVX1 _15367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [7]),
    .Y(_4141_)
);

NOR2X1 _15368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf1 ),
    .B(\datapath.programcounter.pc_mux [7]),
    .Y(_4142_)
);

AOI21X1 _15369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf0 ),
    .B(_4141_),
    .C(_4142_),
    .Y(\datapath.programcounter._1_ [7])
);

INVX2 _15370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [8]),
    .Y(_4143_)
);

NOR2X1 _15371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf7 ),
    .B(\datapath.programcounter.pc_mux [8]),
    .Y(_4144_)
);

AOI21X1 _15372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf6 ),
    .B(_4143_),
    .C(_4144_),
    .Y(\datapath.programcounter._1_ [8])
);

INVX1 _15373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc_mux [9]),
    .Y(_4145_)
);

NAND2X1 _15374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf5 ),
    .B(\datapath.programcounter.pc [9]),
    .Y(_4146_)
);

OAI21X1 _15375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4145_),
    .B(\datapath.pcstall_bF$buf4 ),
    .C(_4146_),
    .Y(\datapath.programcounter._1_ [9])
);

INVX1 _15376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [10]),
    .Y(_4147_)
);

NOR2X1 _15377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf3 ),
    .B(\datapath.programcounter.pc_mux [10]),
    .Y(_4148_)
);

AOI21X1 _15378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf2 ),
    .B(_4147_),
    .C(_4148_),
    .Y(\datapath.programcounter._1_ [10])
);

INVX1 _15379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc_mux [11]),
    .Y(_4149_)
);

NAND2X1 _15380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf1 ),
    .B(\datapath.programcounter.pc [11]),
    .Y(_4150_)
);

OAI21X1 _15381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4149_),
    .B(\datapath.pcstall_bF$buf0 ),
    .C(_4150_),
    .Y(\datapath.programcounter._1_ [11])
);

INVX1 _15382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [12]),
    .Y(_4151_)
);

NOR2X1 _15383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf7 ),
    .B(\datapath.programcounter.pc_mux [12]),
    .Y(_4152_)
);

AOI21X1 _15384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf6 ),
    .B(_4151_),
    .C(_4152_),
    .Y(\datapath.programcounter._1_ [12])
);

INVX2 _15385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [13]),
    .Y(_4153_)
);

NOR2X1 _15386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf5 ),
    .B(\datapath.programcounter.pc_mux [13]),
    .Y(_4154_)
);

AOI21X1 _15387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf4 ),
    .B(_4153_),
    .C(_4154_),
    .Y(\datapath.programcounter._1_ [13])
);

INVX1 _15388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [14]),
    .Y(_4155_)
);

NOR2X1 _15389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf3 ),
    .B(\datapath.programcounter.pc_mux [14]),
    .Y(_4156_)
);

AOI21X1 _15390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf2 ),
    .B(_4155_),
    .C(_4156_),
    .Y(\datapath.programcounter._1_ [14])
);

INVX1 _15391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [15]),
    .Y(_4157_)
);

NOR2X1 _15392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf1 ),
    .B(\datapath.programcounter.pc_mux [15]),
    .Y(_4158_)
);

AOI21X1 _15393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf0 ),
    .B(_4157_),
    .C(_4158_),
    .Y(\datapath.programcounter._1_ [15])
);

INVX1 _15394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [16]),
    .Y(_4159_)
);

NOR2X1 _15395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf7 ),
    .B(\datapath.programcounter.pc_mux [16]),
    .Y(_4160_)
);

AOI21X1 _15396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf6 ),
    .B(_4159_),
    .C(_4160_),
    .Y(\datapath.programcounter._1_ [16])
);

INVX2 _15397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [17]),
    .Y(_4161_)
);

NOR2X1 _15398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf5 ),
    .B(\datapath.programcounter.pc_mux [17]),
    .Y(_4162_)
);

AOI21X1 _15399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf4 ),
    .B(_4161_),
    .C(_4162_),
    .Y(\datapath.programcounter._1_ [17])
);

INVX2 _15400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [18]),
    .Y(_4163_)
);

NOR2X1 _15401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf3 ),
    .B(\datapath.programcounter.pc_mux [18]),
    .Y(_4164_)
);

AOI21X1 _15402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf2 ),
    .B(_4163_),
    .C(_4164_),
    .Y(\datapath.programcounter._1_ [18])
);

INVX1 _15403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [19]),
    .Y(_4165_)
);

NOR2X1 _15404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf1 ),
    .B(\datapath.programcounter.pc_mux [19]),
    .Y(_4166_)
);

AOI21X1 _15405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf0 ),
    .B(_4165_),
    .C(_4166_),
    .Y(\datapath.programcounter._1_ [19])
);

INVX1 _15406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [20]),
    .Y(_4167_)
);

NOR2X1 _15407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf7 ),
    .B(\datapath.programcounter.pc_mux [20]),
    .Y(_4168_)
);

AOI21X1 _15408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf6 ),
    .B(_4167_),
    .C(_4168_),
    .Y(\datapath.programcounter._1_ [20])
);

INVX1 _15409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [21]),
    .Y(_4169_)
);

NOR2X1 _15410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf5 ),
    .B(\datapath.programcounter.pc_mux [21]),
    .Y(_4170_)
);

AOI21X1 _15411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf4 ),
    .B(_4169_),
    .C(_4170_),
    .Y(\datapath.programcounter._1_ [21])
);

INVX2 _15412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [22]),
    .Y(_4171_)
);

NOR2X1 _15413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf3 ),
    .B(\datapath.programcounter.pc_mux [22]),
    .Y(_4172_)
);

AOI21X1 _15414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf2 ),
    .B(_4171_),
    .C(_4172_),
    .Y(\datapath.programcounter._1_ [22])
);

INVX1 _15415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc_mux [23]),
    .Y(_4173_)
);

NAND2X1 _15416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf1 ),
    .B(\datapath.programcounter.pc [23]),
    .Y(_4174_)
);

OAI21X1 _15417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4173_),
    .B(\datapath.pcstall_bF$buf0 ),
    .C(_4174_),
    .Y(\datapath.programcounter._1_ [23])
);

INVX2 _15418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [24]),
    .Y(_4175_)
);

NOR2X1 _15419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf7 ),
    .B(\datapath.programcounter.pc_mux [24]),
    .Y(_4176_)
);

AOI21X1 _15420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf6 ),
    .B(_4175_),
    .C(_4176_),
    .Y(\datapath.programcounter._1_ [24])
);

INVX2 _15421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [25]),
    .Y(_4177_)
);

NOR2X1 _15422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf5 ),
    .B(\datapath.programcounter.pc_mux [25]),
    .Y(_4178_)
);

AOI21X1 _15423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf4 ),
    .B(_4177_),
    .C(_4178_),
    .Y(\datapath.programcounter._1_ [25])
);

INVX2 _15424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [26]),
    .Y(_4179_)
);

NOR2X1 _15425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf3 ),
    .B(\datapath.programcounter.pc_mux [26]),
    .Y(_4180_)
);

AOI21X1 _15426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf2 ),
    .B(_4179_),
    .C(_4180_),
    .Y(\datapath.programcounter._1_ [26])
);

INVX1 _15427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [27]),
    .Y(_4181_)
);

NOR2X1 _15428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf1 ),
    .B(\datapath.programcounter.pc_mux [27]),
    .Y(_4182_)
);

AOI21X1 _15429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf0 ),
    .B(_4181_),
    .C(_4182_),
    .Y(\datapath.programcounter._1_ [27])
);

INVX2 _15430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [28]),
    .Y(_4183_)
);

NOR2X1 _15431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf7 ),
    .B(\datapath.programcounter.pc_mux [28]),
    .Y(_4184_)
);

AOI21X1 _15432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf6 ),
    .B(_4183_),
    .C(_4184_),
    .Y(\datapath.programcounter._1_ [28])
);

INVX1 _15433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [29]),
    .Y(_4185_)
);

NOR2X1 _15434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf5 ),
    .B(\datapath.programcounter.pc_mux [29]),
    .Y(_4186_)
);

AOI21X1 _15435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf4 ),
    .B(_4185_),
    .C(_4186_),
    .Y(\datapath.programcounter._1_ [29])
);

INVX2 _15436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [30]),
    .Y(_4187_)
);

NOR2X1 _15437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf3 ),
    .B(\datapath.programcounter.pc_mux [30]),
    .Y(_4188_)
);

AOI21X1 _15438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf2 ),
    .B(_4187_),
    .C(_4188_),
    .Y(\datapath.programcounter._1_ [30])
);

INVX1 _15439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [31]),
    .Y(_4189_)
);

NOR2X1 _15440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf1 ),
    .B(\datapath.programcounter.pc_mux [31]),
    .Y(_4190_)
);

AOI21X1 _15441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.pcstall_bF$buf0 ),
    .B(_4189_),
    .C(_4190_),
    .Y(\datapath.programcounter._1_ [31])
);

INVX1 _15442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath._62_ ),
    .Y(_4191_)
);

NOR2X1 _15443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath._60_ ),
    .B(_4191_),
    .Y(_4192_)
);

NOR2X1 _15444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath._60_ ),
    .B(\datapath._62_ ),
    .Y(_4193_)
);

AOI22X1 _15445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [0]),
    .B(_4193__bF$buf4),
    .C(_4192__bF$buf4),
    .D(gnd),
    .Y(_4194_)
);

INVX1 _15446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath._60_ ),
    .Y(_4195_)
);

NOR2X1 _15447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath._62_ ),
    .B(_4195_),
    .Y(_4196_)
);

NAND2X1 _15448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [0]),
    .B(_4196__bF$buf4),
    .Y(_4197_)
);

NOR2X1 _15449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4195_),
    .B(_4191_),
    .Y(_4198_)
);

NAND2X1 _15450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_4198__bF$buf4),
    .Y(_4199_)
);

NAND3X1 _15451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4197_),
    .B(_4199_),
    .C(_4194_),
    .Y(\datapath.programcounter.pc_mux [0])
);

AOI22X1 _15452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [1]),
    .B(_4193__bF$buf3),
    .C(_4192__bF$buf3),
    .D(_0__1_bF$buf6),
    .Y(_4200_)
);

NAND2X1 _15453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [1]),
    .B(_4196__bF$buf3),
    .Y(_4201_)
);

NAND2X1 _15454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .B(_4198__bF$buf3),
    .Y(_4202_)
);

NAND3X1 _15455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4201_),
    .B(_4202_),
    .C(_4200_),
    .Y(\datapath.programcounter.pc_mux [1])
);

AOI22X1 _15456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [2]),
    .B(_4193__bF$buf2),
    .C(_4192__bF$buf2),
    .D(_0_[2]),
    .Y(_4203_)
);

AOI22X1 _15457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4196__bF$buf2),
    .B(\datapath.programcounter.jumps [2]),
    .C(\datapath.csr.csr_pcaddr [2]),
    .D(_4198__bF$buf2),
    .Y(_4204_)
);

NAND2X1 _15458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4203_),
    .B(_4204_),
    .Y(\datapath.programcounter.pc_mux [2])
);

NOR2X1 _15459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.nextpc [2]),
    .B(_4133_),
    .Y(_4205_)
);

NOR2X1 _15460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [2]),
    .B(\datapath.programcounter.pc [3]),
    .Y(_4206_)
);

NOR2X1 _15461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4206_),
    .B(_4205_),
    .Y(\datapath.nextpc [3])
);

NAND2X1 _15462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf1),
    .B(\datapath.nextpc [3]),
    .Y(_4207_)
);

NAND2X1 _15463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [3]),
    .B(_4196__bF$buf1),
    .Y(_4208_)
);

AOI22X1 _15464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf1),
    .B(_0_[3]),
    .C(\datapath.csr.csr_pcaddr [3]),
    .D(_4198__bF$buf1),
    .Y(_4209_)
);

NAND3X1 _15465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4208_),
    .B(_4209_),
    .C(_4207_),
    .Y(\datapath.programcounter.pc_mux [3])
);

NAND3X1 _15466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [2]),
    .B(\datapath.programcounter.pc [3]),
    .C(\datapath.programcounter.pc [4]),
    .Y(_4210_)
);

INVX2 _15467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4210_),
    .Y(_4211_)
);

NOR2X1 _15468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [4]),
    .B(_4205_),
    .Y(_4212_)
);

NOR2X1 _15469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4211_),
    .B(_4212_),
    .Y(\datapath.nextpc [4])
);

NAND2X1 _15470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf0),
    .B(\datapath.nextpc [4]),
    .Y(_4213_)
);

NAND2X1 _15471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [4]),
    .B(_4196__bF$buf0),
    .Y(_4214_)
);

AOI22X1 _15472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf0),
    .B(_0_[4]),
    .C(\datapath.csr.csr_pcaddr [4]),
    .D(_4198__bF$buf0),
    .Y(_4215_)
);

NAND3X1 _15473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4214_),
    .B(_4215_),
    .C(_4213_),
    .Y(\datapath.programcounter.pc_mux [4])
);

XNOR2X1 _15474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4210_),
    .B(\datapath.programcounter.pc [5]),
    .Y(\datapath.nextpc [5])
);

NAND2X1 _15475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf4),
    .B(\datapath.nextpc [5]),
    .Y(_4216_)
);

NAND2X1 _15476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [5]),
    .B(_4196__bF$buf4),
    .Y(_4217_)
);

AOI22X1 _15477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf4),
    .B(_0_[5]),
    .C(\datapath.csr.csr_pcaddr [5]),
    .D(_4198__bF$buf4),
    .Y(_4218_)
);

NAND3X1 _15478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4217_),
    .B(_4218_),
    .C(_4216_),
    .Y(\datapath.programcounter.pc_mux [5])
);

NAND2X1 _15479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [5]),
    .B(\datapath.programcounter.pc [6]),
    .Y(_4219_)
);

NOR2X1 _15480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4219_),
    .B(_4210_),
    .Y(_4220_)
);

AOI21X1 _15481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [5]),
    .B(_4211_),
    .C(\datapath.programcounter.pc [6]),
    .Y(_4221_)
);

NOR2X1 _15482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4220_),
    .B(_4221_),
    .Y(\datapath.nextpc [6])
);

NAND2X1 _15483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf3),
    .B(\datapath.nextpc [6]),
    .Y(_4222_)
);

NAND2X1 _15484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [6]),
    .B(_4196__bF$buf3),
    .Y(_4223_)
);

AOI22X1 _15485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf3),
    .B(_0_[6]),
    .C(\datapath.csr.csr_pcaddr [6]),
    .D(_4198__bF$buf3),
    .Y(_4224_)
);

NAND3X1 _15486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4223_),
    .B(_4224_),
    .C(_4222_),
    .Y(\datapath.programcounter.pc_mux [6])
);

OAI21X1 _15487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4210_),
    .B(_4219_),
    .C(_4141_),
    .Y(_4225_)
);

NAND2X1 _15488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [7]),
    .B(_4220_),
    .Y(_4226_)
);

AND2X2 _15489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4226_),
    .B(_4225_),
    .Y(\datapath.nextpc [7])
);

NAND2X1 _15490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf2),
    .B(\datapath.nextpc [7]),
    .Y(_4227_)
);

NAND2X1 _15491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [7]),
    .B(_4196__bF$buf2),
    .Y(_4228_)
);

AOI22X1 _15492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf2),
    .B(_0_[7]),
    .C(\datapath.csr.csr_pcaddr [7]),
    .D(_4198__bF$buf2),
    .Y(_4229_)
);

NAND3X1 _15493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4228_),
    .B(_4229_),
    .C(_4227_),
    .Y(\datapath.programcounter.pc_mux [7])
);

NAND3X1 _15494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [5]),
    .B(\datapath.programcounter.pc [6]),
    .C(\datapath.programcounter.pc [7]),
    .Y(_4230_)
);

OAI21X1 _15495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4210_),
    .B(_4230_),
    .C(_4143_),
    .Y(_4231_)
);

OR2X2 _15496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4210_),
    .B(_4230_),
    .Y(_4232_)
);

NOR2X1 _15497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4143_),
    .B(_4232_),
    .Y(_4233_)
);

INVX1 _15498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4233_),
    .Y(_4234_)
);

AND2X2 _15499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4234_),
    .B(_4231_),
    .Y(\datapath.nextpc [8])
);

NAND2X1 _15500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf1),
    .B(\datapath.nextpc [8]),
    .Y(_4235_)
);

NAND2X1 _15501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [8]),
    .B(_4196__bF$buf1),
    .Y(_4236_)
);

AOI22X1 _15502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf1),
    .B(_0_[8]),
    .C(\datapath.csr.csr_pcaddr [8]),
    .D(_4198__bF$buf1),
    .Y(_4237_)
);

NAND3X1 _15503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4236_),
    .B(_4237_),
    .C(_4235_),
    .Y(\datapath.programcounter.pc_mux [8])
);

XOR2X1 _15504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4233_),
    .B(\datapath.programcounter.pc [9]),
    .Y(\datapath.nextpc [9])
);

NAND2X1 _15505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf0),
    .B(\datapath.nextpc [9]),
    .Y(_4238_)
);

NAND2X1 _15506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [9]),
    .B(_4196__bF$buf0),
    .Y(_4239_)
);

AOI22X1 _15507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf0),
    .B(_0_[9]),
    .C(\datapath.csr.csr_pcaddr [9]),
    .D(_4198__bF$buf0),
    .Y(_4240_)
);

NAND3X1 _15508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4239_),
    .B(_4240_),
    .C(_4238_),
    .Y(\datapath.programcounter.pc_mux [9])
);

NAND2X1 _15509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [8]),
    .B(\datapath.programcounter.pc [9]),
    .Y(_4241_)
);

OAI21X1 _15510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4226_),
    .B(_4241_),
    .C(_4147_),
    .Y(_4242_)
);

NAND3X1 _15511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [9]),
    .B(\datapath.programcounter.pc [10]),
    .C(_4233_),
    .Y(_4243_)
);

AND2X2 _15512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4243_),
    .B(_4242_),
    .Y(\datapath.nextpc [10])
);

NAND2X1 _15513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf4),
    .B(\datapath.nextpc [10]),
    .Y(_4244_)
);

NAND2X1 _15514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [10]),
    .B(_4196__bF$buf4),
    .Y(_4245_)
);

AOI22X1 _15515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf4),
    .B(_0_[10]),
    .C(\datapath.csr.csr_pcaddr [10]),
    .D(_4198__bF$buf4),
    .Y(_4246_)
);

NAND3X1 _15516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4245_),
    .B(_4246_),
    .C(_4244_),
    .Y(\datapath.programcounter.pc_mux [10])
);

XNOR2X1 _15517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4243_),
    .B(\datapath.programcounter.pc [11]),
    .Y(\datapath.nextpc [11])
);

NAND2X1 _15518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf3),
    .B(\datapath.nextpc [11]),
    .Y(_4247_)
);

NAND2X1 _15519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [11]),
    .B(_4196__bF$buf3),
    .Y(_4248_)
);

AOI22X1 _15520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf3),
    .B(_0_[11]),
    .C(\datapath.csr.csr_pcaddr [11]),
    .D(_4198__bF$buf3),
    .Y(_4249_)
);

NAND3X1 _15521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4248_),
    .B(_4249_),
    .C(_4247_),
    .Y(\datapath.programcounter.pc_mux [11])
);

NAND2X1 _15522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [4]),
    .B(\datapath.programcounter.pc [5]),
    .Y(_4250_)
);

NAND2X1 _15523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [6]),
    .B(\datapath.programcounter.pc [7]),
    .Y(_4251_)
);

NOR2X1 _15524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4250_),
    .B(_4251_),
    .Y(_4252_)
);

NAND2X1 _15525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [10]),
    .B(\datapath.programcounter.pc [11]),
    .Y(_4253_)
);

NOR2X1 _15526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4241_),
    .B(_4253_),
    .Y(_4254_)
);

NAND3X1 _15527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4205_),
    .B(_4252_),
    .C(_4254_),
    .Y(_4255_)
);

XNOR2X1 _15528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4255_),
    .B(\datapath.programcounter.pc [12]),
    .Y(\datapath.nextpc [12])
);

NAND2X1 _15529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf2),
    .B(\datapath.nextpc [12]),
    .Y(_4256_)
);

NAND2X1 _15530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [12]),
    .B(_4196__bF$buf2),
    .Y(_4257_)
);

AOI22X1 _15531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf2),
    .B(_0_[12]),
    .C(\datapath.csr.csr_pcaddr [12]),
    .D(_4198__bF$buf2),
    .Y(_4258_)
);

NAND3X1 _15532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4257_),
    .B(_4258_),
    .C(_4256_),
    .Y(\datapath.programcounter.pc_mux [12])
);

NOR2X1 _15533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4210_),
    .B(_4230_),
    .Y(_4259_)
);

NAND3X1 _15534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [12]),
    .B(_4254_),
    .C(_4259_),
    .Y(_4260_)
);

AND2X2 _15535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4260_),
    .B(\datapath.programcounter.pc [13]),
    .Y(_4261_)
);

NOR2X1 _15536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [13]),
    .B(_4260_),
    .Y(_4262_)
);

OR2X2 _15537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4261_),
    .B(_4262_),
    .Y(\datapath.nextpc [13])
);

OAI21X1 _15538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4261_),
    .B(_4262_),
    .C(_4193__bF$buf1),
    .Y(_4263_)
);

NAND2X1 _15539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [13]),
    .B(_4196__bF$buf1),
    .Y(_4264_)
);

AOI22X1 _15540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf1),
    .B(_0_[13]),
    .C(\datapath.csr.csr_pcaddr [13]),
    .D(_4198__bF$buf1),
    .Y(_4265_)
);

NAND3X1 _15541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4264_),
    .B(_4265_),
    .C(_4263_),
    .Y(\datapath.programcounter.pc_mux [13])
);

OAI21X1 _15542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4260_),
    .B(_4153_),
    .C(_4155_),
    .Y(_4266_)
);

NOR2X1 _15543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4153_),
    .B(_4260_),
    .Y(_4267_)
);

NAND2X1 _15544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [14]),
    .B(_4267_),
    .Y(_4268_)
);

NAND2X1 _15545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4266_),
    .B(_4268_),
    .Y(_4269_)
);

INVX1 _15546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4269_),
    .Y(\datapath.nextpc [14])
);

INVX1 _15547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf0),
    .Y(_4270_)
);

NAND2X1 _15548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_pcaddr [14]),
    .B(_4198__bF$buf0),
    .Y(_4271_)
);

NAND2X1 _15549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[14]),
    .B(_4192__bF$buf0),
    .Y(_4272_)
);

NAND2X1 _15550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4272_),
    .B(_4271_),
    .Y(_4273_)
);

AOI21X1 _15551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [14]),
    .B(_4196__bF$buf0),
    .C(_4273_),
    .Y(_4274_)
);

OAI21X1 _15552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4269_),
    .B(_4270_),
    .C(_4274_),
    .Y(\datapath.programcounter.pc_mux [14])
);

NAND2X1 _15553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [12]),
    .B(\datapath.programcounter.pc [13]),
    .Y(_4275_)
);

NOR2X1 _15554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4275_),
    .B(_4255_),
    .Y(_4276_)
);

AOI21X1 _15555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [14]),
    .B(_4276_),
    .C(_4157_),
    .Y(_4277_)
);

NAND2X1 _15556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [14]),
    .B(_4276_),
    .Y(_4278_)
);

NOR2X1 _15557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [15]),
    .B(_4278_),
    .Y(_4279_)
);

OR2X2 _15558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4279_),
    .B(_4277_),
    .Y(\datapath.nextpc [15])
);

OAI21X1 _15559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4279_),
    .B(_4277_),
    .C(_4193__bF$buf4),
    .Y(_4280_)
);

NAND2X1 _15560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_pcaddr [15]),
    .B(_4198__bF$buf4),
    .Y(_4281_)
);

AOI22X1 _15561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf4),
    .B(_0_[15]),
    .C(\datapath.programcounter.jumps [15]),
    .D(_4196__bF$buf4),
    .Y(_4282_)
);

NAND3X1 _15562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4281_),
    .B(_4282_),
    .C(_4280_),
    .Y(\datapath.programcounter.pc_mux [15])
);

NAND2X1 _15563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [14]),
    .B(\datapath.programcounter.pc [15]),
    .Y(_4283_)
);

NOR2X1 _15564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4275_),
    .B(_4283_),
    .Y(_4284_)
);

NAND3X1 _15565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4254_),
    .B(_4284_),
    .C(_4259_),
    .Y(_4285_)
);

INVX1 _15566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4285_),
    .Y(_4286_)
);

NOR2X1 _15567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [16]),
    .B(_4286_),
    .Y(_4287_)
);

NOR2X1 _15568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4159_),
    .B(_4285_),
    .Y(_4288_)
);

NOR2X1 _15569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4288_),
    .B(_4287_),
    .Y(\datapath.nextpc [16])
);

NAND2X1 _15570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf3),
    .B(\datapath.nextpc [16]),
    .Y(_4289_)
);

NAND2X1 _15571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [16]),
    .B(_4196__bF$buf3),
    .Y(_4290_)
);

AOI22X1 _15572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf3),
    .B(_0_[16]),
    .C(\datapath.csr.csr_pcaddr [16]),
    .D(_4198__bF$buf3),
    .Y(_4291_)
);

NAND3X1 _15573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4290_),
    .B(_4291_),
    .C(_4289_),
    .Y(\datapath.programcounter.pc_mux [16])
);

XNOR2X1 _15574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4288_),
    .B(_4161_),
    .Y(\datapath.nextpc [17])
);

NAND2X1 _15575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf2),
    .B(\datapath.nextpc [17]),
    .Y(_4292_)
);

NAND2X1 _15576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [17]),
    .B(_4196__bF$buf2),
    .Y(_4293_)
);

AOI22X1 _15577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf2),
    .B(_0_[17]),
    .C(\datapath.csr.csr_pcaddr [17]),
    .D(_4198__bF$buf2),
    .Y(_4294_)
);

NAND3X1 _15578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4293_),
    .B(_4294_),
    .C(_4292_),
    .Y(\datapath.programcounter.pc_mux [17])
);

NAND3X1 _15579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [7]),
    .B(\datapath.programcounter.pc [14]),
    .C(\datapath.programcounter.pc [15]),
    .Y(_4295_)
);

NOR3X1 _15580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4219_),
    .B(_4275_),
    .C(_4295_),
    .Y(_4296_)
);

AND2X2 _15581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4254_),
    .B(_4211_),
    .Y(_4297_)
);

NAND2X1 _15582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4296_),
    .B(_4297_),
    .Y(_4298_)
);

NAND2X1 _15583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [16]),
    .B(\datapath.programcounter.pc [17]),
    .Y(_4299_)
);

OAI21X1 _15584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4298_),
    .B(_4299_),
    .C(_4163_),
    .Y(_4300_)
);

NAND3X1 _15585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [17]),
    .B(\datapath.programcounter.pc [18]),
    .C(_4288_),
    .Y(_4301_)
);

AND2X2 _15586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4301_),
    .B(_4300_),
    .Y(\datapath.nextpc [18])
);

NAND2X1 _15587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf1),
    .B(\datapath.nextpc [18]),
    .Y(_4302_)
);

NAND2X1 _15588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [18]),
    .B(_4196__bF$buf1),
    .Y(_4303_)
);

AOI22X1 _15589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf1),
    .B(_0_[18]),
    .C(\datapath.csr.csr_pcaddr [18]),
    .D(_4198__bF$buf1),
    .Y(_4304_)
);

NAND3X1 _15590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4303_),
    .B(_4304_),
    .C(_4302_),
    .Y(\datapath.programcounter.pc_mux [18])
);

OR2X2 _15591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4298_),
    .B(_4299_),
    .Y(_4305_)
);

OAI21X1 _15592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4305_),
    .B(_4163_),
    .C(_4165_),
    .Y(_4306_)
);

NOR2X1 _15593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4299_),
    .B(_4298_),
    .Y(_4307_)
);

NAND3X1 _15594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [18]),
    .B(\datapath.programcounter.pc [19]),
    .C(_4307_),
    .Y(_4308_)
);

AND2X2 _15595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4306_),
    .B(_4308_),
    .Y(\datapath.nextpc [19])
);

NAND3X1 _15596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf0),
    .B(_4308_),
    .C(_4306_),
    .Y(_4309_)
);

NAND2X1 _15597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [19]),
    .B(_4196__bF$buf0),
    .Y(_4310_)
);

AOI22X1 _15598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf0),
    .B(_0_[19]),
    .C(\datapath.csr.csr_pcaddr [19]),
    .D(_4198__bF$buf0),
    .Y(_4311_)
);

NAND3X1 _15599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4310_),
    .B(_4311_),
    .C(_4309_),
    .Y(\datapath.programcounter.pc_mux [19])
);

NAND2X1 _15600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [18]),
    .B(\datapath.programcounter.pc [19]),
    .Y(_4312_)
);

NOR2X1 _15601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4299_),
    .B(_4312_),
    .Y(_4313_)
);

NAND3X1 _15602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4296_),
    .B(_4313_),
    .C(_4297_),
    .Y(_4314_)
);

XNOR2X1 _15603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4314_),
    .B(\datapath.programcounter.pc [20]),
    .Y(\datapath.nextpc [20])
);

NAND2X1 _15604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf4),
    .B(\datapath.nextpc [20]),
    .Y(_4315_)
);

NAND2X1 _15605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [20]),
    .B(_4196__bF$buf4),
    .Y(_4316_)
);

AOI22X1 _15606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf4),
    .B(_0_[20]),
    .C(\datapath.csr.csr_pcaddr [20]),
    .D(_4198__bF$buf4),
    .Y(_4317_)
);

NAND3X1 _15607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4316_),
    .B(_4317_),
    .C(_4315_),
    .Y(\datapath.programcounter.pc_mux [20])
);

OAI21X1 _15608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4314_),
    .B(_4167_),
    .C(_4169_),
    .Y(_4318_)
);

INVX1 _15609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4314_),
    .Y(_4319_)
);

NAND2X1 _15610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [20]),
    .B(\datapath.programcounter.pc [21]),
    .Y(_4320_)
);

INVX1 _15611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4320_),
    .Y(_4321_)
);

NAND2X1 _15612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4321_),
    .B(_4319_),
    .Y(_4322_)
);

AND2X2 _15613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4322_),
    .B(_4318_),
    .Y(\datapath.nextpc [21])
);

NAND3X1 _15614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf3),
    .B(_4318_),
    .C(_4322_),
    .Y(_4323_)
);

NAND2X1 _15615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [21]),
    .B(_4196__bF$buf3),
    .Y(_4324_)
);

AOI22X1 _15616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf3),
    .B(_0_[21]),
    .C(\datapath.csr.csr_pcaddr [21]),
    .D(_4198__bF$buf3),
    .Y(_4325_)
);

NAND3X1 _15617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4324_),
    .B(_4325_),
    .C(_4323_),
    .Y(\datapath.programcounter.pc_mux [21])
);

OAI21X1 _15618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4314_),
    .B(_4320_),
    .C(_4171_),
    .Y(_4326_)
);

NOR3X1 _15619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4171_),
    .B(_4320_),
    .C(_4314_),
    .Y(_4327_)
);

INVX1 _15620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4327_),
    .Y(_4328_)
);

AND2X2 _15621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4328_),
    .B(_4326_),
    .Y(\datapath.nextpc [22])
);

NAND3X1 _15622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf2),
    .B(_4326_),
    .C(_4328_),
    .Y(_4329_)
);

NAND2X1 _15623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [22]),
    .B(_4196__bF$buf2),
    .Y(_4330_)
);

AOI22X1 _15624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf2),
    .B(_0_[22]),
    .C(\datapath.csr.csr_pcaddr [22]),
    .D(_4198__bF$buf2),
    .Y(_4331_)
);

NAND3X1 _15625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4330_),
    .B(_4331_),
    .C(_4329_),
    .Y(\datapath.programcounter.pc_mux [22])
);

XNOR2X1 _15626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4327_),
    .B(\datapath.programcounter.pc [23]),
    .Y(_4332_)
);

INVX1 _15627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4332_),
    .Y(\datapath.nextpc [23])
);

INVX1 _15628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [23]),
    .Y(_4333_)
);

INVX2 _15629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4196__bF$buf1),
    .Y(_4334_)
);

NAND2X1 _15630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_pcaddr [23]),
    .B(_4198__bF$buf1),
    .Y(_4335_)
);

OAI21X1 _15631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4334_),
    .B(_4333_),
    .C(_4335_),
    .Y(_4336_)
);

AOI21X1 _15632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[23]),
    .B(_4192__bF$buf1),
    .C(_4336_),
    .Y(_4337_)
);

OAI21X1 _15633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4332_),
    .B(_4270_),
    .C(_4337_),
    .Y(\datapath.programcounter.pc_mux [23])
);

NAND2X1 _15634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [22]),
    .B(\datapath.programcounter.pc [23]),
    .Y(_4338_)
);

NOR2X1 _15635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4320_),
    .B(_4338_),
    .Y(_4339_)
);

AND2X2 _15636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4313_),
    .B(_4339_),
    .Y(_4340_)
);

NAND3X1 _15637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4296_),
    .B(_4297_),
    .C(_4340_),
    .Y(_4341_)
);

XNOR2X1 _15638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4341_),
    .B(\datapath.programcounter.pc [24]),
    .Y(\datapath.nextpc [24])
);

NAND2X1 _15639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf1),
    .B(\datapath.nextpc [24]),
    .Y(_4342_)
);

NAND2X1 _15640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [24]),
    .B(_4196__bF$buf0),
    .Y(_4343_)
);

AOI22X1 _15641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf0),
    .B(_0_[24]),
    .C(\datapath.csr.csr_pcaddr [24]),
    .D(_4198__bF$buf0),
    .Y(_4344_)
);

NAND3X1 _15642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4343_),
    .B(_4344_),
    .C(_4342_),
    .Y(\datapath.programcounter.pc_mux [24])
);

OAI21X1 _15643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4341_),
    .B(_4175_),
    .C(_4177_),
    .Y(_4345_)
);

INVX1 _15644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4295_),
    .Y(_4346_)
);

NOR2X1 _15645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4219_),
    .B(_4275_),
    .Y(_4347_)
);

NAND2X1 _15646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4346_),
    .B(_4347_),
    .Y(_4348_)
);

NAND2X1 _15647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4211_),
    .B(_4254_),
    .Y(_4349_)
);

NAND2X1 _15648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4313_),
    .B(_4339_),
    .Y(_4350_)
);

NOR3X1 _15649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4348_),
    .B(_4349_),
    .C(_4350_),
    .Y(_4351_)
);

NAND3X1 _15650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [24]),
    .B(\datapath.programcounter.pc [25]),
    .C(_4351_),
    .Y(_4352_)
);

AND2X2 _15651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4345_),
    .B(_4352_),
    .Y(\datapath.nextpc [25])
);

NAND2X1 _15652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf0),
    .B(\datapath.nextpc [25]),
    .Y(_4353_)
);

NAND2X1 _15653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [25]),
    .B(_4196__bF$buf4),
    .Y(_4354_)
);

AOI22X1 _15654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf4),
    .B(_0_[25]),
    .C(\datapath.csr.csr_pcaddr [25]),
    .D(_4198__bF$buf4),
    .Y(_4355_)
);

NAND3X1 _15655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4354_),
    .B(_4355_),
    .C(_4353_),
    .Y(\datapath.programcounter.pc_mux [25])
);

NOR2X1 _15656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4175_),
    .B(_4177_),
    .Y(_4356_)
);

INVX2 _15657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4356_),
    .Y(_4357_)
);

OAI21X1 _15658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4341_),
    .B(_4357_),
    .C(_4179_),
    .Y(_4358_)
);

NOR2X1 _15659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4357_),
    .B(_4341_),
    .Y(_4359_)
);

NAND2X1 _15660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [26]),
    .B(_4359_),
    .Y(_4360_)
);

AND2X2 _15661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4360_),
    .B(_4358_),
    .Y(\datapath.nextpc [26])
);

NAND3X1 _15662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf4),
    .B(_4358_),
    .C(_4360_),
    .Y(_4361_)
);

NAND2X1 _15663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [26]),
    .B(_4196__bF$buf3),
    .Y(_4362_)
);

AOI22X1 _15664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf3),
    .B(_0_[26]),
    .C(\datapath.csr.csr_pcaddr [26]),
    .D(_4198__bF$buf3),
    .Y(_4363_)
);

NAND3X1 _15665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362_),
    .B(_4363_),
    .C(_4361_),
    .Y(\datapath.programcounter.pc_mux [26])
);

NAND2X1 _15666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4356_),
    .B(_4351_),
    .Y(_4364_)
);

OAI21X1 _15667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4364_),
    .B(_4179_),
    .C(_4181_),
    .Y(_4365_)
);

NAND3X1 _15668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [26]),
    .B(\datapath.programcounter.pc [27]),
    .C(_4359_),
    .Y(_4366_)
);

AND2X2 _15669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4366_),
    .B(_4365_),
    .Y(\datapath.nextpc [27])
);

NAND3X1 _15670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf3),
    .B(_4365_),
    .C(_4366_),
    .Y(_4367_)
);

NAND2X1 _15671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_pcaddr [27]),
    .B(_4198__bF$buf2),
    .Y(_4368_)
);

AOI22X1 _15672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf2),
    .B(_0_[27]),
    .C(\datapath.programcounter.jumps [27]),
    .D(_4196__bF$buf2),
    .Y(_4369_)
);

NAND3X1 _15673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4368_),
    .B(_4369_),
    .C(_4367_),
    .Y(\datapath.programcounter.pc_mux [27])
);

NAND2X1 _15674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [26]),
    .B(\datapath.programcounter.pc [27]),
    .Y(_4370_)
);

OR2X2 _15675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4357_),
    .B(_4370_),
    .Y(_4371_)
);

OAI21X1 _15676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4341_),
    .B(_4371_),
    .C(_4183_),
    .Y(_4372_)
);

NOR2X1 _15677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4371_),
    .B(_4341_),
    .Y(_4373_)
);

NAND2X1 _15678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [28]),
    .B(_4373_),
    .Y(_4374_)
);

AND2X2 _15679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4374_),
    .B(_4372_),
    .Y(\datapath.nextpc [28])
);

NAND3X1 _15680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf2),
    .B(_4372_),
    .C(_4374_),
    .Y(_4375_)
);

NAND2X1 _15681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [28]),
    .B(_4196__bF$buf1),
    .Y(_4376_)
);

AOI22X1 _15682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf1),
    .B(_0_[28]),
    .C(\datapath.csr.csr_pcaddr [28]),
    .D(_4198__bF$buf1),
    .Y(_4377_)
);

NAND3X1 _15683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4376_),
    .B(_4377_),
    .C(_4375_),
    .Y(\datapath.programcounter.pc_mux [28])
);

NOR2X1 _15684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4370_),
    .B(_4357_),
    .Y(_4378_)
);

NAND2X1 _15685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4378_),
    .B(_4351_),
    .Y(_4379_)
);

OAI21X1 _15686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4379_),
    .B(_4183_),
    .C(_4185_),
    .Y(_4380_)
);

NAND3X1 _15687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [28]),
    .B(\datapath.programcounter.pc [29]),
    .C(_4373_),
    .Y(_4381_)
);

AND2X2 _15688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4381_),
    .B(_4380_),
    .Y(\datapath.nextpc [29])
);

NAND3X1 _15689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf1),
    .B(_4380_),
    .C(_4381_),
    .Y(_4382_)
);

NAND2X1 _15690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_pcaddr [29]),
    .B(_4198__bF$buf0),
    .Y(_4383_)
);

AOI22X1 _15691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4192__bF$buf0),
    .B(_0_[29]),
    .C(\datapath.programcounter.jumps [29]),
    .D(_4196__bF$buf0),
    .Y(_4384_)
);

NAND3X1 _15692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4383_),
    .B(_4384_),
    .C(_4382_),
    .Y(\datapath.programcounter.pc_mux [29])
);

NAND2X1 _15693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [28]),
    .B(\datapath.programcounter.pc [29]),
    .Y(_4385_)
);

OAI21X1 _15694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4379_),
    .B(_4385_),
    .C(_4187_),
    .Y(_4386_)
);

NOR2X1 _15695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4350_),
    .B(_4285_),
    .Y(_4387_)
);

AND2X2 _15696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4387_),
    .B(_4378_),
    .Y(_4388_)
);

INVX1 _15697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4385_),
    .Y(_4389_)
);

NAND3X1 _15698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [30]),
    .B(_4389_),
    .C(_4388_),
    .Y(_4390_)
);

AND2X2 _15699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4390_),
    .B(_4386_),
    .Y(\datapath.nextpc [30])
);

NAND3X1 _15700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf0),
    .B(_4386_),
    .C(_4390_),
    .Y(_4391_)
);

INVX1 _15701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [30]),
    .Y(_4392_)
);

NAND2X1 _15702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[30]),
    .B(_4192__bF$buf4),
    .Y(_4393_)
);

OAI21X1 _15703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4334_),
    .B(_4392_),
    .C(_4393_),
    .Y(_4394_)
);

AOI21X1 _15704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_pcaddr [30]),
    .B(_4198__bF$buf4),
    .C(_4394_),
    .Y(_4395_)
);

NAND2X1 _15705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4395_),
    .B(_4391_),
    .Y(\datapath.programcounter.pc_mux [30])
);

NAND3X1 _15706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4378_),
    .B(_4389_),
    .C(_4351_),
    .Y(_4396_)
);

OAI21X1 _15707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4396_),
    .B(_4187_),
    .C(_4189_),
    .Y(_4397_)
);

NOR3X1 _15708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4371_),
    .B(_4385_),
    .C(_4341_),
    .Y(_4398_)
);

NAND3X1 _15709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [30]),
    .B(\datapath.programcounter.pc [31]),
    .C(_4398_),
    .Y(_4399_)
);

AND2X2 _15710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4399_),
    .B(_4397_),
    .Y(\datapath.nextpc [31])
);

NAND3X1 _15711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193__bF$buf4),
    .B(_4397_),
    .C(_4399_),
    .Y(_4400_)
);

INVX1 _15712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [31]),
    .Y(_4401_)
);

NAND2X1 _15713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_pcaddr [31]),
    .B(_4198__bF$buf3),
    .Y(_4402_)
);

OAI21X1 _15714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4334_),
    .B(_4401_),
    .C(_4402_),
    .Y(_4403_)
);

AOI21X1 _15715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[31]),
    .B(_4192__bF$buf3),
    .C(_4403_),
    .Y(_4404_)
);

NAND2X1 _15716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4404_),
    .B(_4400_),
    .Y(\datapath.programcounter.pc_mux [31])
);

DFFPOSX1 _15717_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf56),
    .D(\datapath.programcounter._1_ [0]),
    .Q(\datapath.programcounter.pc [0])
);

DFFPOSX1 _15718_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf55),
    .D(\datapath.programcounter._1_ [1]),
    .Q(\datapath.programcounter.pc [1])
);

DFFPOSX1 _15719_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf54),
    .D(\datapath.programcounter._1_ [2]),
    .Q(\datapath.programcounter.pc [2])
);

DFFPOSX1 _15720_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf53),
    .D(\datapath.programcounter._1_ [3]),
    .Q(\datapath.programcounter.pc [3])
);

DFFPOSX1 _15721_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf52),
    .D(\datapath.programcounter._1_ [4]),
    .Q(\datapath.programcounter.pc [4])
);

DFFPOSX1 _15722_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf51),
    .D(\datapath.programcounter._1_ [5]),
    .Q(\datapath.programcounter.pc [5])
);

DFFPOSX1 _15723_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf50),
    .D(\datapath.programcounter._1_ [6]),
    .Q(\datapath.programcounter.pc [6])
);

DFFPOSX1 _15724_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf49),
    .D(\datapath.programcounter._1_ [7]),
    .Q(\datapath.programcounter.pc [7])
);

DFFPOSX1 _15725_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf48),
    .D(\datapath.programcounter._1_ [8]),
    .Q(\datapath.programcounter.pc [8])
);

DFFPOSX1 _15726_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf47),
    .D(\datapath.programcounter._1_ [9]),
    .Q(\datapath.programcounter.pc [9])
);

DFFPOSX1 _15727_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf46),
    .D(\datapath.programcounter._1_ [10]),
    .Q(\datapath.programcounter.pc [10])
);

DFFPOSX1 _15728_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf45),
    .D(\datapath.programcounter._1_ [11]),
    .Q(\datapath.programcounter.pc [11])
);

DFFPOSX1 _15729_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf44),
    .D(\datapath.programcounter._1_ [12]),
    .Q(\datapath.programcounter.pc [12])
);

DFFPOSX1 _15730_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf43),
    .D(\datapath.programcounter._1_ [13]),
    .Q(\datapath.programcounter.pc [13])
);

DFFPOSX1 _15731_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf42),
    .D(\datapath.programcounter._1_ [14]),
    .Q(\datapath.programcounter.pc [14])
);

DFFPOSX1 _15732_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf41),
    .D(\datapath.programcounter._1_ [15]),
    .Q(\datapath.programcounter.pc [15])
);

DFFPOSX1 _15733_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf40),
    .D(\datapath.programcounter._1_ [16]),
    .Q(\datapath.programcounter.pc [16])
);

DFFPOSX1 _15734_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf39),
    .D(\datapath.programcounter._1_ [17]),
    .Q(\datapath.programcounter.pc [17])
);

DFFPOSX1 _15735_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf38),
    .D(\datapath.programcounter._1_ [18]),
    .Q(\datapath.programcounter.pc [18])
);

DFFPOSX1 _15736_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf37),
    .D(\datapath.programcounter._1_ [19]),
    .Q(\datapath.programcounter.pc [19])
);

DFFPOSX1 _15737_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf36),
    .D(\datapath.programcounter._1_ [20]),
    .Q(\datapath.programcounter.pc [20])
);

DFFPOSX1 _15738_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf35),
    .D(\datapath.programcounter._1_ [21]),
    .Q(\datapath.programcounter.pc [21])
);

DFFPOSX1 _15739_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf34),
    .D(\datapath.programcounter._1_ [22]),
    .Q(\datapath.programcounter.pc [22])
);

DFFPOSX1 _15740_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf33),
    .D(\datapath.programcounter._1_ [23]),
    .Q(\datapath.programcounter.pc [23])
);

DFFPOSX1 _15741_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf32),
    .D(\datapath.programcounter._1_ [24]),
    .Q(\datapath.programcounter.pc [24])
);

DFFPOSX1 _15742_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf31),
    .D(\datapath.programcounter._1_ [25]),
    .Q(\datapath.programcounter.pc [25])
);

DFFPOSX1 _15743_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf30),
    .D(\datapath.programcounter._1_ [26]),
    .Q(\datapath.programcounter.pc [26])
);

DFFPOSX1 _15744_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf29),
    .D(\datapath.programcounter._1_ [27]),
    .Q(\datapath.programcounter.pc [27])
);

DFFPOSX1 _15745_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf28),
    .D(\datapath.programcounter._1_ [28]),
    .Q(\datapath.programcounter.pc [28])
);

DFFPOSX1 _15746_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf27),
    .D(\datapath.programcounter._1_ [29]),
    .Q(\datapath.programcounter.pc [29])
);

DFFPOSX1 _15747_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf26),
    .D(\datapath.programcounter._1_ [30]),
    .Q(\datapath.programcounter.pc [30])
);

DFFPOSX1 _15748_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf25),
    .D(\datapath.programcounter._1_ [31]),
    .Q(\datapath.programcounter.pc [31])
);

INVX8 _15749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [0]),
    .Y(_5429_)
);

INVX2 _15750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [9]),
    .Y(_5430_)
);

NAND2X1 _15751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [11]),
    .B(\datapath.wbinstr [10]),
    .Y(_5431_)
);

OR2X2 _15752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5431_),
    .B(_5430_),
    .Y(_5432_)
);

INVX1 _15753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf10),
    .Y(_5433_)
);

NAND3X1 _15754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [8]),
    .B(\datapath.wbinstr [7]),
    .C(\controlunit.regfile_wen ),
    .Y(_5434_)
);

INVX4 _15755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5434__bF$buf14),
    .Y(_5435_)
);

NAND2X1 _15756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5435_),
    .B(_5433_),
    .Y(_5436_)
);

OAI21X1 _15757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf9),
    .B(_5434__bF$buf13),
    .C(\datapath.registers.1226[31] [0]),
    .Y(_5437_)
);

OAI21X1 _15758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf4),
    .B(_5429__bF$buf4),
    .C(_5437_),
    .Y(_5173_)
);

INVX8 _15759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [1]),
    .Y(_5438_)
);

OAI21X1 _15760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf8),
    .B(_5434__bF$buf12),
    .C(\datapath.registers.1226[31] [1]),
    .Y(_5439_)
);

OAI21X1 _15761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf3),
    .B(_5438__bF$buf4),
    .C(_5439_),
    .Y(_5184_)
);

INVX8 _15762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [2]),
    .Y(_5440_)
);

OAI21X1 _15763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf7),
    .B(_5434__bF$buf11),
    .C(\datapath.registers.1226[31] [2]),
    .Y(_5441_)
);

OAI21X1 _15764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf2),
    .B(_5440__bF$buf4),
    .C(_5441_),
    .Y(_5195_)
);

INVX8 _15765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [3]),
    .Y(_5442_)
);

OAI21X1 _15766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf6),
    .B(_5434__bF$buf10),
    .C(\datapath.registers.1226[31] [3]),
    .Y(_5443_)
);

OAI21X1 _15767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf1),
    .B(_5442__bF$buf4),
    .C(_5443_),
    .Y(_5198_)
);

INVX8 _15768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [4]),
    .Y(_5444_)
);

OAI21X1 _15769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf5),
    .B(_5434__bF$buf9),
    .C(\datapath.registers.1226[31] [4]),
    .Y(_5445_)
);

OAI21X1 _15770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf0),
    .B(_5444__bF$buf4),
    .C(_5445_),
    .Y(_5199_)
);

INVX8 _15771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [5]),
    .Y(_5446_)
);

OAI21X1 _15772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf4),
    .B(_5434__bF$buf8),
    .C(\datapath.registers.1226[31] [5]),
    .Y(_5447_)
);

OAI21X1 _15773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf4),
    .B(_5446__bF$buf4),
    .C(_5447_),
    .Y(_5200_)
);

INVX8 _15774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [6]),
    .Y(_5448_)
);

OAI21X1 _15775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf3),
    .B(_5434__bF$buf7),
    .C(\datapath.registers.1226[31] [6]),
    .Y(_5449_)
);

OAI21X1 _15776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf3),
    .B(_5448__bF$buf4),
    .C(_5449_),
    .Y(_5201_)
);

INVX8 _15777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [7]),
    .Y(_5450_)
);

OAI21X1 _15778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf2),
    .B(_5434__bF$buf6),
    .C(\datapath.registers.1226[31] [7]),
    .Y(_5451_)
);

OAI21X1 _15779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf2),
    .B(_5450__bF$buf4),
    .C(_5451_),
    .Y(_5202_)
);

INVX8 _15780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [8]),
    .Y(_5452_)
);

OAI21X1 _15781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf1),
    .B(_5434__bF$buf5),
    .C(\datapath.registers.1226[31] [8]),
    .Y(_5453_)
);

OAI21X1 _15782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf1),
    .B(_5452__bF$buf4),
    .C(_5453_),
    .Y(_5203_)
);

INVX8 _15783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [9]),
    .Y(_5454_)
);

OAI21X1 _15784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf0),
    .B(_5434__bF$buf4),
    .C(\datapath.registers.1226[31] [9]),
    .Y(_5455_)
);

OAI21X1 _15785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf0),
    .B(_5454__bF$buf4),
    .C(_5455_),
    .Y(_5204_)
);

INVX8 _15786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [10]),
    .Y(_5456_)
);

OAI21X1 _15787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf10),
    .B(_5434__bF$buf3),
    .C(\datapath.registers.1226[31] [10]),
    .Y(_5457_)
);

OAI21X1 _15788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf4),
    .B(_5456__bF$buf4),
    .C(_5457_),
    .Y(_5174_)
);

INVX8 _15789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [11]),
    .Y(_5458_)
);

OAI21X1 _15790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf9),
    .B(_5434__bF$buf2),
    .C(\datapath.registers.1226[31] [11]),
    .Y(_5459_)
);

OAI21X1 _15791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf3),
    .B(_5458__bF$buf4),
    .C(_5459_),
    .Y(_5175_)
);

INVX8 _15792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [12]),
    .Y(_5460_)
);

OAI21X1 _15793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf8),
    .B(_5434__bF$buf1),
    .C(\datapath.registers.1226[31] [12]),
    .Y(_5461_)
);

OAI21X1 _15794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf2),
    .B(_5460__bF$buf4),
    .C(_5461_),
    .Y(_5176_)
);

INVX8 _15795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [13]),
    .Y(_5462_)
);

OAI21X1 _15796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf7),
    .B(_5434__bF$buf0),
    .C(\datapath.registers.1226[31] [13]),
    .Y(_5463_)
);

OAI21X1 _15797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf1),
    .B(_5462__bF$buf4),
    .C(_5463_),
    .Y(_5177_)
);

INVX8 _15798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [14]),
    .Y(_5464_)
);

OAI21X1 _15799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf6),
    .B(_5434__bF$buf14),
    .C(\datapath.registers.1226[31] [14]),
    .Y(_5465_)
);

OAI21X1 _15800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf0),
    .B(_5464__bF$buf4),
    .C(_5465_),
    .Y(_5178_)
);

INVX8 _15801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [15]),
    .Y(_5466_)
);

OAI21X1 _15802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf5),
    .B(_5434__bF$buf13),
    .C(\datapath.registers.1226[31] [15]),
    .Y(_5467_)
);

OAI21X1 _15803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf4),
    .B(_5466__bF$buf4),
    .C(_5467_),
    .Y(_5179_)
);

INVX8 _15804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [16]),
    .Y(_5468_)
);

OAI21X1 _15805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf4),
    .B(_5434__bF$buf12),
    .C(\datapath.registers.1226[31] [16]),
    .Y(_5469_)
);

OAI21X1 _15806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf3),
    .B(_5468__bF$buf4),
    .C(_5469_),
    .Y(_5180_)
);

INVX8 _15807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [17]),
    .Y(_5470_)
);

OAI21X1 _15808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf3),
    .B(_5434__bF$buf11),
    .C(\datapath.registers.1226[31] [17]),
    .Y(_5471_)
);

OAI21X1 _15809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf2),
    .B(_5470__bF$buf4),
    .C(_5471_),
    .Y(_5181_)
);

INVX8 _15810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [18]),
    .Y(_5472_)
);

OAI21X1 _15811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf2),
    .B(_5434__bF$buf10),
    .C(\datapath.registers.1226[31] [18]),
    .Y(_5473_)
);

OAI21X1 _15812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf1),
    .B(_5472__bF$buf4),
    .C(_5473_),
    .Y(_5182_)
);

INVX8 _15813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [19]),
    .Y(_5474_)
);

OAI21X1 _15814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf1),
    .B(_5434__bF$buf9),
    .C(\datapath.registers.1226[31] [19]),
    .Y(_5475_)
);

OAI21X1 _15815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf0),
    .B(_5474__bF$buf4),
    .C(_5475_),
    .Y(_5183_)
);

INVX8 _15816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [20]),
    .Y(_5476_)
);

OAI21X1 _15817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf0),
    .B(_5434__bF$buf8),
    .C(\datapath.registers.1226[31] [20]),
    .Y(_5477_)
);

OAI21X1 _15818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf4),
    .B(_5476__bF$buf4),
    .C(_5477_),
    .Y(_5185_)
);

INVX8 _15819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [21]),
    .Y(_5478_)
);

OAI21X1 _15820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf10),
    .B(_5434__bF$buf7),
    .C(\datapath.registers.1226[31] [21]),
    .Y(_5479_)
);

OAI21X1 _15821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf3),
    .B(_5478__bF$buf4),
    .C(_5479_),
    .Y(_5186_)
);

INVX8 _15822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [22]),
    .Y(_5480_)
);

OAI21X1 _15823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf9),
    .B(_5434__bF$buf6),
    .C(\datapath.registers.1226[31] [22]),
    .Y(_5481_)
);

OAI21X1 _15824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf2),
    .B(_5480__bF$buf4),
    .C(_5481_),
    .Y(_5187_)
);

INVX8 _15825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [23]),
    .Y(_5482_)
);

OAI21X1 _15826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf8),
    .B(_5434__bF$buf5),
    .C(\datapath.registers.1226[31] [23]),
    .Y(_5483_)
);

OAI21X1 _15827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf1),
    .B(_5482__bF$buf4),
    .C(_5483_),
    .Y(_5188_)
);

INVX8 _15828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [24]),
    .Y(_5484_)
);

OAI21X1 _15829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf7),
    .B(_5434__bF$buf4),
    .C(\datapath.registers.1226[31] [24]),
    .Y(_5485_)
);

OAI21X1 _15830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf0),
    .B(_5484__bF$buf4),
    .C(_5485_),
    .Y(_5189_)
);

INVX8 _15831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [25]),
    .Y(_5486_)
);

OAI21X1 _15832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf6),
    .B(_5434__bF$buf3),
    .C(\datapath.registers.1226[31] [25]),
    .Y(_5487_)
);

OAI21X1 _15833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf4),
    .B(_5486__bF$buf4),
    .C(_5487_),
    .Y(_5190_)
);

INVX8 _15834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [26]),
    .Y(_5488_)
);

OAI21X1 _15835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf5),
    .B(_5434__bF$buf2),
    .C(\datapath.registers.1226[31] [26]),
    .Y(_5489_)
);

OAI21X1 _15836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf3),
    .B(_5488__bF$buf4),
    .C(_5489_),
    .Y(_5191_)
);

INVX8 _15837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [27]),
    .Y(_5490_)
);

OAI21X1 _15838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf4),
    .B(_5434__bF$buf1),
    .C(\datapath.registers.1226[31] [27]),
    .Y(_5491_)
);

OAI21X1 _15839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf2),
    .B(_5490__bF$buf4),
    .C(_5491_),
    .Y(_5192_)
);

INVX8 _15840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [28]),
    .Y(_5492_)
);

OAI21X1 _15841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf3),
    .B(_5434__bF$buf0),
    .C(\datapath.registers.1226[31] [28]),
    .Y(_5493_)
);

OAI21X1 _15842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf1),
    .B(_5492__bF$buf4),
    .C(_5493_),
    .Y(_5193_)
);

INVX8 _15843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [29]),
    .Y(_5494_)
);

OAI21X1 _15844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf2),
    .B(_5434__bF$buf14),
    .C(\datapath.registers.1226[31] [29]),
    .Y(_5495_)
);

OAI21X1 _15845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf0),
    .B(_5494__bF$buf4),
    .C(_5495_),
    .Y(_5194_)
);

INVX8 _15846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [30]),
    .Y(_5496_)
);

OAI21X1 _15847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf1),
    .B(_5434__bF$buf13),
    .C(\datapath.registers.1226[31] [30]),
    .Y(_5497_)
);

OAI21X1 _15848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf4),
    .B(_5496__bF$buf4),
    .C(_5497_),
    .Y(_5196_)
);

INVX8 _15849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [31]),
    .Y(_5498_)
);

OAI21X1 _15850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5432__bF$buf0),
    .B(_5434__bF$buf12),
    .C(\datapath.registers.1226[31] [31]),
    .Y(_5499_)
);

OAI21X1 _15851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436__bF$buf3),
    .B(_5498__bF$buf4),
    .C(_5499_),
    .Y(_5197_)
);

INVX1 _15852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [8]),
    .Y(_5500_)
);

INVX1 _15853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [7]),
    .Y(_5501_)
);

NAND2X1 _15854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5500_),
    .B(_5501_),
    .Y(_5502_)
);

INVX1 _15855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [11]),
    .Y(_5503_)
);

INVX2 _15856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [10]),
    .Y(_5504_)
);

NAND3X1 _15857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5503_),
    .B(_5504_),
    .C(_5430_),
    .Y(_5505_)
);

OAI21X1 _15858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5505__bF$buf7),
    .B(_5502_),
    .C(\controlunit.regfile_wen ),
    .Y(_5506_)
);

NAND2X1 _15859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [8]),
    .B(_5501_),
    .Y(_5507_)
);

NOR2X1 _15860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5507_),
    .B(_5506_),
    .Y(_5508_)
);

NAND2X1 _15861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5433_),
    .B(_5508_),
    .Y(_5509_)
);

INVX8 _15862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5508_),
    .Y(_5510_)
);

OAI21X1 _15863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf15),
    .B(_5432__bF$buf10),
    .C(\datapath.registers.1226[30] [0]),
    .Y(_5511_)
);

OAI21X1 _15864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf3),
    .B(_5509__bF$buf4),
    .C(_5511_),
    .Y(_5141_)
);

OAI21X1 _15865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf14),
    .B(_5432__bF$buf9),
    .C(\datapath.registers.1226[30] [1]),
    .Y(_5512_)
);

OAI21X1 _15866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf3),
    .B(_5509__bF$buf3),
    .C(_5512_),
    .Y(_5152_)
);

OAI21X1 _15867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf13),
    .B(_5432__bF$buf8),
    .C(\datapath.registers.1226[30] [2]),
    .Y(_5513_)
);

OAI21X1 _15868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf3),
    .B(_5509__bF$buf2),
    .C(_5513_),
    .Y(_5163_)
);

OAI21X1 _15869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf12),
    .B(_5432__bF$buf7),
    .C(\datapath.registers.1226[30] [3]),
    .Y(_5514_)
);

OAI21X1 _15870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf3),
    .B(_5509__bF$buf1),
    .C(_5514_),
    .Y(_5166_)
);

OAI21X1 _15871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf11),
    .B(_5432__bF$buf6),
    .C(\datapath.registers.1226[30] [4]),
    .Y(_5515_)
);

OAI21X1 _15872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf3),
    .B(_5509__bF$buf0),
    .C(_5515_),
    .Y(_5167_)
);

OAI21X1 _15873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf10),
    .B(_5432__bF$buf5),
    .C(\datapath.registers.1226[30] [5]),
    .Y(_5516_)
);

OAI21X1 _15874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf3),
    .B(_5509__bF$buf4),
    .C(_5516_),
    .Y(_5168_)
);

OAI21X1 _15875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf9),
    .B(_5432__bF$buf4),
    .C(\datapath.registers.1226[30] [6]),
    .Y(_5517_)
);

OAI21X1 _15876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf3),
    .B(_5509__bF$buf3),
    .C(_5517_),
    .Y(_5169_)
);

OAI21X1 _15877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf8),
    .B(_5432__bF$buf3),
    .C(\datapath.registers.1226[30] [7]),
    .Y(_5518_)
);

OAI21X1 _15878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf3),
    .B(_5509__bF$buf2),
    .C(_5518_),
    .Y(_5170_)
);

OAI21X1 _15879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf7),
    .B(_5432__bF$buf2),
    .C(\datapath.registers.1226[30] [8]),
    .Y(_5519_)
);

OAI21X1 _15880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf3),
    .B(_5509__bF$buf1),
    .C(_5519_),
    .Y(_5171_)
);

OAI21X1 _15881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf6),
    .B(_5432__bF$buf1),
    .C(\datapath.registers.1226[30] [9]),
    .Y(_5520_)
);

OAI21X1 _15882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf3),
    .B(_5509__bF$buf0),
    .C(_5520_),
    .Y(_5172_)
);

OAI21X1 _15883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf5),
    .B(_5432__bF$buf0),
    .C(\datapath.registers.1226[30] [10]),
    .Y(_5521_)
);

OAI21X1 _15884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf3),
    .B(_5509__bF$buf4),
    .C(_5521_),
    .Y(_5142_)
);

OAI21X1 _15885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf4),
    .B(_5432__bF$buf10),
    .C(\datapath.registers.1226[30] [11]),
    .Y(_5522_)
);

OAI21X1 _15886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf3),
    .B(_5509__bF$buf3),
    .C(_5522_),
    .Y(_5143_)
);

OAI21X1 _15887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf3),
    .B(_5432__bF$buf9),
    .C(\datapath.registers.1226[30] [12]),
    .Y(_5523_)
);

OAI21X1 _15888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf3),
    .B(_5509__bF$buf2),
    .C(_5523_),
    .Y(_5144_)
);

OAI21X1 _15889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf2),
    .B(_5432__bF$buf8),
    .C(\datapath.registers.1226[30] [13]),
    .Y(_5524_)
);

OAI21X1 _15890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf3),
    .B(_5509__bF$buf1),
    .C(_5524_),
    .Y(_5145_)
);

OAI21X1 _15891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf1),
    .B(_5432__bF$buf7),
    .C(\datapath.registers.1226[30] [14]),
    .Y(_5525_)
);

OAI21X1 _15892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf3),
    .B(_5509__bF$buf0),
    .C(_5525_),
    .Y(_5146_)
);

OAI21X1 _15893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf0),
    .B(_5432__bF$buf6),
    .C(\datapath.registers.1226[30] [15]),
    .Y(_5526_)
);

OAI21X1 _15894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf3),
    .B(_5509__bF$buf4),
    .C(_5526_),
    .Y(_5147_)
);

OAI21X1 _15895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf15),
    .B(_5432__bF$buf5),
    .C(\datapath.registers.1226[30] [16]),
    .Y(_5527_)
);

OAI21X1 _15896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf3),
    .B(_5509__bF$buf3),
    .C(_5527_),
    .Y(_5148_)
);

OAI21X1 _15897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf14),
    .B(_5432__bF$buf4),
    .C(\datapath.registers.1226[30] [17]),
    .Y(_5528_)
);

OAI21X1 _15898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf3),
    .B(_5509__bF$buf2),
    .C(_5528_),
    .Y(_5149_)
);

OAI21X1 _15899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf13),
    .B(_5432__bF$buf3),
    .C(\datapath.registers.1226[30] [18]),
    .Y(_5529_)
);

OAI21X1 _15900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf3),
    .B(_5509__bF$buf1),
    .C(_5529_),
    .Y(_5150_)
);

OAI21X1 _15901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf12),
    .B(_5432__bF$buf2),
    .C(\datapath.registers.1226[30] [19]),
    .Y(_5530_)
);

OAI21X1 _15902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf3),
    .B(_5509__bF$buf0),
    .C(_5530_),
    .Y(_5151_)
);

OAI21X1 _15903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf11),
    .B(_5432__bF$buf1),
    .C(\datapath.registers.1226[30] [20]),
    .Y(_5531_)
);

OAI21X1 _15904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf3),
    .B(_5509__bF$buf4),
    .C(_5531_),
    .Y(_5153_)
);

OAI21X1 _15905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf10),
    .B(_5432__bF$buf0),
    .C(\datapath.registers.1226[30] [21]),
    .Y(_5532_)
);

OAI21X1 _15906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf3),
    .B(_5509__bF$buf3),
    .C(_5532_),
    .Y(_5154_)
);

OAI21X1 _15907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf9),
    .B(_5432__bF$buf10),
    .C(\datapath.registers.1226[30] [22]),
    .Y(_5533_)
);

OAI21X1 _15908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf3),
    .B(_5509__bF$buf2),
    .C(_5533_),
    .Y(_5155_)
);

OAI21X1 _15909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf8),
    .B(_5432__bF$buf9),
    .C(\datapath.registers.1226[30] [23]),
    .Y(_5534_)
);

OAI21X1 _15910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf3),
    .B(_5509__bF$buf1),
    .C(_5534_),
    .Y(_5156_)
);

OAI21X1 _15911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf7),
    .B(_5432__bF$buf8),
    .C(\datapath.registers.1226[30] [24]),
    .Y(_5535_)
);

OAI21X1 _15912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf3),
    .B(_5509__bF$buf0),
    .C(_5535_),
    .Y(_5157_)
);

OAI21X1 _15913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf6),
    .B(_5432__bF$buf7),
    .C(\datapath.registers.1226[30] [25]),
    .Y(_5536_)
);

OAI21X1 _15914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486__bF$buf3),
    .B(_5509__bF$buf4),
    .C(_5536_),
    .Y(_5158_)
);

OAI21X1 _15915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf5),
    .B(_5432__bF$buf6),
    .C(\datapath.registers.1226[30] [26]),
    .Y(_5537_)
);

OAI21X1 _15916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf3),
    .B(_5509__bF$buf3),
    .C(_5537_),
    .Y(_5159_)
);

OAI21X1 _15917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf4),
    .B(_5432__bF$buf5),
    .C(\datapath.registers.1226[30] [27]),
    .Y(_5538_)
);

OAI21X1 _15918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf3),
    .B(_5509__bF$buf2),
    .C(_5538_),
    .Y(_5160_)
);

OAI21X1 _15919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf3),
    .B(_5432__bF$buf4),
    .C(\datapath.registers.1226[30] [28]),
    .Y(_5539_)
);

OAI21X1 _15920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf3),
    .B(_5509__bF$buf1),
    .C(_5539_),
    .Y(_5161_)
);

OAI21X1 _15921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf2),
    .B(_5432__bF$buf3),
    .C(\datapath.registers.1226[30] [29]),
    .Y(_5540_)
);

OAI21X1 _15922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf3),
    .B(_5509__bF$buf0),
    .C(_5540_),
    .Y(_5162_)
);

OAI21X1 _15923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf1),
    .B(_5432__bF$buf2),
    .C(\datapath.registers.1226[30] [30]),
    .Y(_5541_)
);

OAI21X1 _15924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf3),
    .B(_5509__bF$buf4),
    .C(_5541_),
    .Y(_5164_)
);

OAI21X1 _15925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf0),
    .B(_5432__bF$buf1),
    .C(\datapath.registers.1226[30] [31]),
    .Y(_5542_)
);

OAI21X1 _15926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf3),
    .B(_5509__bF$buf3),
    .C(_5542_),
    .Y(_5165_)
);

NAND2X1 _15927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.regfile_wen ),
    .B(_5500_),
    .Y(_5543_)
);

NOR2X1 _15928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5501_),
    .B(_5543_),
    .Y(_5544_)
);

NAND2X1 _15929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5544_),
    .B(_5433_),
    .Y(_5545_)
);

INVX8 _15930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5544_),
    .Y(_5546_)
);

OAI21X1 _15931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf15),
    .B(_5432__bF$buf0),
    .C(\datapath.registers.1226[29] [0]),
    .Y(_5547_)
);

OAI21X1 _15932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf4),
    .B(_5429__bF$buf2),
    .C(_5547_),
    .Y(_5077_)
);

OAI21X1 _15933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf14),
    .B(_5432__bF$buf10),
    .C(\datapath.registers.1226[29] [1]),
    .Y(_5548_)
);

OAI21X1 _15934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf3),
    .B(_5438__bF$buf2),
    .C(_5548_),
    .Y(_5088_)
);

OAI21X1 _15935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf13),
    .B(_5432__bF$buf9),
    .C(\datapath.registers.1226[29] [2]),
    .Y(_5549_)
);

OAI21X1 _15936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf2),
    .B(_5440__bF$buf2),
    .C(_5549_),
    .Y(_5099_)
);

OAI21X1 _15937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf12),
    .B(_5432__bF$buf8),
    .C(\datapath.registers.1226[29] [3]),
    .Y(_5550_)
);

OAI21X1 _15938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf1),
    .B(_5442__bF$buf2),
    .C(_5550_),
    .Y(_5102_)
);

OAI21X1 _15939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf11),
    .B(_5432__bF$buf7),
    .C(\datapath.registers.1226[29] [4]),
    .Y(_5551_)
);

OAI21X1 _15940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf0),
    .B(_5444__bF$buf2),
    .C(_5551_),
    .Y(_5103_)
);

OAI21X1 _15941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf10),
    .B(_5432__bF$buf6),
    .C(\datapath.registers.1226[29] [5]),
    .Y(_5552_)
);

OAI21X1 _15942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf4),
    .B(_5446__bF$buf2),
    .C(_5552_),
    .Y(_5104_)
);

OAI21X1 _15943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf9),
    .B(_5432__bF$buf5),
    .C(\datapath.registers.1226[29] [6]),
    .Y(_5553_)
);

OAI21X1 _15944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf3),
    .B(_5448__bF$buf2),
    .C(_5553_),
    .Y(_5105_)
);

OAI21X1 _15945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf8),
    .B(_5432__bF$buf4),
    .C(\datapath.registers.1226[29] [7]),
    .Y(_5554_)
);

OAI21X1 _15946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf2),
    .B(_5450__bF$buf2),
    .C(_5554_),
    .Y(_5106_)
);

OAI21X1 _15947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf7),
    .B(_5432__bF$buf3),
    .C(\datapath.registers.1226[29] [8]),
    .Y(_5555_)
);

OAI21X1 _15948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf1),
    .B(_5452__bF$buf2),
    .C(_5555_),
    .Y(_5107_)
);

OAI21X1 _15949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf6),
    .B(_5432__bF$buf2),
    .C(\datapath.registers.1226[29] [9]),
    .Y(_5556_)
);

OAI21X1 _15950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf0),
    .B(_5454__bF$buf2),
    .C(_5556_),
    .Y(_5108_)
);

OAI21X1 _15951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf5),
    .B(_5432__bF$buf1),
    .C(\datapath.registers.1226[29] [10]),
    .Y(_5557_)
);

OAI21X1 _15952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf4),
    .B(_5456__bF$buf2),
    .C(_5557_),
    .Y(_5078_)
);

OAI21X1 _15953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf4),
    .B(_5432__bF$buf0),
    .C(\datapath.registers.1226[29] [11]),
    .Y(_5558_)
);

OAI21X1 _15954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf3),
    .B(_5458__bF$buf2),
    .C(_5558_),
    .Y(_5079_)
);

OAI21X1 _15955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf3),
    .B(_5432__bF$buf10),
    .C(\datapath.registers.1226[29] [12]),
    .Y(_5559_)
);

OAI21X1 _15956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf2),
    .B(_5460__bF$buf2),
    .C(_5559_),
    .Y(_5080_)
);

OAI21X1 _15957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf2),
    .B(_5432__bF$buf9),
    .C(\datapath.registers.1226[29] [13]),
    .Y(_5560_)
);

OAI21X1 _15958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf1),
    .B(_5462__bF$buf2),
    .C(_5560_),
    .Y(_5081_)
);

OAI21X1 _15959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf1),
    .B(_5432__bF$buf8),
    .C(\datapath.registers.1226[29] [14]),
    .Y(_5561_)
);

OAI21X1 _15960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf0),
    .B(_5464__bF$buf2),
    .C(_5561_),
    .Y(_5082_)
);

OAI21X1 _15961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf0),
    .B(_5432__bF$buf7),
    .C(\datapath.registers.1226[29] [15]),
    .Y(_5562_)
);

OAI21X1 _15962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf4),
    .B(_5466__bF$buf2),
    .C(_5562_),
    .Y(_5083_)
);

OAI21X1 _15963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf15),
    .B(_5432__bF$buf6),
    .C(\datapath.registers.1226[29] [16]),
    .Y(_5563_)
);

OAI21X1 _15964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf3),
    .B(_5468__bF$buf2),
    .C(_5563_),
    .Y(_5084_)
);

OAI21X1 _15965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf14),
    .B(_5432__bF$buf5),
    .C(\datapath.registers.1226[29] [17]),
    .Y(_5564_)
);

OAI21X1 _15966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf2),
    .B(_5470__bF$buf2),
    .C(_5564_),
    .Y(_5085_)
);

OAI21X1 _15967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf13),
    .B(_5432__bF$buf4),
    .C(\datapath.registers.1226[29] [18]),
    .Y(_5565_)
);

OAI21X1 _15968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf1),
    .B(_5472__bF$buf2),
    .C(_5565_),
    .Y(_5086_)
);

OAI21X1 _15969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf12),
    .B(_5432__bF$buf3),
    .C(\datapath.registers.1226[29] [19]),
    .Y(_5566_)
);

OAI21X1 _15970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf0),
    .B(_5474__bF$buf2),
    .C(_5566_),
    .Y(_5087_)
);

OAI21X1 _15971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf11),
    .B(_5432__bF$buf2),
    .C(\datapath.registers.1226[29] [20]),
    .Y(_5567_)
);

OAI21X1 _15972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf4),
    .B(_5476__bF$buf2),
    .C(_5567_),
    .Y(_5089_)
);

OAI21X1 _15973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf10),
    .B(_5432__bF$buf1),
    .C(\datapath.registers.1226[29] [21]),
    .Y(_5568_)
);

OAI21X1 _15974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf3),
    .B(_5478__bF$buf2),
    .C(_5568_),
    .Y(_5090_)
);

OAI21X1 _15975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf9),
    .B(_5432__bF$buf0),
    .C(\datapath.registers.1226[29] [22]),
    .Y(_5569_)
);

OAI21X1 _15976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf2),
    .B(_5480__bF$buf2),
    .C(_5569_),
    .Y(_5091_)
);

OAI21X1 _15977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf8),
    .B(_5432__bF$buf10),
    .C(\datapath.registers.1226[29] [23]),
    .Y(_5570_)
);

OAI21X1 _15978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf1),
    .B(_5482__bF$buf2),
    .C(_5570_),
    .Y(_5092_)
);

OAI21X1 _15979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf7),
    .B(_5432__bF$buf9),
    .C(\datapath.registers.1226[29] [24]),
    .Y(_5571_)
);

OAI21X1 _15980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf0),
    .B(_5484__bF$buf2),
    .C(_5571_),
    .Y(_5093_)
);

OAI21X1 _15981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf6),
    .B(_5432__bF$buf8),
    .C(\datapath.registers.1226[29] [25]),
    .Y(_5572_)
);

OAI21X1 _15982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf4),
    .B(_5486__bF$buf2),
    .C(_5572_),
    .Y(_5094_)
);

OAI21X1 _15983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf5),
    .B(_5432__bF$buf7),
    .C(\datapath.registers.1226[29] [26]),
    .Y(_5573_)
);

OAI21X1 _15984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf3),
    .B(_5488__bF$buf2),
    .C(_5573_),
    .Y(_5095_)
);

OAI21X1 _15985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf4),
    .B(_5432__bF$buf6),
    .C(\datapath.registers.1226[29] [27]),
    .Y(_5574_)
);

OAI21X1 _15986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf2),
    .B(_5490__bF$buf2),
    .C(_5574_),
    .Y(_5096_)
);

OAI21X1 _15987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf3),
    .B(_5432__bF$buf5),
    .C(\datapath.registers.1226[29] [28]),
    .Y(_5575_)
);

OAI21X1 _15988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf1),
    .B(_5492__bF$buf2),
    .C(_5575_),
    .Y(_5097_)
);

OAI21X1 _15989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf2),
    .B(_5432__bF$buf4),
    .C(\datapath.registers.1226[29] [29]),
    .Y(_5576_)
);

OAI21X1 _15990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf0),
    .B(_5494__bF$buf2),
    .C(_5576_),
    .Y(_5098_)
);

OAI21X1 _15991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf1),
    .B(_5432__bF$buf3),
    .C(\datapath.registers.1226[29] [30]),
    .Y(_5577_)
);

OAI21X1 _15992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf4),
    .B(_5496__bF$buf2),
    .C(_5577_),
    .Y(_5100_)
);

OAI21X1 _15993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf0),
    .B(_5432__bF$buf2),
    .C(\datapath.registers.1226[29] [31]),
    .Y(_5578_)
);

OAI21X1 _15994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545__bF$buf3),
    .B(_5498__bF$buf2),
    .C(_5578_),
    .Y(_5101_)
);

OR2X2 _15995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5543_),
    .B(\datapath.wbinstr [7]),
    .Y(_5579_)
);

OR2X2 _15996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf5),
    .B(_5432__bF$buf1),
    .Y(_5580_)
);

OAI21X1 _15997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf4),
    .B(_5432__bF$buf0),
    .C(\datapath.registers.1226[28] [0]),
    .Y(_5581_)
);

OAI21X1 _15998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf4),
    .B(_5429__bF$buf1),
    .C(_5581_),
    .Y(_5045_)
);

OAI21X1 _15999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf3),
    .B(_5432__bF$buf10),
    .C(\datapath.registers.1226[28] [1]),
    .Y(_5582_)
);

OAI21X1 _16000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf3),
    .B(_5438__bF$buf1),
    .C(_5582_),
    .Y(_5056_)
);

OAI21X1 _16001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf2),
    .B(_5432__bF$buf9),
    .C(\datapath.registers.1226[28] [2]),
    .Y(_5583_)
);

OAI21X1 _16002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf2),
    .B(_5440__bF$buf1),
    .C(_5583_),
    .Y(_5067_)
);

OAI21X1 _16003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf1),
    .B(_5432__bF$buf8),
    .C(\datapath.registers.1226[28] [3]),
    .Y(_5584_)
);

OAI21X1 _16004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf1),
    .B(_5442__bF$buf1),
    .C(_5584_),
    .Y(_5070_)
);

OAI21X1 _16005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf0),
    .B(_5432__bF$buf7),
    .C(\datapath.registers.1226[28] [4]),
    .Y(_5585_)
);

OAI21X1 _16006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf0),
    .B(_5444__bF$buf1),
    .C(_5585_),
    .Y(_5071_)
);

OAI21X1 _16007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf5),
    .B(_5432__bF$buf6),
    .C(\datapath.registers.1226[28] [5]),
    .Y(_5586_)
);

OAI21X1 _16008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf4),
    .B(_5446__bF$buf1),
    .C(_5586_),
    .Y(_5072_)
);

OAI21X1 _16009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf4),
    .B(_5432__bF$buf5),
    .C(\datapath.registers.1226[28] [6]),
    .Y(_5587_)
);

OAI21X1 _16010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf3),
    .B(_5448__bF$buf1),
    .C(_5587_),
    .Y(_5073_)
);

OAI21X1 _16011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf3),
    .B(_5432__bF$buf4),
    .C(\datapath.registers.1226[28] [7]),
    .Y(_5588_)
);

OAI21X1 _16012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf2),
    .B(_5450__bF$buf1),
    .C(_5588_),
    .Y(_5074_)
);

OAI21X1 _16013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf2),
    .B(_5432__bF$buf3),
    .C(\datapath.registers.1226[28] [8]),
    .Y(_5589_)
);

OAI21X1 _16014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf1),
    .B(_5452__bF$buf1),
    .C(_5589_),
    .Y(_5075_)
);

OAI21X1 _16015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf1),
    .B(_5432__bF$buf2),
    .C(\datapath.registers.1226[28] [9]),
    .Y(_5590_)
);

OAI21X1 _16016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf0),
    .B(_5454__bF$buf1),
    .C(_5590_),
    .Y(_5076_)
);

OAI21X1 _16017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf0),
    .B(_5432__bF$buf1),
    .C(\datapath.registers.1226[28] [10]),
    .Y(_5591_)
);

OAI21X1 _16018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf4),
    .B(_5456__bF$buf1),
    .C(_5591_),
    .Y(_5046_)
);

OAI21X1 _16019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf5),
    .B(_5432__bF$buf0),
    .C(\datapath.registers.1226[28] [11]),
    .Y(_5592_)
);

OAI21X1 _16020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf3),
    .B(_5458__bF$buf1),
    .C(_5592_),
    .Y(_5047_)
);

OAI21X1 _16021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf4),
    .B(_5432__bF$buf10),
    .C(\datapath.registers.1226[28] [12]),
    .Y(_5593_)
);

OAI21X1 _16022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf2),
    .B(_5460__bF$buf1),
    .C(_5593_),
    .Y(_5048_)
);

OAI21X1 _16023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf3),
    .B(_5432__bF$buf9),
    .C(\datapath.registers.1226[28] [13]),
    .Y(_5594_)
);

OAI21X1 _16024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf1),
    .B(_5462__bF$buf1),
    .C(_5594_),
    .Y(_5049_)
);

OAI21X1 _16025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf2),
    .B(_5432__bF$buf8),
    .C(\datapath.registers.1226[28] [14]),
    .Y(_5595_)
);

OAI21X1 _16026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf0),
    .B(_5464__bF$buf1),
    .C(_5595_),
    .Y(_5050_)
);

OAI21X1 _16027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf1),
    .B(_5432__bF$buf7),
    .C(\datapath.registers.1226[28] [15]),
    .Y(_5596_)
);

OAI21X1 _16028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf4),
    .B(_5466__bF$buf1),
    .C(_5596_),
    .Y(_5051_)
);

OAI21X1 _16029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf0),
    .B(_5432__bF$buf6),
    .C(\datapath.registers.1226[28] [16]),
    .Y(_5597_)
);

OAI21X1 _16030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf3),
    .B(_5468__bF$buf1),
    .C(_5597_),
    .Y(_5052_)
);

OAI21X1 _16031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf5),
    .B(_5432__bF$buf5),
    .C(\datapath.registers.1226[28] [17]),
    .Y(_5598_)
);

OAI21X1 _16032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf2),
    .B(_5470__bF$buf1),
    .C(_5598_),
    .Y(_5053_)
);

OAI21X1 _16033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf4),
    .B(_5432__bF$buf4),
    .C(\datapath.registers.1226[28] [18]),
    .Y(_5599_)
);

OAI21X1 _16034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf1),
    .B(_5472__bF$buf1),
    .C(_5599_),
    .Y(_5054_)
);

OAI21X1 _16035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf3),
    .B(_5432__bF$buf3),
    .C(\datapath.registers.1226[28] [19]),
    .Y(_5600_)
);

OAI21X1 _16036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf0),
    .B(_5474__bF$buf1),
    .C(_5600_),
    .Y(_5055_)
);

OAI21X1 _16037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf2),
    .B(_5432__bF$buf2),
    .C(\datapath.registers.1226[28] [20]),
    .Y(_5601_)
);

OAI21X1 _16038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf4),
    .B(_5476__bF$buf1),
    .C(_5601_),
    .Y(_5057_)
);

OAI21X1 _16039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf1),
    .B(_5432__bF$buf1),
    .C(\datapath.registers.1226[28] [21]),
    .Y(_5602_)
);

OAI21X1 _16040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf3),
    .B(_5478__bF$buf1),
    .C(_5602_),
    .Y(_5058_)
);

OAI21X1 _16041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf0),
    .B(_5432__bF$buf0),
    .C(\datapath.registers.1226[28] [22]),
    .Y(_5603_)
);

OAI21X1 _16042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf2),
    .B(_5480__bF$buf1),
    .C(_5603_),
    .Y(_5059_)
);

OAI21X1 _16043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf5),
    .B(_5432__bF$buf10),
    .C(\datapath.registers.1226[28] [23]),
    .Y(_5604_)
);

OAI21X1 _16044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf1),
    .B(_5482__bF$buf1),
    .C(_5604_),
    .Y(_5060_)
);

OAI21X1 _16045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf4),
    .B(_5432__bF$buf9),
    .C(\datapath.registers.1226[28] [24]),
    .Y(_5605_)
);

OAI21X1 _16046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf0),
    .B(_5484__bF$buf1),
    .C(_5605_),
    .Y(_5061_)
);

OAI21X1 _16047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf3),
    .B(_5432__bF$buf8),
    .C(\datapath.registers.1226[28] [25]),
    .Y(_5606_)
);

OAI21X1 _16048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf4),
    .B(_5486__bF$buf1),
    .C(_5606_),
    .Y(_5062_)
);

OAI21X1 _16049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf2),
    .B(_5432__bF$buf7),
    .C(\datapath.registers.1226[28] [26]),
    .Y(_5607_)
);

OAI21X1 _16050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf3),
    .B(_5488__bF$buf1),
    .C(_5607_),
    .Y(_5063_)
);

OAI21X1 _16051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf1),
    .B(_5432__bF$buf6),
    .C(\datapath.registers.1226[28] [27]),
    .Y(_5608_)
);

OAI21X1 _16052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf2),
    .B(_5490__bF$buf1),
    .C(_5608_),
    .Y(_5064_)
);

OAI21X1 _16053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf0),
    .B(_5432__bF$buf5),
    .C(\datapath.registers.1226[28] [28]),
    .Y(_5609_)
);

OAI21X1 _16054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf1),
    .B(_5492__bF$buf1),
    .C(_5609_),
    .Y(_5065_)
);

OAI21X1 _16055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf5),
    .B(_5432__bF$buf4),
    .C(\datapath.registers.1226[28] [29]),
    .Y(_5610_)
);

OAI21X1 _16056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf0),
    .B(_5494__bF$buf1),
    .C(_5610_),
    .Y(_5066_)
);

OAI21X1 _16057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf4),
    .B(_5432__bF$buf3),
    .C(\datapath.registers.1226[28] [30]),
    .Y(_5611_)
);

OAI21X1 _16058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf4),
    .B(_5496__bF$buf1),
    .C(_5611_),
    .Y(_5068_)
);

OAI21X1 _16059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf3),
    .B(_5432__bF$buf2),
    .C(\datapath.registers.1226[28] [31]),
    .Y(_5612_)
);

OAI21X1 _16060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5580__bF$buf3),
    .B(_5498__bF$buf1),
    .C(_5612_),
    .Y(_5069_)
);

NOR2X1 _16061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [9]),
    .B(_5431_),
    .Y(_5613_)
);

NAND2X1 _16062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5435_),
    .B(_5613_),
    .Y(_5614_)
);

INVX8 _16063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5613_),
    .Y(_5615_)
);

OAI21X1 _16064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf8),
    .B(_5434__bF$buf11),
    .C(\datapath.registers.1226[27] [0]),
    .Y(_5616_)
);

OAI21X1 _16065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf4),
    .B(_5429__bF$buf0),
    .C(_5616_),
    .Y(_5013_)
);

OAI21X1 _16066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf7),
    .B(_5434__bF$buf10),
    .C(\datapath.registers.1226[27] [1]),
    .Y(_5617_)
);

OAI21X1 _16067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf3),
    .B(_5438__bF$buf0),
    .C(_5617_),
    .Y(_5024_)
);

OAI21X1 _16068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf6),
    .B(_5434__bF$buf9),
    .C(\datapath.registers.1226[27] [2]),
    .Y(_5618_)
);

OAI21X1 _16069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf2),
    .B(_5440__bF$buf0),
    .C(_5618_),
    .Y(_5035_)
);

OAI21X1 _16070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf5),
    .B(_5434__bF$buf8),
    .C(\datapath.registers.1226[27] [3]),
    .Y(_5619_)
);

OAI21X1 _16071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf1),
    .B(_5442__bF$buf0),
    .C(_5619_),
    .Y(_5038_)
);

OAI21X1 _16072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf4),
    .B(_5434__bF$buf7),
    .C(\datapath.registers.1226[27] [4]),
    .Y(_5620_)
);

OAI21X1 _16073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf0),
    .B(_5444__bF$buf0),
    .C(_5620_),
    .Y(_5039_)
);

OAI21X1 _16074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf3),
    .B(_5434__bF$buf6),
    .C(\datapath.registers.1226[27] [5]),
    .Y(_5621_)
);

OAI21X1 _16075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf4),
    .B(_5446__bF$buf0),
    .C(_5621_),
    .Y(_5040_)
);

OAI21X1 _16076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf2),
    .B(_5434__bF$buf5),
    .C(\datapath.registers.1226[27] [6]),
    .Y(_5622_)
);

OAI21X1 _16077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf3),
    .B(_5448__bF$buf0),
    .C(_5622_),
    .Y(_5041_)
);

OAI21X1 _16078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf1),
    .B(_5434__bF$buf4),
    .C(\datapath.registers.1226[27] [7]),
    .Y(_5623_)
);

OAI21X1 _16079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf2),
    .B(_5450__bF$buf0),
    .C(_5623_),
    .Y(_5042_)
);

OAI21X1 _16080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf0),
    .B(_5434__bF$buf3),
    .C(\datapath.registers.1226[27] [8]),
    .Y(_5624_)
);

OAI21X1 _16081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf1),
    .B(_5452__bF$buf0),
    .C(_5624_),
    .Y(_5043_)
);

OAI21X1 _16082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf8),
    .B(_5434__bF$buf2),
    .C(\datapath.registers.1226[27] [9]),
    .Y(_5625_)
);

OAI21X1 _16083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf0),
    .B(_5454__bF$buf0),
    .C(_5625_),
    .Y(_5044_)
);

OAI21X1 _16084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf7),
    .B(_5434__bF$buf1),
    .C(\datapath.registers.1226[27] [10]),
    .Y(_5626_)
);

OAI21X1 _16085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf4),
    .B(_5456__bF$buf0),
    .C(_5626_),
    .Y(_5014_)
);

OAI21X1 _16086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf6),
    .B(_5434__bF$buf0),
    .C(\datapath.registers.1226[27] [11]),
    .Y(_5627_)
);

OAI21X1 _16087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf3),
    .B(_5458__bF$buf0),
    .C(_5627_),
    .Y(_5015_)
);

OAI21X1 _16088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf5),
    .B(_5434__bF$buf14),
    .C(\datapath.registers.1226[27] [12]),
    .Y(_5628_)
);

OAI21X1 _16089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf2),
    .B(_5460__bF$buf0),
    .C(_5628_),
    .Y(_5016_)
);

OAI21X1 _16090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf4),
    .B(_5434__bF$buf13),
    .C(\datapath.registers.1226[27] [13]),
    .Y(_5629_)
);

OAI21X1 _16091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf1),
    .B(_5462__bF$buf0),
    .C(_5629_),
    .Y(_5017_)
);

OAI21X1 _16092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf3),
    .B(_5434__bF$buf12),
    .C(\datapath.registers.1226[27] [14]),
    .Y(_5630_)
);

OAI21X1 _16093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf0),
    .B(_5464__bF$buf0),
    .C(_5630_),
    .Y(_5018_)
);

OAI21X1 _16094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf2),
    .B(_5434__bF$buf11),
    .C(\datapath.registers.1226[27] [15]),
    .Y(_5631_)
);

OAI21X1 _16095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf4),
    .B(_5466__bF$buf0),
    .C(_5631_),
    .Y(_5019_)
);

OAI21X1 _16096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf1),
    .B(_5434__bF$buf10),
    .C(\datapath.registers.1226[27] [16]),
    .Y(_5632_)
);

OAI21X1 _16097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf3),
    .B(_5468__bF$buf0),
    .C(_5632_),
    .Y(_5020_)
);

OAI21X1 _16098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf0),
    .B(_5434__bF$buf9),
    .C(\datapath.registers.1226[27] [17]),
    .Y(_5633_)
);

OAI21X1 _16099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf2),
    .B(_5470__bF$buf0),
    .C(_5633_),
    .Y(_5021_)
);

OAI21X1 _16100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf8),
    .B(_5434__bF$buf8),
    .C(\datapath.registers.1226[27] [18]),
    .Y(_5634_)
);

OAI21X1 _16101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf1),
    .B(_5472__bF$buf0),
    .C(_5634_),
    .Y(_5022_)
);

OAI21X1 _16102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf7),
    .B(_5434__bF$buf7),
    .C(\datapath.registers.1226[27] [19]),
    .Y(_5635_)
);

OAI21X1 _16103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf0),
    .B(_5474__bF$buf0),
    .C(_5635_),
    .Y(_5023_)
);

OAI21X1 _16104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf6),
    .B(_5434__bF$buf6),
    .C(\datapath.registers.1226[27] [20]),
    .Y(_5636_)
);

OAI21X1 _16105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf4),
    .B(_5476__bF$buf0),
    .C(_5636_),
    .Y(_5025_)
);

OAI21X1 _16106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf5),
    .B(_5434__bF$buf5),
    .C(\datapath.registers.1226[27] [21]),
    .Y(_5637_)
);

OAI21X1 _16107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf3),
    .B(_5478__bF$buf0),
    .C(_5637_),
    .Y(_5026_)
);

OAI21X1 _16108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf4),
    .B(_5434__bF$buf4),
    .C(\datapath.registers.1226[27] [22]),
    .Y(_5638_)
);

OAI21X1 _16109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf2),
    .B(_5480__bF$buf0),
    .C(_5638_),
    .Y(_5027_)
);

OAI21X1 _16110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf3),
    .B(_5434__bF$buf3),
    .C(\datapath.registers.1226[27] [23]),
    .Y(_5639_)
);

OAI21X1 _16111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf1),
    .B(_5482__bF$buf0),
    .C(_5639_),
    .Y(_5028_)
);

OAI21X1 _16112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf2),
    .B(_5434__bF$buf2),
    .C(\datapath.registers.1226[27] [24]),
    .Y(_5640_)
);

OAI21X1 _16113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf0),
    .B(_5484__bF$buf0),
    .C(_5640_),
    .Y(_5029_)
);

OAI21X1 _16114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf1),
    .B(_5434__bF$buf1),
    .C(\datapath.registers.1226[27] [25]),
    .Y(_5641_)
);

OAI21X1 _16115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf4),
    .B(_5486__bF$buf0),
    .C(_5641_),
    .Y(_5030_)
);

OAI21X1 _16116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf0),
    .B(_5434__bF$buf0),
    .C(\datapath.registers.1226[27] [26]),
    .Y(_5642_)
);

OAI21X1 _16117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf3),
    .B(_5488__bF$buf0),
    .C(_5642_),
    .Y(_5031_)
);

OAI21X1 _16118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf8),
    .B(_5434__bF$buf14),
    .C(\datapath.registers.1226[27] [27]),
    .Y(_5643_)
);

OAI21X1 _16119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf2),
    .B(_5490__bF$buf0),
    .C(_5643_),
    .Y(_5032_)
);

OAI21X1 _16120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf7),
    .B(_5434__bF$buf13),
    .C(\datapath.registers.1226[27] [28]),
    .Y(_5644_)
);

OAI21X1 _16121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf1),
    .B(_5492__bF$buf0),
    .C(_5644_),
    .Y(_5033_)
);

OAI21X1 _16122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf6),
    .B(_5434__bF$buf12),
    .C(\datapath.registers.1226[27] [29]),
    .Y(_5645_)
);

OAI21X1 _16123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf0),
    .B(_5494__bF$buf0),
    .C(_5645_),
    .Y(_5034_)
);

OAI21X1 _16124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf5),
    .B(_5434__bF$buf11),
    .C(\datapath.registers.1226[27] [30]),
    .Y(_5646_)
);

OAI21X1 _16125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf4),
    .B(_5496__bF$buf0),
    .C(_5646_),
    .Y(_5036_)
);

OAI21X1 _16126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf4),
    .B(_5434__bF$buf10),
    .C(\datapath.registers.1226[27] [31]),
    .Y(_5647_)
);

OAI21X1 _16127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614__bF$buf3),
    .B(_5498__bF$buf0),
    .C(_5647_),
    .Y(_5037_)
);

NAND2X1 _16128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5613_),
    .B(_5508_),
    .Y(_5648_)
);

OAI21X1 _16129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf15),
    .B(_5615__bF$buf3),
    .C(\datapath.registers.1226[26] [0]),
    .Y(_5649_)
);

OAI21X1 _16130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf4),
    .B(_5648__bF$buf4),
    .C(_5649_),
    .Y(_4981_)
);

OAI21X1 _16131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf14),
    .B(_5615__bF$buf2),
    .C(\datapath.registers.1226[26] [1]),
    .Y(_5650_)
);

OAI21X1 _16132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf4),
    .B(_5648__bF$buf3),
    .C(_5650_),
    .Y(_4992_)
);

OAI21X1 _16133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf13),
    .B(_5615__bF$buf1),
    .C(\datapath.registers.1226[26] [2]),
    .Y(_5651_)
);

OAI21X1 _16134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf4),
    .B(_5648__bF$buf2),
    .C(_5651_),
    .Y(_5003_)
);

OAI21X1 _16135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf12),
    .B(_5615__bF$buf0),
    .C(\datapath.registers.1226[26] [3]),
    .Y(_5652_)
);

OAI21X1 _16136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf4),
    .B(_5648__bF$buf1),
    .C(_5652_),
    .Y(_5006_)
);

OAI21X1 _16137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf11),
    .B(_5615__bF$buf8),
    .C(\datapath.registers.1226[26] [4]),
    .Y(_5653_)
);

OAI21X1 _16138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf4),
    .B(_5648__bF$buf0),
    .C(_5653_),
    .Y(_5007_)
);

OAI21X1 _16139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf10),
    .B(_5615__bF$buf7),
    .C(\datapath.registers.1226[26] [5]),
    .Y(_5654_)
);

OAI21X1 _16140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf4),
    .B(_5648__bF$buf4),
    .C(_5654_),
    .Y(_5008_)
);

OAI21X1 _16141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf9),
    .B(_5615__bF$buf6),
    .C(\datapath.registers.1226[26] [6]),
    .Y(_5655_)
);

OAI21X1 _16142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf4),
    .B(_5648__bF$buf3),
    .C(_5655_),
    .Y(_5009_)
);

OAI21X1 _16143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf8),
    .B(_5615__bF$buf5),
    .C(\datapath.registers.1226[26] [7]),
    .Y(_5656_)
);

OAI21X1 _16144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf4),
    .B(_5648__bF$buf2),
    .C(_5656_),
    .Y(_5010_)
);

OAI21X1 _16145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf7),
    .B(_5615__bF$buf4),
    .C(\datapath.registers.1226[26] [8]),
    .Y(_5657_)
);

OAI21X1 _16146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf4),
    .B(_5648__bF$buf1),
    .C(_5657_),
    .Y(_5011_)
);

OAI21X1 _16147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf6),
    .B(_5615__bF$buf3),
    .C(\datapath.registers.1226[26] [9]),
    .Y(_5658_)
);

OAI21X1 _16148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf4),
    .B(_5648__bF$buf0),
    .C(_5658_),
    .Y(_5012_)
);

OAI21X1 _16149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf5),
    .B(_5615__bF$buf2),
    .C(\datapath.registers.1226[26] [10]),
    .Y(_5659_)
);

OAI21X1 _16150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf4),
    .B(_5648__bF$buf4),
    .C(_5659_),
    .Y(_4982_)
);

OAI21X1 _16151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf4),
    .B(_5615__bF$buf1),
    .C(\datapath.registers.1226[26] [11]),
    .Y(_5660_)
);

OAI21X1 _16152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf4),
    .B(_5648__bF$buf3),
    .C(_5660_),
    .Y(_4983_)
);

OAI21X1 _16153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf3),
    .B(_5615__bF$buf0),
    .C(\datapath.registers.1226[26] [12]),
    .Y(_5661_)
);

OAI21X1 _16154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf4),
    .B(_5648__bF$buf2),
    .C(_5661_),
    .Y(_4984_)
);

OAI21X1 _16155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf2),
    .B(_5615__bF$buf8),
    .C(\datapath.registers.1226[26] [13]),
    .Y(_5662_)
);

OAI21X1 _16156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf4),
    .B(_5648__bF$buf1),
    .C(_5662_),
    .Y(_4985_)
);

OAI21X1 _16157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf1),
    .B(_5615__bF$buf7),
    .C(\datapath.registers.1226[26] [14]),
    .Y(_5663_)
);

OAI21X1 _16158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf4),
    .B(_5648__bF$buf0),
    .C(_5663_),
    .Y(_4986_)
);

OAI21X1 _16159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf0),
    .B(_5615__bF$buf6),
    .C(\datapath.registers.1226[26] [15]),
    .Y(_5664_)
);

OAI21X1 _16160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf4),
    .B(_5648__bF$buf4),
    .C(_5664_),
    .Y(_4987_)
);

OAI21X1 _16161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf15),
    .B(_5615__bF$buf5),
    .C(\datapath.registers.1226[26] [16]),
    .Y(_5665_)
);

OAI21X1 _16162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf4),
    .B(_5648__bF$buf3),
    .C(_5665_),
    .Y(_4988_)
);

OAI21X1 _16163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf14),
    .B(_5615__bF$buf4),
    .C(\datapath.registers.1226[26] [17]),
    .Y(_5666_)
);

OAI21X1 _16164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf4),
    .B(_5648__bF$buf2),
    .C(_5666_),
    .Y(_4989_)
);

OAI21X1 _16165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf13),
    .B(_5615__bF$buf3),
    .C(\datapath.registers.1226[26] [18]),
    .Y(_5667_)
);

OAI21X1 _16166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf4),
    .B(_5648__bF$buf1),
    .C(_5667_),
    .Y(_4990_)
);

OAI21X1 _16167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf12),
    .B(_5615__bF$buf2),
    .C(\datapath.registers.1226[26] [19]),
    .Y(_5668_)
);

OAI21X1 _16168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf4),
    .B(_5648__bF$buf0),
    .C(_5668_),
    .Y(_4991_)
);

OAI21X1 _16169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf11),
    .B(_5615__bF$buf1),
    .C(\datapath.registers.1226[26] [20]),
    .Y(_5669_)
);

OAI21X1 _16170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf4),
    .B(_5648__bF$buf4),
    .C(_5669_),
    .Y(_4993_)
);

OAI21X1 _16171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf10),
    .B(_5615__bF$buf0),
    .C(\datapath.registers.1226[26] [21]),
    .Y(_5670_)
);

OAI21X1 _16172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf4),
    .B(_5648__bF$buf3),
    .C(_5670_),
    .Y(_4994_)
);

OAI21X1 _16173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf9),
    .B(_5615__bF$buf8),
    .C(\datapath.registers.1226[26] [22]),
    .Y(_5671_)
);

OAI21X1 _16174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf4),
    .B(_5648__bF$buf2),
    .C(_5671_),
    .Y(_4995_)
);

OAI21X1 _16175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf8),
    .B(_5615__bF$buf7),
    .C(\datapath.registers.1226[26] [23]),
    .Y(_5672_)
);

OAI21X1 _16176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf4),
    .B(_5648__bF$buf1),
    .C(_5672_),
    .Y(_4996_)
);

OAI21X1 _16177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf7),
    .B(_5615__bF$buf6),
    .C(\datapath.registers.1226[26] [24]),
    .Y(_5673_)
);

OAI21X1 _16178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf4),
    .B(_5648__bF$buf0),
    .C(_5673_),
    .Y(_4997_)
);

OAI21X1 _16179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf6),
    .B(_5615__bF$buf5),
    .C(\datapath.registers.1226[26] [25]),
    .Y(_5674_)
);

OAI21X1 _16180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486__bF$buf4),
    .B(_5648__bF$buf4),
    .C(_5674_),
    .Y(_4998_)
);

OAI21X1 _16181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf5),
    .B(_5615__bF$buf4),
    .C(\datapath.registers.1226[26] [26]),
    .Y(_5675_)
);

OAI21X1 _16182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf4),
    .B(_5648__bF$buf3),
    .C(_5675_),
    .Y(_4999_)
);

OAI21X1 _16183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf4),
    .B(_5615__bF$buf3),
    .C(\datapath.registers.1226[26] [27]),
    .Y(_5676_)
);

OAI21X1 _16184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf4),
    .B(_5648__bF$buf2),
    .C(_5676_),
    .Y(_5000_)
);

OAI21X1 _16185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf3),
    .B(_5615__bF$buf2),
    .C(\datapath.registers.1226[26] [28]),
    .Y(_5677_)
);

OAI21X1 _16186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf4),
    .B(_5648__bF$buf1),
    .C(_5677_),
    .Y(_5001_)
);

OAI21X1 _16187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf2),
    .B(_5615__bF$buf1),
    .C(\datapath.registers.1226[26] [29]),
    .Y(_5678_)
);

OAI21X1 _16188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf4),
    .B(_5648__bF$buf0),
    .C(_5678_),
    .Y(_5002_)
);

OAI21X1 _16189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf1),
    .B(_5615__bF$buf0),
    .C(\datapath.registers.1226[26] [30]),
    .Y(_5679_)
);

OAI21X1 _16190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf4),
    .B(_5648__bF$buf4),
    .C(_5679_),
    .Y(_5004_)
);

OAI21X1 _16191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf0),
    .B(_5615__bF$buf8),
    .C(\datapath.registers.1226[26] [31]),
    .Y(_5680_)
);

OAI21X1 _16192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf4),
    .B(_5648__bF$buf3),
    .C(_5680_),
    .Y(_5005_)
);

NAND2X1 _16193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5613_),
    .B(_5544_),
    .Y(_5681_)
);

OAI21X1 _16194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf15),
    .B(_5615__bF$buf7),
    .C(\datapath.registers.1226[25] [0]),
    .Y(_5682_)
);

OAI21X1 _16195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf3),
    .B(_5681__bF$buf4),
    .C(_5682_),
    .Y(_4949_)
);

OAI21X1 _16196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf14),
    .B(_5615__bF$buf6),
    .C(\datapath.registers.1226[25] [1]),
    .Y(_5683_)
);

OAI21X1 _16197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf3),
    .B(_5681__bF$buf3),
    .C(_5683_),
    .Y(_4960_)
);

OAI21X1 _16198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf13),
    .B(_5615__bF$buf5),
    .C(\datapath.registers.1226[25] [2]),
    .Y(_5684_)
);

OAI21X1 _16199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf3),
    .B(_5681__bF$buf2),
    .C(_5684_),
    .Y(_4971_)
);

OAI21X1 _16200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf12),
    .B(_5615__bF$buf4),
    .C(\datapath.registers.1226[25] [3]),
    .Y(_5685_)
);

OAI21X1 _16201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf3),
    .B(_5681__bF$buf1),
    .C(_5685_),
    .Y(_4974_)
);

OAI21X1 _16202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf11),
    .B(_5615__bF$buf3),
    .C(\datapath.registers.1226[25] [4]),
    .Y(_5686_)
);

OAI21X1 _16203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf3),
    .B(_5681__bF$buf0),
    .C(_5686_),
    .Y(_4975_)
);

OAI21X1 _16204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf10),
    .B(_5615__bF$buf2),
    .C(\datapath.registers.1226[25] [5]),
    .Y(_5687_)
);

OAI21X1 _16205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf3),
    .B(_5681__bF$buf4),
    .C(_5687_),
    .Y(_4976_)
);

OAI21X1 _16206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf9),
    .B(_5615__bF$buf1),
    .C(\datapath.registers.1226[25] [6]),
    .Y(_5688_)
);

OAI21X1 _16207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf3),
    .B(_5681__bF$buf3),
    .C(_5688_),
    .Y(_4977_)
);

OAI21X1 _16208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf8),
    .B(_5615__bF$buf0),
    .C(\datapath.registers.1226[25] [7]),
    .Y(_5689_)
);

OAI21X1 _16209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf3),
    .B(_5681__bF$buf2),
    .C(_5689_),
    .Y(_4978_)
);

OAI21X1 _16210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf7),
    .B(_5615__bF$buf8),
    .C(\datapath.registers.1226[25] [8]),
    .Y(_5690_)
);

OAI21X1 _16211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf3),
    .B(_5681__bF$buf1),
    .C(_5690_),
    .Y(_4979_)
);

OAI21X1 _16212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf6),
    .B(_5615__bF$buf7),
    .C(\datapath.registers.1226[25] [9]),
    .Y(_5691_)
);

OAI21X1 _16213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf3),
    .B(_5681__bF$buf0),
    .C(_5691_),
    .Y(_4980_)
);

OAI21X1 _16214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf5),
    .B(_5615__bF$buf6),
    .C(\datapath.registers.1226[25] [10]),
    .Y(_5692_)
);

OAI21X1 _16215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf3),
    .B(_5681__bF$buf4),
    .C(_5692_),
    .Y(_4950_)
);

OAI21X1 _16216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf4),
    .B(_5615__bF$buf5),
    .C(\datapath.registers.1226[25] [11]),
    .Y(_5693_)
);

OAI21X1 _16217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf3),
    .B(_5681__bF$buf3),
    .C(_5693_),
    .Y(_4951_)
);

OAI21X1 _16218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf3),
    .B(_5615__bF$buf4),
    .C(\datapath.registers.1226[25] [12]),
    .Y(_5694_)
);

OAI21X1 _16219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf3),
    .B(_5681__bF$buf2),
    .C(_5694_),
    .Y(_4952_)
);

OAI21X1 _16220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf2),
    .B(_5615__bF$buf3),
    .C(\datapath.registers.1226[25] [13]),
    .Y(_5695_)
);

OAI21X1 _16221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf3),
    .B(_5681__bF$buf1),
    .C(_5695_),
    .Y(_4953_)
);

OAI21X1 _16222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf1),
    .B(_5615__bF$buf2),
    .C(\datapath.registers.1226[25] [14]),
    .Y(_5696_)
);

OAI21X1 _16223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf3),
    .B(_5681__bF$buf0),
    .C(_5696_),
    .Y(_4954_)
);

OAI21X1 _16224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf0),
    .B(_5615__bF$buf1),
    .C(\datapath.registers.1226[25] [15]),
    .Y(_5697_)
);

OAI21X1 _16225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf3),
    .B(_5681__bF$buf4),
    .C(_5697_),
    .Y(_4955_)
);

OAI21X1 _16226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf15),
    .B(_5615__bF$buf0),
    .C(\datapath.registers.1226[25] [16]),
    .Y(_5698_)
);

OAI21X1 _16227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf3),
    .B(_5681__bF$buf3),
    .C(_5698_),
    .Y(_4956_)
);

OAI21X1 _16228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf14),
    .B(_5615__bF$buf8),
    .C(\datapath.registers.1226[25] [17]),
    .Y(_5699_)
);

OAI21X1 _16229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf3),
    .B(_5681__bF$buf2),
    .C(_5699_),
    .Y(_4957_)
);

OAI21X1 _16230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf13),
    .B(_5615__bF$buf7),
    .C(\datapath.registers.1226[25] [18]),
    .Y(_5700_)
);

OAI21X1 _16231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf3),
    .B(_5681__bF$buf1),
    .C(_5700_),
    .Y(_4958_)
);

OAI21X1 _16232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf12),
    .B(_5615__bF$buf6),
    .C(\datapath.registers.1226[25] [19]),
    .Y(_5701_)
);

OAI21X1 _16233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf3),
    .B(_5681__bF$buf0),
    .C(_5701_),
    .Y(_4959_)
);

OAI21X1 _16234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf11),
    .B(_5615__bF$buf5),
    .C(\datapath.registers.1226[25] [20]),
    .Y(_5702_)
);

OAI21X1 _16235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf3),
    .B(_5681__bF$buf4),
    .C(_5702_),
    .Y(_4961_)
);

OAI21X1 _16236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf10),
    .B(_5615__bF$buf4),
    .C(\datapath.registers.1226[25] [21]),
    .Y(_5703_)
);

OAI21X1 _16237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf3),
    .B(_5681__bF$buf3),
    .C(_5703_),
    .Y(_4962_)
);

OAI21X1 _16238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf9),
    .B(_5615__bF$buf3),
    .C(\datapath.registers.1226[25] [22]),
    .Y(_5704_)
);

OAI21X1 _16239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf3),
    .B(_5681__bF$buf2),
    .C(_5704_),
    .Y(_4963_)
);

OAI21X1 _16240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf8),
    .B(_5615__bF$buf2),
    .C(\datapath.registers.1226[25] [23]),
    .Y(_5705_)
);

OAI21X1 _16241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf3),
    .B(_5681__bF$buf1),
    .C(_5705_),
    .Y(_4964_)
);

OAI21X1 _16242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf7),
    .B(_5615__bF$buf1),
    .C(\datapath.registers.1226[25] [24]),
    .Y(_5706_)
);

OAI21X1 _16243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf3),
    .B(_5681__bF$buf0),
    .C(_5706_),
    .Y(_4965_)
);

OAI21X1 _16244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf6),
    .B(_5615__bF$buf0),
    .C(\datapath.registers.1226[25] [25]),
    .Y(_5707_)
);

OAI21X1 _16245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486__bF$buf3),
    .B(_5681__bF$buf4),
    .C(_5707_),
    .Y(_4966_)
);

OAI21X1 _16246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf5),
    .B(_5615__bF$buf8),
    .C(\datapath.registers.1226[25] [26]),
    .Y(_5708_)
);

OAI21X1 _16247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf3),
    .B(_5681__bF$buf3),
    .C(_5708_),
    .Y(_4967_)
);

OAI21X1 _16248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf4),
    .B(_5615__bF$buf7),
    .C(\datapath.registers.1226[25] [27]),
    .Y(_5709_)
);

OAI21X1 _16249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf3),
    .B(_5681__bF$buf2),
    .C(_5709_),
    .Y(_4968_)
);

OAI21X1 _16250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf3),
    .B(_5615__bF$buf6),
    .C(\datapath.registers.1226[25] [28]),
    .Y(_5710_)
);

OAI21X1 _16251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf3),
    .B(_5681__bF$buf1),
    .C(_5710_),
    .Y(_4969_)
);

OAI21X1 _16252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf2),
    .B(_5615__bF$buf5),
    .C(\datapath.registers.1226[25] [29]),
    .Y(_5711_)
);

OAI21X1 _16253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf3),
    .B(_5681__bF$buf0),
    .C(_5711_),
    .Y(_4970_)
);

OAI21X1 _16254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf1),
    .B(_5615__bF$buf4),
    .C(\datapath.registers.1226[25] [30]),
    .Y(_5712_)
);

OAI21X1 _16255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf3),
    .B(_5681__bF$buf4),
    .C(_5712_),
    .Y(_4972_)
);

OAI21X1 _16256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf0),
    .B(_5615__bF$buf3),
    .C(\datapath.registers.1226[25] [31]),
    .Y(_5713_)
);

OAI21X1 _16257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf3),
    .B(_5681__bF$buf3),
    .C(_5713_),
    .Y(_4973_)
);

INVX1 _16258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [0]),
    .Y(_5714_)
);

NOR2X1 _16259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5615__bF$buf2),
    .B(_5579__bF$buf2),
    .Y(_5715_)
);

NAND2X1 _16260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [0]),
    .B(_5715__bF$buf7),
    .Y(_5716_)
);

OAI21X1 _16261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5714_),
    .B(_5715__bF$buf6),
    .C(_5716_),
    .Y(_4917_)
);

NOR2X1 _16262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [1]),
    .B(_5715__bF$buf5),
    .Y(_5717_)
);

AOI21X1 _16263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf2),
    .B(_5715__bF$buf4),
    .C(_5717_),
    .Y(_4928_)
);

NOR2X1 _16264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [2]),
    .B(_5715__bF$buf3),
    .Y(_5718_)
);

AOI21X1 _16265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf2),
    .B(_5715__bF$buf2),
    .C(_5718_),
    .Y(_4939_)
);

INVX1 _16266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [3]),
    .Y(_5719_)
);

NAND2X1 _16267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [3]),
    .B(_5715__bF$buf1),
    .Y(_5720_)
);

OAI21X1 _16268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5719_),
    .B(_5715__bF$buf0),
    .C(_5720_),
    .Y(_4942_)
);

NOR2X1 _16269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [4]),
    .B(_5715__bF$buf7),
    .Y(_5721_)
);

AOI21X1 _16270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf2),
    .B(_5715__bF$buf6),
    .C(_5721_),
    .Y(_4943_)
);

NOR2X1 _16271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [5]),
    .B(_5715__bF$buf5),
    .Y(_5722_)
);

AOI21X1 _16272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf2),
    .B(_5715__bF$buf4),
    .C(_5722_),
    .Y(_4944_)
);

NOR2X1 _16273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [6]),
    .B(_5715__bF$buf3),
    .Y(_5723_)
);

AOI21X1 _16274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf2),
    .B(_5715__bF$buf2),
    .C(_5723_),
    .Y(_4945_)
);

NOR2X1 _16275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [7]),
    .B(_5715__bF$buf1),
    .Y(_5724_)
);

AOI21X1 _16276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf2),
    .B(_5715__bF$buf0),
    .C(_5724_),
    .Y(_4946_)
);

NOR2X1 _16277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [8]),
    .B(_5715__bF$buf7),
    .Y(_5725_)
);

AOI21X1 _16278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf2),
    .B(_5715__bF$buf6),
    .C(_5725_),
    .Y(_4947_)
);

NOR2X1 _16279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [9]),
    .B(_5715__bF$buf5),
    .Y(_5726_)
);

AOI21X1 _16280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf2),
    .B(_5715__bF$buf4),
    .C(_5726_),
    .Y(_4948_)
);

INVX1 _16281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [10]),
    .Y(_5727_)
);

NAND2X1 _16282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [10]),
    .B(_5715__bF$buf3),
    .Y(_5728_)
);

OAI21X1 _16283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5727_),
    .B(_5715__bF$buf2),
    .C(_5728_),
    .Y(_4918_)
);

NOR2X1 _16284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [11]),
    .B(_5715__bF$buf1),
    .Y(_5729_)
);

AOI21X1 _16285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf2),
    .B(_5715__bF$buf0),
    .C(_5729_),
    .Y(_4919_)
);

NOR2X1 _16286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [12]),
    .B(_5715__bF$buf7),
    .Y(_5730_)
);

AOI21X1 _16287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf2),
    .B(_5715__bF$buf6),
    .C(_5730_),
    .Y(_4920_)
);

NOR2X1 _16288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [13]),
    .B(_5715__bF$buf5),
    .Y(_5731_)
);

AOI21X1 _16289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf2),
    .B(_5715__bF$buf4),
    .C(_5731_),
    .Y(_4921_)
);

NOR2X1 _16290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [14]),
    .B(_5715__bF$buf3),
    .Y(_5732_)
);

AOI21X1 _16291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf2),
    .B(_5715__bF$buf2),
    .C(_5732_),
    .Y(_4922_)
);

NOR2X1 _16292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [15]),
    .B(_5715__bF$buf1),
    .Y(_5733_)
);

AOI21X1 _16293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf2),
    .B(_5715__bF$buf0),
    .C(_5733_),
    .Y(_4923_)
);

INVX1 _16294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [16]),
    .Y(_5734_)
);

NAND2X1 _16295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [16]),
    .B(_5715__bF$buf7),
    .Y(_5735_)
);

OAI21X1 _16296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5734_),
    .B(_5715__bF$buf6),
    .C(_5735_),
    .Y(_4924_)
);

INVX1 _16297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [17]),
    .Y(_5736_)
);

NAND2X1 _16298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [17]),
    .B(_5715__bF$buf5),
    .Y(_5737_)
);

OAI21X1 _16299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5736_),
    .B(_5715__bF$buf4),
    .C(_5737_),
    .Y(_4925_)
);

NOR2X1 _16300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [18]),
    .B(_5715__bF$buf3),
    .Y(_5738_)
);

AOI21X1 _16301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf2),
    .B(_5715__bF$buf2),
    .C(_5738_),
    .Y(_4926_)
);

NOR2X1 _16302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [19]),
    .B(_5715__bF$buf1),
    .Y(_5739_)
);

AOI21X1 _16303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf2),
    .B(_5715__bF$buf0),
    .C(_5739_),
    .Y(_4927_)
);

INVX1 _16304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [20]),
    .Y(_5740_)
);

NAND2X1 _16305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [20]),
    .B(_5715__bF$buf7),
    .Y(_5741_)
);

OAI21X1 _16306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5740_),
    .B(_5715__bF$buf6),
    .C(_5741_),
    .Y(_4929_)
);

INVX1 _16307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [21]),
    .Y(_5742_)
);

NAND2X1 _16308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [21]),
    .B(_5715__bF$buf5),
    .Y(_5743_)
);

OAI21X1 _16309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5742_),
    .B(_5715__bF$buf4),
    .C(_5743_),
    .Y(_4930_)
);

NOR2X1 _16310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [22]),
    .B(_5715__bF$buf3),
    .Y(_5744_)
);

AOI21X1 _16311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf2),
    .B(_5715__bF$buf2),
    .C(_5744_),
    .Y(_4931_)
);

NOR2X1 _16312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [23]),
    .B(_5715__bF$buf1),
    .Y(_5745_)
);

AOI21X1 _16313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf2),
    .B(_5715__bF$buf0),
    .C(_5745_),
    .Y(_4932_)
);

NOR2X1 _16314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [24]),
    .B(_5715__bF$buf7),
    .Y(_5746_)
);

AOI21X1 _16315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf2),
    .B(_5715__bF$buf6),
    .C(_5746_),
    .Y(_4933_)
);

INVX1 _16316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [25]),
    .Y(_5747_)
);

NAND2X1 _16317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [25]),
    .B(_5715__bF$buf5),
    .Y(_5748_)
);

OAI21X1 _16318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5747_),
    .B(_5715__bF$buf4),
    .C(_5748_),
    .Y(_4934_)
);

NOR2X1 _16319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [26]),
    .B(_5715__bF$buf3),
    .Y(_5749_)
);

AOI21X1 _16320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf2),
    .B(_5715__bF$buf2),
    .C(_5749_),
    .Y(_4935_)
);

NOR2X1 _16321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [27]),
    .B(_5715__bF$buf1),
    .Y(_5750_)
);

AOI21X1 _16322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf2),
    .B(_5715__bF$buf0),
    .C(_5750_),
    .Y(_4936_)
);

INVX1 _16323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [28]),
    .Y(_5751_)
);

NAND2X1 _16324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [28]),
    .B(_5715__bF$buf7),
    .Y(_5752_)
);

OAI21X1 _16325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5751_),
    .B(_5715__bF$buf6),
    .C(_5752_),
    .Y(_4937_)
);

NOR2X1 _16326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [29]),
    .B(_5715__bF$buf5),
    .Y(_5753_)
);

AOI21X1 _16327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf2),
    .B(_5715__bF$buf4),
    .C(_5753_),
    .Y(_4938_)
);

NOR2X1 _16328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [30]),
    .B(_5715__bF$buf3),
    .Y(_5754_)
);

AOI21X1 _16329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf2),
    .B(_5715__bF$buf2),
    .C(_5754_),
    .Y(_4940_)
);

INVX1 _16330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[24] [31]),
    .Y(_5755_)
);

NAND2X1 _16331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [31]),
    .B(_5715__bF$buf1),
    .Y(_5756_)
);

OAI21X1 _16332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5755_),
    .B(_5715__bF$buf0),
    .C(_5756_),
    .Y(_4941_)
);

NAND2X1 _16333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [11]),
    .B(_5504_),
    .Y(_5757_)
);

NOR2X1 _16334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5430_),
    .B(_5757_),
    .Y(_5758_)
);

NAND2X1 _16335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5435_),
    .B(_5758_),
    .Y(_5759_)
);

INVX8 _16336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5758_),
    .Y(_5760_)
);

OAI21X1 _16337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf8),
    .B(_5434__bF$buf9),
    .C(\datapath.registers.1226[23] [0]),
    .Y(_5761_)
);

OAI21X1 _16338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf4),
    .B(_5429__bF$buf2),
    .C(_5761_),
    .Y(_4885_)
);

OAI21X1 _16339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf7),
    .B(_5434__bF$buf8),
    .C(\datapath.registers.1226[23] [1]),
    .Y(_5762_)
);

OAI21X1 _16340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf3),
    .B(_5438__bF$buf1),
    .C(_5762_),
    .Y(_4896_)
);

OAI21X1 _16341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf6),
    .B(_5434__bF$buf7),
    .C(\datapath.registers.1226[23] [2]),
    .Y(_5763_)
);

OAI21X1 _16342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf2),
    .B(_5440__bF$buf1),
    .C(_5763_),
    .Y(_4907_)
);

OAI21X1 _16343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf5),
    .B(_5434__bF$buf6),
    .C(\datapath.registers.1226[23] [3]),
    .Y(_5764_)
);

OAI21X1 _16344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf1),
    .B(_5442__bF$buf2),
    .C(_5764_),
    .Y(_4910_)
);

OAI21X1 _16345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf4),
    .B(_5434__bF$buf5),
    .C(\datapath.registers.1226[23] [4]),
    .Y(_5765_)
);

OAI21X1 _16346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf0),
    .B(_5444__bF$buf1),
    .C(_5765_),
    .Y(_4911_)
);

OAI21X1 _16347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf3),
    .B(_5434__bF$buf4),
    .C(\datapath.registers.1226[23] [5]),
    .Y(_5766_)
);

OAI21X1 _16348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf4),
    .B(_5446__bF$buf1),
    .C(_5766_),
    .Y(_4912_)
);

OAI21X1 _16349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf2),
    .B(_5434__bF$buf3),
    .C(\datapath.registers.1226[23] [6]),
    .Y(_5767_)
);

OAI21X1 _16350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf3),
    .B(_5448__bF$buf1),
    .C(_5767_),
    .Y(_4913_)
);

OAI21X1 _16351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf1),
    .B(_5434__bF$buf2),
    .C(\datapath.registers.1226[23] [7]),
    .Y(_5768_)
);

OAI21X1 _16352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf2),
    .B(_5450__bF$buf1),
    .C(_5768_),
    .Y(_4914_)
);

OAI21X1 _16353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf0),
    .B(_5434__bF$buf1),
    .C(\datapath.registers.1226[23] [8]),
    .Y(_5769_)
);

OAI21X1 _16354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf1),
    .B(_5452__bF$buf1),
    .C(_5769_),
    .Y(_4915_)
);

OAI21X1 _16355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf8),
    .B(_5434__bF$buf0),
    .C(\datapath.registers.1226[23] [9]),
    .Y(_5770_)
);

OAI21X1 _16356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf0),
    .B(_5454__bF$buf1),
    .C(_5770_),
    .Y(_4916_)
);

OAI21X1 _16357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf7),
    .B(_5434__bF$buf14),
    .C(\datapath.registers.1226[23] [10]),
    .Y(_5771_)
);

OAI21X1 _16358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf4),
    .B(_5456__bF$buf2),
    .C(_5771_),
    .Y(_4886_)
);

OAI21X1 _16359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf6),
    .B(_5434__bF$buf13),
    .C(\datapath.registers.1226[23] [11]),
    .Y(_5772_)
);

OAI21X1 _16360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf3),
    .B(_5458__bF$buf1),
    .C(_5772_),
    .Y(_4887_)
);

OAI21X1 _16361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf5),
    .B(_5434__bF$buf12),
    .C(\datapath.registers.1226[23] [12]),
    .Y(_5773_)
);

OAI21X1 _16362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf2),
    .B(_5460__bF$buf1),
    .C(_5773_),
    .Y(_4888_)
);

OAI21X1 _16363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf4),
    .B(_5434__bF$buf11),
    .C(\datapath.registers.1226[23] [13]),
    .Y(_5774_)
);

OAI21X1 _16364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf1),
    .B(_5462__bF$buf1),
    .C(_5774_),
    .Y(_4889_)
);

OAI21X1 _16365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf3),
    .B(_5434__bF$buf10),
    .C(\datapath.registers.1226[23] [14]),
    .Y(_5775_)
);

OAI21X1 _16366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf0),
    .B(_5464__bF$buf1),
    .C(_5775_),
    .Y(_4890_)
);

OAI21X1 _16367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf2),
    .B(_5434__bF$buf9),
    .C(\datapath.registers.1226[23] [15]),
    .Y(_5776_)
);

OAI21X1 _16368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf4),
    .B(_5466__bF$buf1),
    .C(_5776_),
    .Y(_4891_)
);

OAI21X1 _16369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf1),
    .B(_5434__bF$buf8),
    .C(\datapath.registers.1226[23] [16]),
    .Y(_5777_)
);

OAI21X1 _16370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf3),
    .B(_5468__bF$buf2),
    .C(_5777_),
    .Y(_4892_)
);

OAI21X1 _16371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf0),
    .B(_5434__bF$buf7),
    .C(\datapath.registers.1226[23] [17]),
    .Y(_5778_)
);

OAI21X1 _16372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf2),
    .B(_5470__bF$buf2),
    .C(_5778_),
    .Y(_4893_)
);

OAI21X1 _16373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf8),
    .B(_5434__bF$buf6),
    .C(\datapath.registers.1226[23] [18]),
    .Y(_5779_)
);

OAI21X1 _16374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf1),
    .B(_5472__bF$buf1),
    .C(_5779_),
    .Y(_4894_)
);

OAI21X1 _16375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf7),
    .B(_5434__bF$buf5),
    .C(\datapath.registers.1226[23] [19]),
    .Y(_5780_)
);

OAI21X1 _16376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf0),
    .B(_5474__bF$buf1),
    .C(_5780_),
    .Y(_4895_)
);

OAI21X1 _16377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf6),
    .B(_5434__bF$buf4),
    .C(\datapath.registers.1226[23] [20]),
    .Y(_5781_)
);

OAI21X1 _16378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf4),
    .B(_5476__bF$buf2),
    .C(_5781_),
    .Y(_4897_)
);

OAI21X1 _16379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf5),
    .B(_5434__bF$buf3),
    .C(\datapath.registers.1226[23] [21]),
    .Y(_5782_)
);

OAI21X1 _16380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf3),
    .B(_5478__bF$buf2),
    .C(_5782_),
    .Y(_4898_)
);

OAI21X1 _16381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf4),
    .B(_5434__bF$buf2),
    .C(\datapath.registers.1226[23] [22]),
    .Y(_5783_)
);

OAI21X1 _16382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf2),
    .B(_5480__bF$buf1),
    .C(_5783_),
    .Y(_4899_)
);

OAI21X1 _16383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf3),
    .B(_5434__bF$buf1),
    .C(\datapath.registers.1226[23] [23]),
    .Y(_5784_)
);

OAI21X1 _16384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf1),
    .B(_5482__bF$buf1),
    .C(_5784_),
    .Y(_4900_)
);

OAI21X1 _16385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf2),
    .B(_5434__bF$buf0),
    .C(\datapath.registers.1226[23] [24]),
    .Y(_5785_)
);

OAI21X1 _16386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf0),
    .B(_5484__bF$buf1),
    .C(_5785_),
    .Y(_4901_)
);

OAI21X1 _16387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf1),
    .B(_5434__bF$buf14),
    .C(\datapath.registers.1226[23] [25]),
    .Y(_5786_)
);

OAI21X1 _16388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf4),
    .B(_5486__bF$buf2),
    .C(_5786_),
    .Y(_4902_)
);

OAI21X1 _16389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf0),
    .B(_5434__bF$buf13),
    .C(\datapath.registers.1226[23] [26]),
    .Y(_5787_)
);

OAI21X1 _16390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf3),
    .B(_5488__bF$buf1),
    .C(_5787_),
    .Y(_4903_)
);

OAI21X1 _16391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf8),
    .B(_5434__bF$buf12),
    .C(\datapath.registers.1226[23] [27]),
    .Y(_5788_)
);

OAI21X1 _16392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf2),
    .B(_5490__bF$buf1),
    .C(_5788_),
    .Y(_4904_)
);

OAI21X1 _16393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf7),
    .B(_5434__bF$buf11),
    .C(\datapath.registers.1226[23] [28]),
    .Y(_5789_)
);

OAI21X1 _16394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf1),
    .B(_5492__bF$buf2),
    .C(_5789_),
    .Y(_4905_)
);

OAI21X1 _16395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf6),
    .B(_5434__bF$buf10),
    .C(\datapath.registers.1226[23] [29]),
    .Y(_5790_)
);

OAI21X1 _16396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf0),
    .B(_5494__bF$buf1),
    .C(_5790_),
    .Y(_4906_)
);

OAI21X1 _16397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf5),
    .B(_5434__bF$buf9),
    .C(\datapath.registers.1226[23] [30]),
    .Y(_5791_)
);

OAI21X1 _16398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf4),
    .B(_5496__bF$buf1),
    .C(_5791_),
    .Y(_4908_)
);

OAI21X1 _16399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5760__bF$buf4),
    .B(_5434__bF$buf8),
    .C(\datapath.registers.1226[23] [31]),
    .Y(_5792_)
);

OAI21X1 _16400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759__bF$buf3),
    .B(_5498__bF$buf2),
    .C(_5792_),
    .Y(_4909_)
);

NAND2X1 _16401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5758_),
    .B(_5508_),
    .Y(_5793_)
);

OAI21X1 _16402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf15),
    .B(_5760__bF$buf3),
    .C(\datapath.registers.1226[22] [0]),
    .Y(_5794_)
);

OAI21X1 _16403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf1),
    .B(_5793__bF$buf4),
    .C(_5794_),
    .Y(_4853_)
);

OAI21X1 _16404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf14),
    .B(_5760__bF$buf2),
    .C(\datapath.registers.1226[22] [1]),
    .Y(_5795_)
);

OAI21X1 _16405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf0),
    .B(_5793__bF$buf3),
    .C(_5795_),
    .Y(_4864_)
);

OAI21X1 _16406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf13),
    .B(_5760__bF$buf1),
    .C(\datapath.registers.1226[22] [2]),
    .Y(_5796_)
);

OAI21X1 _16407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf0),
    .B(_5793__bF$buf2),
    .C(_5796_),
    .Y(_4875_)
);

OAI21X1 _16408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf12),
    .B(_5760__bF$buf0),
    .C(\datapath.registers.1226[22] [3]),
    .Y(_5797_)
);

OAI21X1 _16409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf1),
    .B(_5793__bF$buf1),
    .C(_5797_),
    .Y(_4878_)
);

OAI21X1 _16410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf11),
    .B(_5760__bF$buf8),
    .C(\datapath.registers.1226[22] [4]),
    .Y(_5798_)
);

OAI21X1 _16411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf0),
    .B(_5793__bF$buf0),
    .C(_5798_),
    .Y(_4879_)
);

OAI21X1 _16412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf10),
    .B(_5760__bF$buf7),
    .C(\datapath.registers.1226[22] [5]),
    .Y(_5799_)
);

OAI21X1 _16413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf0),
    .B(_5793__bF$buf4),
    .C(_5799_),
    .Y(_4880_)
);

OAI21X1 _16414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf9),
    .B(_5760__bF$buf6),
    .C(\datapath.registers.1226[22] [6]),
    .Y(_5800_)
);

OAI21X1 _16415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf0),
    .B(_5793__bF$buf3),
    .C(_5800_),
    .Y(_4881_)
);

OAI21X1 _16416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf8),
    .B(_5760__bF$buf5),
    .C(\datapath.registers.1226[22] [7]),
    .Y(_5801_)
);

OAI21X1 _16417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf0),
    .B(_5793__bF$buf2),
    .C(_5801_),
    .Y(_4882_)
);

OAI21X1 _16418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf7),
    .B(_5760__bF$buf4),
    .C(\datapath.registers.1226[22] [8]),
    .Y(_5802_)
);

OAI21X1 _16419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf0),
    .B(_5793__bF$buf1),
    .C(_5802_),
    .Y(_4883_)
);

OAI21X1 _16420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf6),
    .B(_5760__bF$buf3),
    .C(\datapath.registers.1226[22] [9]),
    .Y(_5803_)
);

OAI21X1 _16421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf0),
    .B(_5793__bF$buf0),
    .C(_5803_),
    .Y(_4884_)
);

OAI21X1 _16422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf5),
    .B(_5760__bF$buf2),
    .C(\datapath.registers.1226[22] [10]),
    .Y(_5804_)
);

OAI21X1 _16423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf1),
    .B(_5793__bF$buf4),
    .C(_5804_),
    .Y(_4854_)
);

OAI21X1 _16424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf4),
    .B(_5760__bF$buf1),
    .C(\datapath.registers.1226[22] [11]),
    .Y(_5805_)
);

OAI21X1 _16425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf0),
    .B(_5793__bF$buf3),
    .C(_5805_),
    .Y(_4855_)
);

OAI21X1 _16426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf3),
    .B(_5760__bF$buf0),
    .C(\datapath.registers.1226[22] [12]),
    .Y(_5806_)
);

OAI21X1 _16427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf0),
    .B(_5793__bF$buf2),
    .C(_5806_),
    .Y(_4856_)
);

OAI21X1 _16428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf2),
    .B(_5760__bF$buf8),
    .C(\datapath.registers.1226[22] [13]),
    .Y(_5807_)
);

OAI21X1 _16429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf0),
    .B(_5793__bF$buf1),
    .C(_5807_),
    .Y(_4857_)
);

OAI21X1 _16430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf1),
    .B(_5760__bF$buf7),
    .C(\datapath.registers.1226[22] [14]),
    .Y(_5808_)
);

OAI21X1 _16431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf0),
    .B(_5793__bF$buf0),
    .C(_5808_),
    .Y(_4858_)
);

OAI21X1 _16432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf0),
    .B(_5760__bF$buf6),
    .C(\datapath.registers.1226[22] [15]),
    .Y(_5809_)
);

OAI21X1 _16433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf0),
    .B(_5793__bF$buf4),
    .C(_5809_),
    .Y(_4859_)
);

OAI21X1 _16434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf15),
    .B(_5760__bF$buf5),
    .C(\datapath.registers.1226[22] [16]),
    .Y(_5810_)
);

OAI21X1 _16435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf1),
    .B(_5793__bF$buf3),
    .C(_5810_),
    .Y(_4860_)
);

OAI21X1 _16436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf14),
    .B(_5760__bF$buf4),
    .C(\datapath.registers.1226[22] [17]),
    .Y(_5811_)
);

OAI21X1 _16437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf1),
    .B(_5793__bF$buf2),
    .C(_5811_),
    .Y(_4861_)
);

OAI21X1 _16438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf13),
    .B(_5760__bF$buf3),
    .C(\datapath.registers.1226[22] [18]),
    .Y(_5812_)
);

OAI21X1 _16439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf0),
    .B(_5793__bF$buf1),
    .C(_5812_),
    .Y(_4862_)
);

OAI21X1 _16440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf12),
    .B(_5760__bF$buf2),
    .C(\datapath.registers.1226[22] [19]),
    .Y(_5813_)
);

OAI21X1 _16441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf0),
    .B(_5793__bF$buf0),
    .C(_5813_),
    .Y(_4863_)
);

OAI21X1 _16442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf11),
    .B(_5760__bF$buf1),
    .C(\datapath.registers.1226[22] [20]),
    .Y(_5814_)
);

OAI21X1 _16443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf1),
    .B(_5793__bF$buf4),
    .C(_5814_),
    .Y(_4865_)
);

OAI21X1 _16444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf10),
    .B(_5760__bF$buf0),
    .C(\datapath.registers.1226[22] [21]),
    .Y(_5815_)
);

OAI21X1 _16445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf1),
    .B(_5793__bF$buf3),
    .C(_5815_),
    .Y(_4866_)
);

OAI21X1 _16446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf9),
    .B(_5760__bF$buf8),
    .C(\datapath.registers.1226[22] [22]),
    .Y(_5816_)
);

OAI21X1 _16447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf0),
    .B(_5793__bF$buf2),
    .C(_5816_),
    .Y(_4867_)
);

OAI21X1 _16448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf8),
    .B(_5760__bF$buf7),
    .C(\datapath.registers.1226[22] [23]),
    .Y(_5817_)
);

OAI21X1 _16449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf0),
    .B(_5793__bF$buf1),
    .C(_5817_),
    .Y(_4868_)
);

OAI21X1 _16450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf7),
    .B(_5760__bF$buf6),
    .C(\datapath.registers.1226[22] [24]),
    .Y(_5818_)
);

OAI21X1 _16451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf0),
    .B(_5793__bF$buf0),
    .C(_5818_),
    .Y(_4869_)
);

OAI21X1 _16452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf6),
    .B(_5760__bF$buf5),
    .C(\datapath.registers.1226[22] [25]),
    .Y(_5819_)
);

OAI21X1 _16453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486__bF$buf1),
    .B(_5793__bF$buf4),
    .C(_5819_),
    .Y(_4870_)
);

OAI21X1 _16454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf5),
    .B(_5760__bF$buf4),
    .C(\datapath.registers.1226[22] [26]),
    .Y(_5820_)
);

OAI21X1 _16455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf0),
    .B(_5793__bF$buf3),
    .C(_5820_),
    .Y(_4871_)
);

OAI21X1 _16456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf4),
    .B(_5760__bF$buf3),
    .C(\datapath.registers.1226[22] [27]),
    .Y(_5821_)
);

OAI21X1 _16457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf0),
    .B(_5793__bF$buf2),
    .C(_5821_),
    .Y(_4872_)
);

OAI21X1 _16458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf3),
    .B(_5760__bF$buf2),
    .C(\datapath.registers.1226[22] [28]),
    .Y(_5822_)
);

OAI21X1 _16459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf1),
    .B(_5793__bF$buf1),
    .C(_5822_),
    .Y(_4873_)
);

OAI21X1 _16460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf2),
    .B(_5760__bF$buf1),
    .C(\datapath.registers.1226[22] [29]),
    .Y(_5823_)
);

OAI21X1 _16461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf0),
    .B(_5793__bF$buf0),
    .C(_5823_),
    .Y(_4874_)
);

OAI21X1 _16462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf1),
    .B(_5760__bF$buf0),
    .C(\datapath.registers.1226[22] [30]),
    .Y(_5824_)
);

OAI21X1 _16463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf0),
    .B(_5793__bF$buf4),
    .C(_5824_),
    .Y(_4876_)
);

OAI21X1 _16464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf0),
    .B(_5760__bF$buf8),
    .C(\datapath.registers.1226[22] [31]),
    .Y(_5825_)
);

OAI21X1 _16465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf1),
    .B(_5793__bF$buf3),
    .C(_5825_),
    .Y(_4877_)
);

NAND2X1 _16466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5758_),
    .B(_5544_),
    .Y(_5826_)
);

OAI21X1 _16467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf15),
    .B(_5760__bF$buf7),
    .C(\datapath.registers.1226[21] [0]),
    .Y(_5827_)
);

OAI21X1 _16468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf0),
    .B(_5826__bF$buf4),
    .C(_5827_),
    .Y(_4821_)
);

OAI21X1 _16469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf14),
    .B(_5760__bF$buf6),
    .C(\datapath.registers.1226[21] [1]),
    .Y(_5828_)
);

OAI21X1 _16470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf4),
    .B(_5826__bF$buf3),
    .C(_5828_),
    .Y(_4832_)
);

OAI21X1 _16471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf13),
    .B(_5760__bF$buf5),
    .C(\datapath.registers.1226[21] [2]),
    .Y(_5829_)
);

OAI21X1 _16472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf4),
    .B(_5826__bF$buf2),
    .C(_5829_),
    .Y(_4843_)
);

OAI21X1 _16473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf12),
    .B(_5760__bF$buf4),
    .C(\datapath.registers.1226[21] [3]),
    .Y(_5830_)
);

OAI21X1 _16474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf0),
    .B(_5826__bF$buf1),
    .C(_5830_),
    .Y(_4846_)
);

OAI21X1 _16475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf11),
    .B(_5760__bF$buf3),
    .C(\datapath.registers.1226[21] [4]),
    .Y(_5831_)
);

OAI21X1 _16476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf4),
    .B(_5826__bF$buf0),
    .C(_5831_),
    .Y(_4847_)
);

OAI21X1 _16477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf10),
    .B(_5760__bF$buf2),
    .C(\datapath.registers.1226[21] [5]),
    .Y(_5832_)
);

OAI21X1 _16478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf4),
    .B(_5826__bF$buf4),
    .C(_5832_),
    .Y(_4848_)
);

OAI21X1 _16479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf9),
    .B(_5760__bF$buf1),
    .C(\datapath.registers.1226[21] [6]),
    .Y(_5833_)
);

OAI21X1 _16480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf4),
    .B(_5826__bF$buf3),
    .C(_5833_),
    .Y(_4849_)
);

OAI21X1 _16481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf8),
    .B(_5760__bF$buf0),
    .C(\datapath.registers.1226[21] [7]),
    .Y(_5834_)
);

OAI21X1 _16482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf4),
    .B(_5826__bF$buf2),
    .C(_5834_),
    .Y(_4850_)
);

OAI21X1 _16483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf7),
    .B(_5760__bF$buf8),
    .C(\datapath.registers.1226[21] [8]),
    .Y(_5835_)
);

OAI21X1 _16484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf4),
    .B(_5826__bF$buf1),
    .C(_5835_),
    .Y(_4851_)
);

OAI21X1 _16485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf6),
    .B(_5760__bF$buf7),
    .C(\datapath.registers.1226[21] [9]),
    .Y(_5836_)
);

OAI21X1 _16486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf4),
    .B(_5826__bF$buf0),
    .C(_5836_),
    .Y(_4852_)
);

OAI21X1 _16487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf5),
    .B(_5760__bF$buf6),
    .C(\datapath.registers.1226[21] [10]),
    .Y(_5837_)
);

OAI21X1 _16488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf0),
    .B(_5826__bF$buf4),
    .C(_5837_),
    .Y(_4822_)
);

OAI21X1 _16489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf4),
    .B(_5760__bF$buf5),
    .C(\datapath.registers.1226[21] [11]),
    .Y(_5838_)
);

OAI21X1 _16490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf4),
    .B(_5826__bF$buf3),
    .C(_5838_),
    .Y(_4823_)
);

OAI21X1 _16491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf3),
    .B(_5760__bF$buf4),
    .C(\datapath.registers.1226[21] [12]),
    .Y(_5839_)
);

OAI21X1 _16492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf4),
    .B(_5826__bF$buf2),
    .C(_5839_),
    .Y(_4824_)
);

OAI21X1 _16493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf2),
    .B(_5760__bF$buf3),
    .C(\datapath.registers.1226[21] [13]),
    .Y(_5840_)
);

OAI21X1 _16494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf4),
    .B(_5826__bF$buf1),
    .C(_5840_),
    .Y(_4825_)
);

OAI21X1 _16495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf1),
    .B(_5760__bF$buf2),
    .C(\datapath.registers.1226[21] [14]),
    .Y(_5841_)
);

OAI21X1 _16496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf4),
    .B(_5826__bF$buf0),
    .C(_5841_),
    .Y(_4826_)
);

OAI21X1 _16497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf0),
    .B(_5760__bF$buf1),
    .C(\datapath.registers.1226[21] [15]),
    .Y(_5842_)
);

OAI21X1 _16498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf4),
    .B(_5826__bF$buf4),
    .C(_5842_),
    .Y(_4827_)
);

OAI21X1 _16499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf15),
    .B(_5760__bF$buf0),
    .C(\datapath.registers.1226[21] [16]),
    .Y(_5843_)
);

OAI21X1 _16500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf0),
    .B(_5826__bF$buf3),
    .C(_5843_),
    .Y(_4828_)
);

OAI21X1 _16501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf14),
    .B(_5760__bF$buf8),
    .C(\datapath.registers.1226[21] [17]),
    .Y(_5844_)
);

OAI21X1 _16502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf0),
    .B(_5826__bF$buf2),
    .C(_5844_),
    .Y(_4829_)
);

OAI21X1 _16503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf13),
    .B(_5760__bF$buf7),
    .C(\datapath.registers.1226[21] [18]),
    .Y(_5845_)
);

OAI21X1 _16504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf4),
    .B(_5826__bF$buf1),
    .C(_5845_),
    .Y(_4830_)
);

OAI21X1 _16505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf12),
    .B(_5760__bF$buf6),
    .C(\datapath.registers.1226[21] [19]),
    .Y(_5846_)
);

OAI21X1 _16506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf4),
    .B(_5826__bF$buf0),
    .C(_5846_),
    .Y(_4831_)
);

OAI21X1 _16507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf11),
    .B(_5760__bF$buf5),
    .C(\datapath.registers.1226[21] [20]),
    .Y(_5847_)
);

OAI21X1 _16508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf0),
    .B(_5826__bF$buf4),
    .C(_5847_),
    .Y(_4833_)
);

OAI21X1 _16509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf10),
    .B(_5760__bF$buf4),
    .C(\datapath.registers.1226[21] [21]),
    .Y(_5848_)
);

OAI21X1 _16510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf0),
    .B(_5826__bF$buf3),
    .C(_5848_),
    .Y(_4834_)
);

OAI21X1 _16511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf9),
    .B(_5760__bF$buf3),
    .C(\datapath.registers.1226[21] [22]),
    .Y(_5849_)
);

OAI21X1 _16512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf4),
    .B(_5826__bF$buf2),
    .C(_5849_),
    .Y(_4835_)
);

OAI21X1 _16513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf8),
    .B(_5760__bF$buf2),
    .C(\datapath.registers.1226[21] [23]),
    .Y(_5850_)
);

OAI21X1 _16514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf4),
    .B(_5826__bF$buf1),
    .C(_5850_),
    .Y(_4836_)
);

OAI21X1 _16515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf7),
    .B(_5760__bF$buf1),
    .C(\datapath.registers.1226[21] [24]),
    .Y(_5851_)
);

OAI21X1 _16516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf4),
    .B(_5826__bF$buf0),
    .C(_5851_),
    .Y(_4837_)
);

OAI21X1 _16517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf6),
    .B(_5760__bF$buf0),
    .C(\datapath.registers.1226[21] [25]),
    .Y(_5852_)
);

OAI21X1 _16518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486__bF$buf0),
    .B(_5826__bF$buf4),
    .C(_5852_),
    .Y(_4838_)
);

OAI21X1 _16519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf5),
    .B(_5760__bF$buf8),
    .C(\datapath.registers.1226[21] [26]),
    .Y(_5853_)
);

OAI21X1 _16520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf4),
    .B(_5826__bF$buf3),
    .C(_5853_),
    .Y(_4839_)
);

OAI21X1 _16521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf4),
    .B(_5760__bF$buf7),
    .C(\datapath.registers.1226[21] [27]),
    .Y(_5854_)
);

OAI21X1 _16522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf4),
    .B(_5826__bF$buf2),
    .C(_5854_),
    .Y(_4840_)
);

OAI21X1 _16523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf3),
    .B(_5760__bF$buf6),
    .C(\datapath.registers.1226[21] [28]),
    .Y(_5855_)
);

OAI21X1 _16524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf0),
    .B(_5826__bF$buf1),
    .C(_5855_),
    .Y(_4841_)
);

OAI21X1 _16525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf2),
    .B(_5760__bF$buf5),
    .C(\datapath.registers.1226[21] [29]),
    .Y(_5856_)
);

OAI21X1 _16526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf4),
    .B(_5826__bF$buf0),
    .C(_5856_),
    .Y(_4842_)
);

OAI21X1 _16527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf1),
    .B(_5760__bF$buf4),
    .C(\datapath.registers.1226[21] [30]),
    .Y(_5857_)
);

OAI21X1 _16528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf4),
    .B(_5826__bF$buf4),
    .C(_5857_),
    .Y(_4844_)
);

OAI21X1 _16529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf0),
    .B(_5760__bF$buf3),
    .C(\datapath.registers.1226[21] [31]),
    .Y(_5858_)
);

OAI21X1 _16530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf0),
    .B(_5826__bF$buf3),
    .C(_5858_),
    .Y(_4845_)
);

NOR2X1 _16531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf1),
    .B(_5760__bF$buf2),
    .Y(_5859_)
);

NOR2X1 _16532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [0]),
    .B(_5859__bF$buf7),
    .Y(_5860_)
);

AOI21X1 _16533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf4),
    .B(_5859__bF$buf6),
    .C(_5860_),
    .Y(_4789_)
);

NOR2X1 _16534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [1]),
    .B(_5859__bF$buf5),
    .Y(_5861_)
);

AOI21X1 _16535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf3),
    .B(_5859__bF$buf4),
    .C(_5861_),
    .Y(_4800_)
);

NOR2X1 _16536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [2]),
    .B(_5859__bF$buf3),
    .Y(_5862_)
);

AOI21X1 _16537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf3),
    .B(_5859__bF$buf2),
    .C(_5862_),
    .Y(_4811_)
);

NOR2X1 _16538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [3]),
    .B(_5859__bF$buf1),
    .Y(_5863_)
);

AOI21X1 _16539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf4),
    .B(_5859__bF$buf0),
    .C(_5863_),
    .Y(_4814_)
);

NOR2X1 _16540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [4]),
    .B(_5859__bF$buf7),
    .Y(_5864_)
);

AOI21X1 _16541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf3),
    .B(_5859__bF$buf6),
    .C(_5864_),
    .Y(_4815_)
);

NOR2X1 _16542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [5]),
    .B(_5859__bF$buf5),
    .Y(_5865_)
);

AOI21X1 _16543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf3),
    .B(_5859__bF$buf4),
    .C(_5865_),
    .Y(_4816_)
);

NOR2X1 _16544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [6]),
    .B(_5859__bF$buf3),
    .Y(_5866_)
);

AOI21X1 _16545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf3),
    .B(_5859__bF$buf2),
    .C(_5866_),
    .Y(_4817_)
);

NOR2X1 _16546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [7]),
    .B(_5859__bF$buf1),
    .Y(_5867_)
);

AOI21X1 _16547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf3),
    .B(_5859__bF$buf0),
    .C(_5867_),
    .Y(_4818_)
);

NOR2X1 _16548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [8]),
    .B(_5859__bF$buf7),
    .Y(_5868_)
);

AOI21X1 _16549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf3),
    .B(_5859__bF$buf6),
    .C(_5868_),
    .Y(_4819_)
);

NOR2X1 _16550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [9]),
    .B(_5859__bF$buf5),
    .Y(_5869_)
);

AOI21X1 _16551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf3),
    .B(_5859__bF$buf4),
    .C(_5869_),
    .Y(_4820_)
);

NOR2X1 _16552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [10]),
    .B(_5859__bF$buf3),
    .Y(_5870_)
);

AOI21X1 _16553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf4),
    .B(_5859__bF$buf2),
    .C(_5870_),
    .Y(_4790_)
);

NOR2X1 _16554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [11]),
    .B(_5859__bF$buf1),
    .Y(_5871_)
);

AOI21X1 _16555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf3),
    .B(_5859__bF$buf0),
    .C(_5871_),
    .Y(_4791_)
);

NOR2X1 _16556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [12]),
    .B(_5859__bF$buf7),
    .Y(_5872_)
);

AOI21X1 _16557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf3),
    .B(_5859__bF$buf6),
    .C(_5872_),
    .Y(_4792_)
);

NOR2X1 _16558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [13]),
    .B(_5859__bF$buf5),
    .Y(_5873_)
);

AOI21X1 _16559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf3),
    .B(_5859__bF$buf4),
    .C(_5873_),
    .Y(_4793_)
);

NOR2X1 _16560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [14]),
    .B(_5859__bF$buf3),
    .Y(_5874_)
);

AOI21X1 _16561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf3),
    .B(_5859__bF$buf2),
    .C(_5874_),
    .Y(_4794_)
);

NOR2X1 _16562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [15]),
    .B(_5859__bF$buf1),
    .Y(_5875_)
);

AOI21X1 _16563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf3),
    .B(_5859__bF$buf0),
    .C(_5875_),
    .Y(_4795_)
);

NOR2X1 _16564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [16]),
    .B(_5859__bF$buf7),
    .Y(_5876_)
);

AOI21X1 _16565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf4),
    .B(_5859__bF$buf6),
    .C(_5876_),
    .Y(_4796_)
);

NOR2X1 _16566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [17]),
    .B(_5859__bF$buf5),
    .Y(_5877_)
);

AOI21X1 _16567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf4),
    .B(_5859__bF$buf4),
    .C(_5877_),
    .Y(_4797_)
);

NOR2X1 _16568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [18]),
    .B(_5859__bF$buf3),
    .Y(_5878_)
);

AOI21X1 _16569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf3),
    .B(_5859__bF$buf2),
    .C(_5878_),
    .Y(_4798_)
);

NOR2X1 _16570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [19]),
    .B(_5859__bF$buf1),
    .Y(_5879_)
);

AOI21X1 _16571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf3),
    .B(_5859__bF$buf0),
    .C(_5879_),
    .Y(_4799_)
);

NOR2X1 _16572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [20]),
    .B(_5859__bF$buf7),
    .Y(_5880_)
);

AOI21X1 _16573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf4),
    .B(_5859__bF$buf6),
    .C(_5880_),
    .Y(_4801_)
);

NOR2X1 _16574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [21]),
    .B(_5859__bF$buf5),
    .Y(_5881_)
);

AOI21X1 _16575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf4),
    .B(_5859__bF$buf4),
    .C(_5881_),
    .Y(_4802_)
);

NOR2X1 _16576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [22]),
    .B(_5859__bF$buf3),
    .Y(_5882_)
);

AOI21X1 _16577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf3),
    .B(_5859__bF$buf2),
    .C(_5882_),
    .Y(_4803_)
);

NOR2X1 _16578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [23]),
    .B(_5859__bF$buf1),
    .Y(_5883_)
);

AOI21X1 _16579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf3),
    .B(_5859__bF$buf0),
    .C(_5883_),
    .Y(_4804_)
);

NOR2X1 _16580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [24]),
    .B(_5859__bF$buf7),
    .Y(_5884_)
);

AOI21X1 _16581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf3),
    .B(_5859__bF$buf6),
    .C(_5884_),
    .Y(_4805_)
);

NOR2X1 _16582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [25]),
    .B(_5859__bF$buf5),
    .Y(_5885_)
);

AOI21X1 _16583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486__bF$buf4),
    .B(_5859__bF$buf4),
    .C(_5885_),
    .Y(_4806_)
);

NOR2X1 _16584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [26]),
    .B(_5859__bF$buf3),
    .Y(_5886_)
);

AOI21X1 _16585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf3),
    .B(_5859__bF$buf2),
    .C(_5886_),
    .Y(_4807_)
);

NOR2X1 _16586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [27]),
    .B(_5859__bF$buf1),
    .Y(_5887_)
);

AOI21X1 _16587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf3),
    .B(_5859__bF$buf0),
    .C(_5887_),
    .Y(_4808_)
);

NOR2X1 _16588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [28]),
    .B(_5859__bF$buf7),
    .Y(_5888_)
);

AOI21X1 _16589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf4),
    .B(_5859__bF$buf6),
    .C(_5888_),
    .Y(_4809_)
);

NOR2X1 _16590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [29]),
    .B(_5859__bF$buf5),
    .Y(_5889_)
);

AOI21X1 _16591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf3),
    .B(_5859__bF$buf4),
    .C(_5889_),
    .Y(_4810_)
);

NOR2X1 _16592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [30]),
    .B(_5859__bF$buf3),
    .Y(_5890_)
);

AOI21X1 _16593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf3),
    .B(_5859__bF$buf2),
    .C(_5890_),
    .Y(_4812_)
);

NOR2X1 _16594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [31]),
    .B(_5859__bF$buf1),
    .Y(_5891_)
);

AOI21X1 _16595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf4),
    .B(_5859__bF$buf0),
    .C(_5891_),
    .Y(_4813_)
);

NOR2X1 _16596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [9]),
    .B(_5757_),
    .Y(_5892_)
);

NAND2X1 _16597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5435_),
    .B(_5892_),
    .Y(_5893_)
);

INVX8 _16598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5892_),
    .Y(_5894_)
);

OAI21X1 _16599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf8),
    .B(_5434__bF$buf7),
    .C(\datapath.registers.1226[19] [0]),
    .Y(_5895_)
);

OAI21X1 _16600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf4),
    .B(_5429__bF$buf3),
    .C(_5895_),
    .Y(_4725_)
);

OAI21X1 _16601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf7),
    .B(_5434__bF$buf6),
    .C(\datapath.registers.1226[19] [1]),
    .Y(_5896_)
);

OAI21X1 _16602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf3),
    .B(_5438__bF$buf2),
    .C(_5896_),
    .Y(_4736_)
);

OAI21X1 _16603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf6),
    .B(_5434__bF$buf5),
    .C(\datapath.registers.1226[19] [2]),
    .Y(_5897_)
);

OAI21X1 _16604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf2),
    .B(_5440__bF$buf2),
    .C(_5897_),
    .Y(_4747_)
);

OAI21X1 _16605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf5),
    .B(_5434__bF$buf4),
    .C(\datapath.registers.1226[19] [3]),
    .Y(_5898_)
);

OAI21X1 _16606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf1),
    .B(_5442__bF$buf3),
    .C(_5898_),
    .Y(_4750_)
);

OAI21X1 _16607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf4),
    .B(_5434__bF$buf3),
    .C(\datapath.registers.1226[19] [4]),
    .Y(_5899_)
);

OAI21X1 _16608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf0),
    .B(_5444__bF$buf2),
    .C(_5899_),
    .Y(_4751_)
);

OAI21X1 _16609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf3),
    .B(_5434__bF$buf2),
    .C(\datapath.registers.1226[19] [5]),
    .Y(_5900_)
);

OAI21X1 _16610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf4),
    .B(_5446__bF$buf2),
    .C(_5900_),
    .Y(_4752_)
);

OAI21X1 _16611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf2),
    .B(_5434__bF$buf1),
    .C(\datapath.registers.1226[19] [6]),
    .Y(_5901_)
);

OAI21X1 _16612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf3),
    .B(_5448__bF$buf2),
    .C(_5901_),
    .Y(_4753_)
);

OAI21X1 _16613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf1),
    .B(_5434__bF$buf0),
    .C(\datapath.registers.1226[19] [7]),
    .Y(_5902_)
);

OAI21X1 _16614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf2),
    .B(_5450__bF$buf2),
    .C(_5902_),
    .Y(_4754_)
);

OAI21X1 _16615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf0),
    .B(_5434__bF$buf14),
    .C(\datapath.registers.1226[19] [8]),
    .Y(_5903_)
);

OAI21X1 _16616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf1),
    .B(_5452__bF$buf2),
    .C(_5903_),
    .Y(_4755_)
);

OAI21X1 _16617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf8),
    .B(_5434__bF$buf13),
    .C(\datapath.registers.1226[19] [9]),
    .Y(_5904_)
);

OAI21X1 _16618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf0),
    .B(_5454__bF$buf2),
    .C(_5904_),
    .Y(_4756_)
);

OAI21X1 _16619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf7),
    .B(_5434__bF$buf12),
    .C(\datapath.registers.1226[19] [10]),
    .Y(_5905_)
);

OAI21X1 _16620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf4),
    .B(_5456__bF$buf3),
    .C(_5905_),
    .Y(_4726_)
);

OAI21X1 _16621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf6),
    .B(_5434__bF$buf11),
    .C(\datapath.registers.1226[19] [11]),
    .Y(_5906_)
);

OAI21X1 _16622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf3),
    .B(_5458__bF$buf2),
    .C(_5906_),
    .Y(_4727_)
);

OAI21X1 _16623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf5),
    .B(_5434__bF$buf10),
    .C(\datapath.registers.1226[19] [12]),
    .Y(_5907_)
);

OAI21X1 _16624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf2),
    .B(_5460__bF$buf2),
    .C(_5907_),
    .Y(_4728_)
);

OAI21X1 _16625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf4),
    .B(_5434__bF$buf9),
    .C(\datapath.registers.1226[19] [13]),
    .Y(_5908_)
);

OAI21X1 _16626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf1),
    .B(_5462__bF$buf2),
    .C(_5908_),
    .Y(_4729_)
);

OAI21X1 _16627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf3),
    .B(_5434__bF$buf8),
    .C(\datapath.registers.1226[19] [14]),
    .Y(_5909_)
);

OAI21X1 _16628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf0),
    .B(_5464__bF$buf2),
    .C(_5909_),
    .Y(_4730_)
);

OAI21X1 _16629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf2),
    .B(_5434__bF$buf7),
    .C(\datapath.registers.1226[19] [15]),
    .Y(_5910_)
);

OAI21X1 _16630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf4),
    .B(_5466__bF$buf2),
    .C(_5910_),
    .Y(_4731_)
);

OAI21X1 _16631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf1),
    .B(_5434__bF$buf6),
    .C(\datapath.registers.1226[19] [16]),
    .Y(_5911_)
);

OAI21X1 _16632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf3),
    .B(_5468__bF$buf3),
    .C(_5911_),
    .Y(_4732_)
);

OAI21X1 _16633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf0),
    .B(_5434__bF$buf5),
    .C(\datapath.registers.1226[19] [17]),
    .Y(_5912_)
);

OAI21X1 _16634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf2),
    .B(_5470__bF$buf3),
    .C(_5912_),
    .Y(_4733_)
);

OAI21X1 _16635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf8),
    .B(_5434__bF$buf4),
    .C(\datapath.registers.1226[19] [18]),
    .Y(_5913_)
);

OAI21X1 _16636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf1),
    .B(_5472__bF$buf2),
    .C(_5913_),
    .Y(_4734_)
);

OAI21X1 _16637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf7),
    .B(_5434__bF$buf3),
    .C(\datapath.registers.1226[19] [19]),
    .Y(_5914_)
);

OAI21X1 _16638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf0),
    .B(_5474__bF$buf2),
    .C(_5914_),
    .Y(_4735_)
);

OAI21X1 _16639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf6),
    .B(_5434__bF$buf2),
    .C(\datapath.registers.1226[19] [20]),
    .Y(_5915_)
);

OAI21X1 _16640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf4),
    .B(_5476__bF$buf3),
    .C(_5915_),
    .Y(_4737_)
);

OAI21X1 _16641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf5),
    .B(_5434__bF$buf1),
    .C(\datapath.registers.1226[19] [21]),
    .Y(_5916_)
);

OAI21X1 _16642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf3),
    .B(_5478__bF$buf3),
    .C(_5916_),
    .Y(_4738_)
);

OAI21X1 _16643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf4),
    .B(_5434__bF$buf0),
    .C(\datapath.registers.1226[19] [22]),
    .Y(_5917_)
);

OAI21X1 _16644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf2),
    .B(_5480__bF$buf2),
    .C(_5917_),
    .Y(_4739_)
);

OAI21X1 _16645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf3),
    .B(_5434__bF$buf14),
    .C(\datapath.registers.1226[19] [23]),
    .Y(_5918_)
);

OAI21X1 _16646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf1),
    .B(_5482__bF$buf2),
    .C(_5918_),
    .Y(_4740_)
);

OAI21X1 _16647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf2),
    .B(_5434__bF$buf13),
    .C(\datapath.registers.1226[19] [24]),
    .Y(_5919_)
);

OAI21X1 _16648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf0),
    .B(_5484__bF$buf2),
    .C(_5919_),
    .Y(_4741_)
);

OAI21X1 _16649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf1),
    .B(_5434__bF$buf12),
    .C(\datapath.registers.1226[19] [25]),
    .Y(_5920_)
);

OAI21X1 _16650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf4),
    .B(_5486__bF$buf3),
    .C(_5920_),
    .Y(_4742_)
);

OAI21X1 _16651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf0),
    .B(_5434__bF$buf11),
    .C(\datapath.registers.1226[19] [26]),
    .Y(_5921_)
);

OAI21X1 _16652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf3),
    .B(_5488__bF$buf2),
    .C(_5921_),
    .Y(_4743_)
);

OAI21X1 _16653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf8),
    .B(_5434__bF$buf10),
    .C(\datapath.registers.1226[19] [27]),
    .Y(_5922_)
);

OAI21X1 _16654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf2),
    .B(_5490__bF$buf2),
    .C(_5922_),
    .Y(_4744_)
);

OAI21X1 _16655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf7),
    .B(_5434__bF$buf9),
    .C(\datapath.registers.1226[19] [28]),
    .Y(_5923_)
);

OAI21X1 _16656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf1),
    .B(_5492__bF$buf3),
    .C(_5923_),
    .Y(_4745_)
);

OAI21X1 _16657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf6),
    .B(_5434__bF$buf8),
    .C(\datapath.registers.1226[19] [29]),
    .Y(_5924_)
);

OAI21X1 _16658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf0),
    .B(_5494__bF$buf2),
    .C(_5924_),
    .Y(_4746_)
);

OAI21X1 _16659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf5),
    .B(_5434__bF$buf7),
    .C(\datapath.registers.1226[19] [30]),
    .Y(_5925_)
);

OAI21X1 _16660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf4),
    .B(_5496__bF$buf2),
    .C(_5925_),
    .Y(_4748_)
);

OAI21X1 _16661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5894__bF$buf4),
    .B(_5434__bF$buf6),
    .C(\datapath.registers.1226[19] [31]),
    .Y(_5926_)
);

OAI21X1 _16662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893__bF$buf3),
    .B(_5498__bF$buf3),
    .C(_5926_),
    .Y(_4749_)
);

NAND2X1 _16663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5892_),
    .B(_5508_),
    .Y(_5927_)
);

OAI21X1 _16664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf15),
    .B(_5894__bF$buf3),
    .C(\datapath.registers.1226[18] [0]),
    .Y(_5928_)
);

OAI21X1 _16665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf2),
    .B(_5927__bF$buf4),
    .C(_5928_),
    .Y(_4693_)
);

OAI21X1 _16666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf14),
    .B(_5894__bF$buf2),
    .C(\datapath.registers.1226[18] [1]),
    .Y(_5929_)
);

OAI21X1 _16667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf1),
    .B(_5927__bF$buf3),
    .C(_5929_),
    .Y(_4704_)
);

OAI21X1 _16668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf13),
    .B(_5894__bF$buf1),
    .C(\datapath.registers.1226[18] [2]),
    .Y(_5930_)
);

OAI21X1 _16669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf1),
    .B(_5927__bF$buf2),
    .C(_5930_),
    .Y(_4715_)
);

OAI21X1 _16670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf12),
    .B(_5894__bF$buf0),
    .C(\datapath.registers.1226[18] [3]),
    .Y(_5931_)
);

OAI21X1 _16671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf2),
    .B(_5927__bF$buf1),
    .C(_5931_),
    .Y(_4718_)
);

OAI21X1 _16672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf11),
    .B(_5894__bF$buf8),
    .C(\datapath.registers.1226[18] [4]),
    .Y(_5932_)
);

OAI21X1 _16673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf1),
    .B(_5927__bF$buf0),
    .C(_5932_),
    .Y(_4719_)
);

OAI21X1 _16674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf10),
    .B(_5894__bF$buf7),
    .C(\datapath.registers.1226[18] [5]),
    .Y(_5933_)
);

OAI21X1 _16675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf1),
    .B(_5927__bF$buf4),
    .C(_5933_),
    .Y(_4720_)
);

OAI21X1 _16676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf9),
    .B(_5894__bF$buf6),
    .C(\datapath.registers.1226[18] [6]),
    .Y(_5934_)
);

OAI21X1 _16677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf1),
    .B(_5927__bF$buf3),
    .C(_5934_),
    .Y(_4721_)
);

OAI21X1 _16678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf8),
    .B(_5894__bF$buf5),
    .C(\datapath.registers.1226[18] [7]),
    .Y(_5935_)
);

OAI21X1 _16679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf1),
    .B(_5927__bF$buf2),
    .C(_5935_),
    .Y(_4722_)
);

OAI21X1 _16680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf7),
    .B(_5894__bF$buf4),
    .C(\datapath.registers.1226[18] [8]),
    .Y(_5936_)
);

OAI21X1 _16681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf1),
    .B(_5927__bF$buf1),
    .C(_5936_),
    .Y(_4723_)
);

OAI21X1 _16682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf6),
    .B(_5894__bF$buf3),
    .C(\datapath.registers.1226[18] [9]),
    .Y(_5937_)
);

OAI21X1 _16683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf1),
    .B(_5927__bF$buf0),
    .C(_5937_),
    .Y(_4724_)
);

OAI21X1 _16684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf5),
    .B(_5894__bF$buf2),
    .C(\datapath.registers.1226[18] [10]),
    .Y(_5938_)
);

OAI21X1 _16685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf2),
    .B(_5927__bF$buf4),
    .C(_5938_),
    .Y(_4694_)
);

OAI21X1 _16686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf4),
    .B(_5894__bF$buf1),
    .C(\datapath.registers.1226[18] [11]),
    .Y(_5939_)
);

OAI21X1 _16687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf1),
    .B(_5927__bF$buf3),
    .C(_5939_),
    .Y(_4695_)
);

OAI21X1 _16688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf3),
    .B(_5894__bF$buf0),
    .C(\datapath.registers.1226[18] [12]),
    .Y(_5940_)
);

OAI21X1 _16689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf1),
    .B(_5927__bF$buf2),
    .C(_5940_),
    .Y(_4696_)
);

OAI21X1 _16690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf2),
    .B(_5894__bF$buf8),
    .C(\datapath.registers.1226[18] [13]),
    .Y(_5941_)
);

OAI21X1 _16691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf1),
    .B(_5927__bF$buf1),
    .C(_5941_),
    .Y(_4697_)
);

OAI21X1 _16692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf1),
    .B(_5894__bF$buf7),
    .C(\datapath.registers.1226[18] [14]),
    .Y(_5942_)
);

OAI21X1 _16693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf1),
    .B(_5927__bF$buf0),
    .C(_5942_),
    .Y(_4698_)
);

OAI21X1 _16694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf0),
    .B(_5894__bF$buf6),
    .C(\datapath.registers.1226[18] [15]),
    .Y(_5943_)
);

OAI21X1 _16695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf1),
    .B(_5927__bF$buf4),
    .C(_5943_),
    .Y(_4699_)
);

OAI21X1 _16696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf15),
    .B(_5894__bF$buf5),
    .C(\datapath.registers.1226[18] [16]),
    .Y(_5944_)
);

OAI21X1 _16697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf2),
    .B(_5927__bF$buf3),
    .C(_5944_),
    .Y(_4700_)
);

OAI21X1 _16698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf14),
    .B(_5894__bF$buf4),
    .C(\datapath.registers.1226[18] [17]),
    .Y(_5945_)
);

OAI21X1 _16699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf2),
    .B(_5927__bF$buf2),
    .C(_5945_),
    .Y(_4701_)
);

OAI21X1 _16700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf13),
    .B(_5894__bF$buf3),
    .C(\datapath.registers.1226[18] [18]),
    .Y(_5946_)
);

OAI21X1 _16701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf1),
    .B(_5927__bF$buf1),
    .C(_5946_),
    .Y(_4702_)
);

OAI21X1 _16702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf12),
    .B(_5894__bF$buf2),
    .C(\datapath.registers.1226[18] [19]),
    .Y(_5947_)
);

OAI21X1 _16703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf1),
    .B(_5927__bF$buf0),
    .C(_5947_),
    .Y(_4703_)
);

OAI21X1 _16704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf11),
    .B(_5894__bF$buf1),
    .C(\datapath.registers.1226[18] [20]),
    .Y(_5948_)
);

OAI21X1 _16705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf2),
    .B(_5927__bF$buf4),
    .C(_5948_),
    .Y(_4705_)
);

OAI21X1 _16706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf10),
    .B(_5894__bF$buf0),
    .C(\datapath.registers.1226[18] [21]),
    .Y(_5949_)
);

OAI21X1 _16707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf2),
    .B(_5927__bF$buf3),
    .C(_5949_),
    .Y(_4706_)
);

OAI21X1 _16708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf9),
    .B(_5894__bF$buf8),
    .C(\datapath.registers.1226[18] [22]),
    .Y(_5950_)
);

OAI21X1 _16709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf1),
    .B(_5927__bF$buf2),
    .C(_5950_),
    .Y(_4707_)
);

OAI21X1 _16710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf8),
    .B(_5894__bF$buf7),
    .C(\datapath.registers.1226[18] [23]),
    .Y(_5951_)
);

OAI21X1 _16711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf1),
    .B(_5927__bF$buf1),
    .C(_5951_),
    .Y(_4708_)
);

OAI21X1 _16712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf7),
    .B(_5894__bF$buf6),
    .C(\datapath.registers.1226[18] [24]),
    .Y(_5952_)
);

OAI21X1 _16713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf1),
    .B(_5927__bF$buf0),
    .C(_5952_),
    .Y(_4709_)
);

OAI21X1 _16714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf6),
    .B(_5894__bF$buf5),
    .C(\datapath.registers.1226[18] [25]),
    .Y(_5953_)
);

OAI21X1 _16715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486__bF$buf2),
    .B(_5927__bF$buf4),
    .C(_5953_),
    .Y(_4710_)
);

OAI21X1 _16716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf5),
    .B(_5894__bF$buf4),
    .C(\datapath.registers.1226[18] [26]),
    .Y(_5954_)
);

OAI21X1 _16717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf1),
    .B(_5927__bF$buf3),
    .C(_5954_),
    .Y(_4711_)
);

OAI21X1 _16718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf4),
    .B(_5894__bF$buf3),
    .C(\datapath.registers.1226[18] [27]),
    .Y(_5955_)
);

OAI21X1 _16719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf1),
    .B(_5927__bF$buf2),
    .C(_5955_),
    .Y(_4712_)
);

OAI21X1 _16720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf3),
    .B(_5894__bF$buf2),
    .C(\datapath.registers.1226[18] [28]),
    .Y(_5956_)
);

OAI21X1 _16721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf2),
    .B(_5927__bF$buf1),
    .C(_5956_),
    .Y(_4713_)
);

OAI21X1 _16722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf2),
    .B(_5894__bF$buf1),
    .C(\datapath.registers.1226[18] [29]),
    .Y(_5957_)
);

OAI21X1 _16723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf1),
    .B(_5927__bF$buf0),
    .C(_5957_),
    .Y(_4714_)
);

OAI21X1 _16724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf1),
    .B(_5894__bF$buf0),
    .C(\datapath.registers.1226[18] [30]),
    .Y(_5958_)
);

OAI21X1 _16725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf1),
    .B(_5927__bF$buf4),
    .C(_5958_),
    .Y(_4716_)
);

OAI21X1 _16726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf0),
    .B(_5894__bF$buf8),
    .C(\datapath.registers.1226[18] [31]),
    .Y(_5959_)
);

OAI21X1 _16727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf2),
    .B(_5927__bF$buf3),
    .C(_5959_),
    .Y(_4717_)
);

NAND2X1 _16728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5892_),
    .B(_5544_),
    .Y(_5960_)
);

OAI21X1 _16729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf15),
    .B(_5894__bF$buf7),
    .C(\datapath.registers.1226[17] [0]),
    .Y(_5961_)
);

OAI21X1 _16730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf1),
    .B(_5960__bF$buf4),
    .C(_5961_),
    .Y(_4661_)
);

OAI21X1 _16731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf14),
    .B(_5894__bF$buf6),
    .C(\datapath.registers.1226[17] [1]),
    .Y(_5962_)
);

OAI21X1 _16732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf0),
    .B(_5960__bF$buf3),
    .C(_5962_),
    .Y(_4672_)
);

OAI21X1 _16733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf13),
    .B(_5894__bF$buf5),
    .C(\datapath.registers.1226[17] [2]),
    .Y(_5963_)
);

OAI21X1 _16734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf0),
    .B(_5960__bF$buf2),
    .C(_5963_),
    .Y(_4683_)
);

OAI21X1 _16735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf12),
    .B(_5894__bF$buf4),
    .C(\datapath.registers.1226[17] [3]),
    .Y(_5964_)
);

OAI21X1 _16736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf1),
    .B(_5960__bF$buf1),
    .C(_5964_),
    .Y(_4686_)
);

OAI21X1 _16737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf11),
    .B(_5894__bF$buf3),
    .C(\datapath.registers.1226[17] [4]),
    .Y(_5965_)
);

OAI21X1 _16738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf0),
    .B(_5960__bF$buf0),
    .C(_5965_),
    .Y(_4687_)
);

OAI21X1 _16739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf10),
    .B(_5894__bF$buf2),
    .C(\datapath.registers.1226[17] [5]),
    .Y(_5966_)
);

OAI21X1 _16740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf0),
    .B(_5960__bF$buf4),
    .C(_5966_),
    .Y(_4688_)
);

OAI21X1 _16741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf9),
    .B(_5894__bF$buf1),
    .C(\datapath.registers.1226[17] [6]),
    .Y(_5967_)
);

OAI21X1 _16742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf0),
    .B(_5960__bF$buf3),
    .C(_5967_),
    .Y(_4689_)
);

OAI21X1 _16743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf8),
    .B(_5894__bF$buf0),
    .C(\datapath.registers.1226[17] [7]),
    .Y(_5968_)
);

OAI21X1 _16744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf0),
    .B(_5960__bF$buf2),
    .C(_5968_),
    .Y(_4690_)
);

OAI21X1 _16745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf7),
    .B(_5894__bF$buf8),
    .C(\datapath.registers.1226[17] [8]),
    .Y(_5969_)
);

OAI21X1 _16746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf0),
    .B(_5960__bF$buf1),
    .C(_5969_),
    .Y(_4691_)
);

OAI21X1 _16747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf6),
    .B(_5894__bF$buf7),
    .C(\datapath.registers.1226[17] [9]),
    .Y(_5970_)
);

OAI21X1 _16748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf0),
    .B(_5960__bF$buf0),
    .C(_5970_),
    .Y(_4692_)
);

OAI21X1 _16749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf5),
    .B(_5894__bF$buf6),
    .C(\datapath.registers.1226[17] [10]),
    .Y(_5971_)
);

OAI21X1 _16750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf1),
    .B(_5960__bF$buf4),
    .C(_5971_),
    .Y(_4662_)
);

OAI21X1 _16751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf4),
    .B(_5894__bF$buf5),
    .C(\datapath.registers.1226[17] [11]),
    .Y(_5972_)
);

OAI21X1 _16752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf0),
    .B(_5960__bF$buf3),
    .C(_5972_),
    .Y(_4663_)
);

OAI21X1 _16753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf3),
    .B(_5894__bF$buf4),
    .C(\datapath.registers.1226[17] [12]),
    .Y(_5973_)
);

OAI21X1 _16754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf0),
    .B(_5960__bF$buf2),
    .C(_5973_),
    .Y(_4664_)
);

OAI21X1 _16755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf2),
    .B(_5894__bF$buf3),
    .C(\datapath.registers.1226[17] [13]),
    .Y(_5974_)
);

OAI21X1 _16756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf0),
    .B(_5960__bF$buf1),
    .C(_5974_),
    .Y(_4665_)
);

OAI21X1 _16757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf1),
    .B(_5894__bF$buf2),
    .C(\datapath.registers.1226[17] [14]),
    .Y(_5975_)
);

OAI21X1 _16758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf0),
    .B(_5960__bF$buf0),
    .C(_5975_),
    .Y(_4666_)
);

OAI21X1 _16759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf0),
    .B(_5894__bF$buf1),
    .C(\datapath.registers.1226[17] [15]),
    .Y(_5976_)
);

OAI21X1 _16760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf0),
    .B(_5960__bF$buf4),
    .C(_5976_),
    .Y(_4667_)
);

OAI21X1 _16761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf15),
    .B(_5894__bF$buf0),
    .C(\datapath.registers.1226[17] [16]),
    .Y(_5977_)
);

OAI21X1 _16762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf1),
    .B(_5960__bF$buf3),
    .C(_5977_),
    .Y(_4668_)
);

OAI21X1 _16763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf14),
    .B(_5894__bF$buf8),
    .C(\datapath.registers.1226[17] [17]),
    .Y(_5978_)
);

OAI21X1 _16764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf1),
    .B(_5960__bF$buf2),
    .C(_5978_),
    .Y(_4669_)
);

OAI21X1 _16765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf13),
    .B(_5894__bF$buf7),
    .C(\datapath.registers.1226[17] [18]),
    .Y(_5979_)
);

OAI21X1 _16766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf0),
    .B(_5960__bF$buf1),
    .C(_5979_),
    .Y(_4670_)
);

OAI21X1 _16767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf12),
    .B(_5894__bF$buf6),
    .C(\datapath.registers.1226[17] [19]),
    .Y(_5980_)
);

OAI21X1 _16768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf0),
    .B(_5960__bF$buf0),
    .C(_5980_),
    .Y(_4671_)
);

OAI21X1 _16769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf11),
    .B(_5894__bF$buf5),
    .C(\datapath.registers.1226[17] [20]),
    .Y(_5981_)
);

OAI21X1 _16770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf1),
    .B(_5960__bF$buf4),
    .C(_5981_),
    .Y(_4673_)
);

OAI21X1 _16771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf10),
    .B(_5894__bF$buf4),
    .C(\datapath.registers.1226[17] [21]),
    .Y(_5982_)
);

OAI21X1 _16772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf1),
    .B(_5960__bF$buf3),
    .C(_5982_),
    .Y(_4674_)
);

OAI21X1 _16773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf9),
    .B(_5894__bF$buf3),
    .C(\datapath.registers.1226[17] [22]),
    .Y(_5983_)
);

OAI21X1 _16774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf0),
    .B(_5960__bF$buf2),
    .C(_5983_),
    .Y(_4675_)
);

OAI21X1 _16775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf8),
    .B(_5894__bF$buf2),
    .C(\datapath.registers.1226[17] [23]),
    .Y(_5984_)
);

OAI21X1 _16776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf0),
    .B(_5960__bF$buf1),
    .C(_5984_),
    .Y(_4676_)
);

OAI21X1 _16777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf7),
    .B(_5894__bF$buf1),
    .C(\datapath.registers.1226[17] [24]),
    .Y(_5985_)
);

OAI21X1 _16778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf0),
    .B(_5960__bF$buf0),
    .C(_5985_),
    .Y(_4677_)
);

OAI21X1 _16779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf6),
    .B(_5894__bF$buf0),
    .C(\datapath.registers.1226[17] [25]),
    .Y(_5986_)
);

OAI21X1 _16780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486__bF$buf1),
    .B(_5960__bF$buf4),
    .C(_5986_),
    .Y(_4678_)
);

OAI21X1 _16781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf5),
    .B(_5894__bF$buf8),
    .C(\datapath.registers.1226[17] [26]),
    .Y(_5987_)
);

OAI21X1 _16782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf0),
    .B(_5960__bF$buf3),
    .C(_5987_),
    .Y(_4679_)
);

OAI21X1 _16783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf4),
    .B(_5894__bF$buf7),
    .C(\datapath.registers.1226[17] [27]),
    .Y(_5988_)
);

OAI21X1 _16784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf0),
    .B(_5960__bF$buf2),
    .C(_5988_),
    .Y(_4680_)
);

OAI21X1 _16785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf3),
    .B(_5894__bF$buf6),
    .C(\datapath.registers.1226[17] [28]),
    .Y(_5989_)
);

OAI21X1 _16786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf1),
    .B(_5960__bF$buf1),
    .C(_5989_),
    .Y(_4681_)
);

OAI21X1 _16787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf2),
    .B(_5894__bF$buf5),
    .C(\datapath.registers.1226[17] [29]),
    .Y(_5990_)
);

OAI21X1 _16788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf0),
    .B(_5960__bF$buf0),
    .C(_5990_),
    .Y(_4682_)
);

OAI21X1 _16789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf1),
    .B(_5894__bF$buf4),
    .C(\datapath.registers.1226[17] [30]),
    .Y(_5991_)
);

OAI21X1 _16790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf0),
    .B(_5960__bF$buf4),
    .C(_5991_),
    .Y(_4684_)
);

OAI21X1 _16791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf0),
    .B(_5894__bF$buf3),
    .C(\datapath.registers.1226[17] [31]),
    .Y(_5992_)
);

OAI21X1 _16792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf1),
    .B(_5960__bF$buf3),
    .C(_5992_),
    .Y(_4685_)
);

NOR2X1 _16793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf0),
    .B(_5894__bF$buf2),
    .Y(_5993_)
);

NOR2X1 _16794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [0]),
    .B(_5993__bF$buf7),
    .Y(_5994_)
);

AOI21X1 _16795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf0),
    .B(_5993__bF$buf6),
    .C(_5994_),
    .Y(_4629_)
);

INVX1 _16796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [1]),
    .Y(_5995_)
);

NAND2X1 _16797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [1]),
    .B(_5993__bF$buf5),
    .Y(_5996_)
);

OAI21X1 _16798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5995_),
    .B(_5993__bF$buf4),
    .C(_5996_),
    .Y(_4640_)
);

NOR2X1 _16799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [2]),
    .B(_5993__bF$buf3),
    .Y(_5997_)
);

AOI21X1 _16800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf4),
    .B(_5993__bF$buf2),
    .C(_5997_),
    .Y(_4651_)
);

INVX1 _16801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [3]),
    .Y(_5998_)
);

NAND2X1 _16802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [3]),
    .B(_5993__bF$buf1),
    .Y(_5999_)
);

OAI21X1 _16803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5998_),
    .B(_5993__bF$buf0),
    .C(_5999_),
    .Y(_4654_)
);

NOR2X1 _16804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [4]),
    .B(_5993__bF$buf7),
    .Y(_6000_)
);

AOI21X1 _16805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf4),
    .B(_5993__bF$buf6),
    .C(_6000_),
    .Y(_4655_)
);

NOR2X1 _16806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [5]),
    .B(_5993__bF$buf5),
    .Y(_6001_)
);

AOI21X1 _16807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf4),
    .B(_5993__bF$buf4),
    .C(_6001_),
    .Y(_4656_)
);

INVX2 _16808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [6]),
    .Y(_6002_)
);

NAND2X1 _16809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [6]),
    .B(_5993__bF$buf3),
    .Y(_6003_)
);

OAI21X1 _16810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6002_),
    .B(_5993__bF$buf2),
    .C(_6003_),
    .Y(_4657_)
);

INVX1 _16811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [7]),
    .Y(_6004_)
);

NAND2X1 _16812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [7]),
    .B(_5993__bF$buf1),
    .Y(_6005_)
);

OAI21X1 _16813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6004_),
    .B(_5993__bF$buf0),
    .C(_6005_),
    .Y(_4658_)
);

INVX1 _16814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [8]),
    .Y(_6006_)
);

NAND2X1 _16815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [8]),
    .B(_5993__bF$buf7),
    .Y(_6007_)
);

OAI21X1 _16816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6006_),
    .B(_5993__bF$buf6),
    .C(_6007_),
    .Y(_4659_)
);

NOR2X1 _16817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [9]),
    .B(_5993__bF$buf5),
    .Y(_6008_)
);

AOI21X1 _16818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf4),
    .B(_5993__bF$buf4),
    .C(_6008_),
    .Y(_4660_)
);

INVX1 _16819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [10]),
    .Y(_6009_)
);

NAND2X1 _16820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [10]),
    .B(_5993__bF$buf3),
    .Y(_6010_)
);

OAI21X1 _16821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6009_),
    .B(_5993__bF$buf2),
    .C(_6010_),
    .Y(_4630_)
);

NOR2X1 _16822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [11]),
    .B(_5993__bF$buf1),
    .Y(_6011_)
);

AOI21X1 _16823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf4),
    .B(_5993__bF$buf0),
    .C(_6011_),
    .Y(_4631_)
);

INVX1 _16824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [12]),
    .Y(_6012_)
);

NAND2X1 _16825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [12]),
    .B(_5993__bF$buf7),
    .Y(_6013_)
);

OAI21X1 _16826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6012_),
    .B(_5993__bF$buf6),
    .C(_6013_),
    .Y(_4632_)
);

INVX1 _16827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [13]),
    .Y(_6014_)
);

NAND2X1 _16828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [13]),
    .B(_5993__bF$buf5),
    .Y(_6015_)
);

OAI21X1 _16829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6014_),
    .B(_5993__bF$buf4),
    .C(_6015_),
    .Y(_4633_)
);

NOR2X1 _16830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [14]),
    .B(_5993__bF$buf3),
    .Y(_6016_)
);

AOI21X1 _16831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf4),
    .B(_5993__bF$buf2),
    .C(_6016_),
    .Y(_4634_)
);

NOR2X1 _16832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [15]),
    .B(_5993__bF$buf1),
    .Y(_6017_)
);

AOI21X1 _16833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf4),
    .B(_5993__bF$buf0),
    .C(_6017_),
    .Y(_4635_)
);

INVX1 _16834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [16]),
    .Y(_6018_)
);

NAND2X1 _16835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [16]),
    .B(_5993__bF$buf7),
    .Y(_6019_)
);

OAI21X1 _16836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6018_),
    .B(_5993__bF$buf6),
    .C(_6019_),
    .Y(_4636_)
);

NOR2X1 _16837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [17]),
    .B(_5993__bF$buf5),
    .Y(_6020_)
);

AOI21X1 _16838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf0),
    .B(_5993__bF$buf4),
    .C(_6020_),
    .Y(_4637_)
);

NOR2X1 _16839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [18]),
    .B(_5993__bF$buf3),
    .Y(_6021_)
);

AOI21X1 _16840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf4),
    .B(_5993__bF$buf2),
    .C(_6021_),
    .Y(_4638_)
);

NOR2X1 _16841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [19]),
    .B(_5993__bF$buf1),
    .Y(_6022_)
);

AOI21X1 _16842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf4),
    .B(_5993__bF$buf0),
    .C(_6022_),
    .Y(_4639_)
);

NOR2X1 _16843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [20]),
    .B(_5993__bF$buf7),
    .Y(_6023_)
);

AOI21X1 _16844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf0),
    .B(_5993__bF$buf6),
    .C(_6023_),
    .Y(_4641_)
);

INVX1 _16845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [21]),
    .Y(_6024_)
);

NAND2X1 _16846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [21]),
    .B(_5993__bF$buf5),
    .Y(_6025_)
);

OAI21X1 _16847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6024_),
    .B(_5993__bF$buf4),
    .C(_6025_),
    .Y(_4642_)
);

INVX1 _16848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [22]),
    .Y(_6026_)
);

NAND2X1 _16849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [22]),
    .B(_5993__bF$buf3),
    .Y(_6027_)
);

OAI21X1 _16850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6026_),
    .B(_5993__bF$buf2),
    .C(_6027_),
    .Y(_4643_)
);

NOR2X1 _16851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [23]),
    .B(_5993__bF$buf1),
    .Y(_6028_)
);

AOI21X1 _16852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf4),
    .B(_5993__bF$buf0),
    .C(_6028_),
    .Y(_4644_)
);

NOR2X1 _16853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [24]),
    .B(_5993__bF$buf7),
    .Y(_6029_)
);

AOI21X1 _16854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf4),
    .B(_5993__bF$buf6),
    .C(_6029_),
    .Y(_4645_)
);

NOR2X1 _16855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [25]),
    .B(_5993__bF$buf5),
    .Y(_6030_)
);

AOI21X1 _16856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486__bF$buf0),
    .B(_5993__bF$buf4),
    .C(_6030_),
    .Y(_4646_)
);

NOR2X1 _16857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [26]),
    .B(_5993__bF$buf3),
    .Y(_6031_)
);

AOI21X1 _16858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf4),
    .B(_5993__bF$buf2),
    .C(_6031_),
    .Y(_4647_)
);

INVX1 _16859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [27]),
    .Y(_6032_)
);

NAND2X1 _16860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [27]),
    .B(_5993__bF$buf1),
    .Y(_6033_)
);

OAI21X1 _16861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6032_),
    .B(_5993__bF$buf0),
    .C(_6033_),
    .Y(_4648_)
);

NOR2X1 _16862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [28]),
    .B(_5993__bF$buf7),
    .Y(_6034_)
);

AOI21X1 _16863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf0),
    .B(_5993__bF$buf6),
    .C(_6034_),
    .Y(_4649_)
);

NOR2X1 _16864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [29]),
    .B(_5993__bF$buf5),
    .Y(_6035_)
);

AOI21X1 _16865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf4),
    .B(_5993__bF$buf4),
    .C(_6035_),
    .Y(_4650_)
);

NOR2X1 _16866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [30]),
    .B(_5993__bF$buf3),
    .Y(_6036_)
);

AOI21X1 _16867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf4),
    .B(_5993__bF$buf2),
    .C(_6036_),
    .Y(_4652_)
);

NOR2X1 _16868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[16] [31]),
    .B(_5993__bF$buf1),
    .Y(_6037_)
);

AOI21X1 _16869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf0),
    .B(_5993__bF$buf0),
    .C(_6037_),
    .Y(_4653_)
);

NAND2X1 _16870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [10]),
    .B(_5503_),
    .Y(_6038_)
);

NOR2X1 _16871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5430_),
    .B(_6038_),
    .Y(_6039_)
);

NAND2X1 _16872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5435_),
    .B(_6039_),
    .Y(_6040_)
);

INVX8 _16873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6039_),
    .Y(_6041_)
);

OAI21X1 _16874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf8),
    .B(_5434__bF$buf5),
    .C(\datapath.registers.1226[15] [0]),
    .Y(_6042_)
);

OAI21X1 _16875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf4),
    .B(_5429__bF$buf4),
    .C(_6042_),
    .Y(_4597_)
);

OAI21X1 _16876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf7),
    .B(_5434__bF$buf4),
    .C(\datapath.registers.1226[15] [1]),
    .Y(_6043_)
);

OAI21X1 _16877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf3),
    .B(_5438__bF$buf4),
    .C(_6043_),
    .Y(_4608_)
);

OAI21X1 _16878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf6),
    .B(_5434__bF$buf3),
    .C(\datapath.registers.1226[15] [2]),
    .Y(_6044_)
);

OAI21X1 _16879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf2),
    .B(_5440__bF$buf3),
    .C(_6044_),
    .Y(_4619_)
);

OAI21X1 _16880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf5),
    .B(_5434__bF$buf2),
    .C(\datapath.registers.1226[15] [3]),
    .Y(_6045_)
);

OAI21X1 _16881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf1),
    .B(_5442__bF$buf0),
    .C(_6045_),
    .Y(_4622_)
);

OAI21X1 _16882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf4),
    .B(_5434__bF$buf1),
    .C(\datapath.registers.1226[15] [4]),
    .Y(_6046_)
);

OAI21X1 _16883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf0),
    .B(_5444__bF$buf3),
    .C(_6046_),
    .Y(_4623_)
);

OAI21X1 _16884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf3),
    .B(_5434__bF$buf0),
    .C(\datapath.registers.1226[15] [5]),
    .Y(_6047_)
);

OAI21X1 _16885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf4),
    .B(_5446__bF$buf3),
    .C(_6047_),
    .Y(_4624_)
);

OAI21X1 _16886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf2),
    .B(_5434__bF$buf14),
    .C(\datapath.registers.1226[15] [6]),
    .Y(_6048_)
);

OAI21X1 _16887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf3),
    .B(_5448__bF$buf4),
    .C(_6048_),
    .Y(_4625_)
);

OAI21X1 _16888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf1),
    .B(_5434__bF$buf13),
    .C(\datapath.registers.1226[15] [7]),
    .Y(_6049_)
);

OAI21X1 _16889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf2),
    .B(_5450__bF$buf4),
    .C(_6049_),
    .Y(_4626_)
);

OAI21X1 _16890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf0),
    .B(_5434__bF$buf12),
    .C(\datapath.registers.1226[15] [8]),
    .Y(_6050_)
);

OAI21X1 _16891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf1),
    .B(_5452__bF$buf4),
    .C(_6050_),
    .Y(_4627_)
);

OAI21X1 _16892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf8),
    .B(_5434__bF$buf11),
    .C(\datapath.registers.1226[15] [9]),
    .Y(_6051_)
);

OAI21X1 _16893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf0),
    .B(_5454__bF$buf3),
    .C(_6051_),
    .Y(_4628_)
);

OAI21X1 _16894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf7),
    .B(_5434__bF$buf10),
    .C(\datapath.registers.1226[15] [10]),
    .Y(_6052_)
);

OAI21X1 _16895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf4),
    .B(_5456__bF$buf0),
    .C(_6052_),
    .Y(_4598_)
);

OAI21X1 _16896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf6),
    .B(_5434__bF$buf9),
    .C(\datapath.registers.1226[15] [11]),
    .Y(_6053_)
);

OAI21X1 _16897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf3),
    .B(_5458__bF$buf3),
    .C(_6053_),
    .Y(_4599_)
);

OAI21X1 _16898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf5),
    .B(_5434__bF$buf8),
    .C(\datapath.registers.1226[15] [12]),
    .Y(_6054_)
);

OAI21X1 _16899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf2),
    .B(_5460__bF$buf4),
    .C(_6054_),
    .Y(_4600_)
);

OAI21X1 _16900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf4),
    .B(_5434__bF$buf7),
    .C(\datapath.registers.1226[15] [13]),
    .Y(_6055_)
);

OAI21X1 _16901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf1),
    .B(_5462__bF$buf4),
    .C(_6055_),
    .Y(_4601_)
);

OAI21X1 _16902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf3),
    .B(_5434__bF$buf6),
    .C(\datapath.registers.1226[15] [14]),
    .Y(_6056_)
);

OAI21X1 _16903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf0),
    .B(_5464__bF$buf3),
    .C(_6056_),
    .Y(_4602_)
);

OAI21X1 _16904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf2),
    .B(_5434__bF$buf5),
    .C(\datapath.registers.1226[15] [15]),
    .Y(_6057_)
);

OAI21X1 _16905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf4),
    .B(_5466__bF$buf3),
    .C(_6057_),
    .Y(_4603_)
);

OAI21X1 _16906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf1),
    .B(_5434__bF$buf4),
    .C(\datapath.registers.1226[15] [16]),
    .Y(_6058_)
);

OAI21X1 _16907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf3),
    .B(_5468__bF$buf0),
    .C(_6058_),
    .Y(_4604_)
);

OAI21X1 _16908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf0),
    .B(_5434__bF$buf3),
    .C(\datapath.registers.1226[15] [17]),
    .Y(_6059_)
);

OAI21X1 _16909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf2),
    .B(_5470__bF$buf4),
    .C(_6059_),
    .Y(_4605_)
);

OAI21X1 _16910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf8),
    .B(_5434__bF$buf2),
    .C(\datapath.registers.1226[15] [18]),
    .Y(_6060_)
);

OAI21X1 _16911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf1),
    .B(_5472__bF$buf3),
    .C(_6060_),
    .Y(_4606_)
);

OAI21X1 _16912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf7),
    .B(_5434__bF$buf1),
    .C(\datapath.registers.1226[15] [19]),
    .Y(_6061_)
);

OAI21X1 _16913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf0),
    .B(_5474__bF$buf3),
    .C(_6061_),
    .Y(_4607_)
);

OAI21X1 _16914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf6),
    .B(_5434__bF$buf0),
    .C(\datapath.registers.1226[15] [20]),
    .Y(_6062_)
);

OAI21X1 _16915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf4),
    .B(_5476__bF$buf4),
    .C(_6062_),
    .Y(_4609_)
);

OAI21X1 _16916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf5),
    .B(_5434__bF$buf14),
    .C(\datapath.registers.1226[15] [21]),
    .Y(_6063_)
);

OAI21X1 _16917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf3),
    .B(_5478__bF$buf0),
    .C(_6063_),
    .Y(_4610_)
);

OAI21X1 _16918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf4),
    .B(_5434__bF$buf13),
    .C(\datapath.registers.1226[15] [22]),
    .Y(_6064_)
);

OAI21X1 _16919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf2),
    .B(_5480__bF$buf4),
    .C(_6064_),
    .Y(_4611_)
);

OAI21X1 _16920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf3),
    .B(_5434__bF$buf12),
    .C(\datapath.registers.1226[15] [23]),
    .Y(_6065_)
);

OAI21X1 _16921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf1),
    .B(_5482__bF$buf3),
    .C(_6065_),
    .Y(_4612_)
);

OAI21X1 _16922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf2),
    .B(_5434__bF$buf11),
    .C(\datapath.registers.1226[15] [24]),
    .Y(_6066_)
);

OAI21X1 _16923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf0),
    .B(_5484__bF$buf3),
    .C(_6066_),
    .Y(_4613_)
);

OAI21X1 _16924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf1),
    .B(_5434__bF$buf10),
    .C(\datapath.registers.1226[15] [25]),
    .Y(_6067_)
);

OAI21X1 _16925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf4),
    .B(_5486__bF$buf4),
    .C(_6067_),
    .Y(_4614_)
);

OAI21X1 _16926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf0),
    .B(_5434__bF$buf9),
    .C(\datapath.registers.1226[15] [26]),
    .Y(_6068_)
);

OAI21X1 _16927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf3),
    .B(_5488__bF$buf3),
    .C(_6068_),
    .Y(_4615_)
);

OAI21X1 _16928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf8),
    .B(_5434__bF$buf8),
    .C(\datapath.registers.1226[15] [27]),
    .Y(_6069_)
);

OAI21X1 _16929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf2),
    .B(_5490__bF$buf4),
    .C(_6069_),
    .Y(_4616_)
);

OAI21X1 _16930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf7),
    .B(_5434__bF$buf7),
    .C(\datapath.registers.1226[15] [28]),
    .Y(_6070_)
);

OAI21X1 _16931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf1),
    .B(_5492__bF$buf4),
    .C(_6070_),
    .Y(_4617_)
);

OAI21X1 _16932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf6),
    .B(_5434__bF$buf6),
    .C(\datapath.registers.1226[15] [29]),
    .Y(_6071_)
);

OAI21X1 _16933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf0),
    .B(_5494__bF$buf3),
    .C(_6071_),
    .Y(_4618_)
);

OAI21X1 _16934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf5),
    .B(_5434__bF$buf5),
    .C(\datapath.registers.1226[15] [30]),
    .Y(_6072_)
);

OAI21X1 _16935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf4),
    .B(_5496__bF$buf3),
    .C(_6072_),
    .Y(_4620_)
);

OAI21X1 _16936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6041__bF$buf4),
    .B(_5434__bF$buf4),
    .C(\datapath.registers.1226[15] [31]),
    .Y(_6073_)
);

OAI21X1 _16937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040__bF$buf3),
    .B(_5498__bF$buf4),
    .C(_6073_),
    .Y(_4621_)
);

NAND2X1 _16938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6039_),
    .B(_5508_),
    .Y(_6074_)
);

OAI21X1 _16939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf15),
    .B(_6041__bF$buf3),
    .C(\datapath.registers.1226[14] [0]),
    .Y(_6075_)
);

OAI21X1 _16940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf3),
    .B(_6074__bF$buf4),
    .C(_6075_),
    .Y(_4565_)
);

OAI21X1 _16941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf14),
    .B(_6041__bF$buf2),
    .C(\datapath.registers.1226[14] [1]),
    .Y(_6076_)
);

OAI21X1 _16942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf3),
    .B(_6074__bF$buf3),
    .C(_6076_),
    .Y(_4576_)
);

OAI21X1 _16943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf13),
    .B(_6041__bF$buf1),
    .C(\datapath.registers.1226[14] [2]),
    .Y(_6077_)
);

OAI21X1 _16944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf2),
    .B(_6074__bF$buf2),
    .C(_6077_),
    .Y(_4587_)
);

OAI21X1 _16945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf12),
    .B(_6041__bF$buf0),
    .C(\datapath.registers.1226[14] [3]),
    .Y(_6078_)
);

OAI21X1 _16946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf4),
    .B(_6074__bF$buf1),
    .C(_6078_),
    .Y(_4590_)
);

OAI21X1 _16947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf11),
    .B(_6041__bF$buf8),
    .C(\datapath.registers.1226[14] [4]),
    .Y(_6079_)
);

OAI21X1 _16948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf2),
    .B(_6074__bF$buf0),
    .C(_6079_),
    .Y(_4591_)
);

OAI21X1 _16949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf10),
    .B(_6041__bF$buf7),
    .C(\datapath.registers.1226[14] [5]),
    .Y(_6080_)
);

OAI21X1 _16950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf2),
    .B(_6074__bF$buf4),
    .C(_6080_),
    .Y(_4592_)
);

OAI21X1 _16951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf9),
    .B(_6041__bF$buf6),
    .C(\datapath.registers.1226[14] [6]),
    .Y(_6081_)
);

OAI21X1 _16952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf3),
    .B(_6074__bF$buf3),
    .C(_6081_),
    .Y(_4593_)
);

OAI21X1 _16953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf8),
    .B(_6041__bF$buf5),
    .C(\datapath.registers.1226[14] [7]),
    .Y(_6082_)
);

OAI21X1 _16954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf3),
    .B(_6074__bF$buf2),
    .C(_6082_),
    .Y(_4594_)
);

OAI21X1 _16955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf7),
    .B(_6041__bF$buf4),
    .C(\datapath.registers.1226[14] [8]),
    .Y(_6083_)
);

OAI21X1 _16956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf3),
    .B(_6074__bF$buf1),
    .C(_6083_),
    .Y(_4595_)
);

OAI21X1 _16957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf6),
    .B(_6041__bF$buf3),
    .C(\datapath.registers.1226[14] [9]),
    .Y(_6084_)
);

OAI21X1 _16958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf2),
    .B(_6074__bF$buf0),
    .C(_6084_),
    .Y(_4596_)
);

OAI21X1 _16959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf5),
    .B(_6041__bF$buf2),
    .C(\datapath.registers.1226[14] [10]),
    .Y(_6085_)
);

OAI21X1 _16960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf4),
    .B(_6074__bF$buf4),
    .C(_6085_),
    .Y(_4566_)
);

OAI21X1 _16961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf4),
    .B(_6041__bF$buf1),
    .C(\datapath.registers.1226[14] [11]),
    .Y(_6086_)
);

OAI21X1 _16962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf2),
    .B(_6074__bF$buf3),
    .C(_6086_),
    .Y(_4567_)
);

OAI21X1 _16963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf3),
    .B(_6041__bF$buf0),
    .C(\datapath.registers.1226[14] [12]),
    .Y(_6087_)
);

OAI21X1 _16964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf3),
    .B(_6074__bF$buf2),
    .C(_6087_),
    .Y(_4568_)
);

OAI21X1 _16965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf2),
    .B(_6041__bF$buf8),
    .C(\datapath.registers.1226[14] [13]),
    .Y(_6088_)
);

OAI21X1 _16966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf3),
    .B(_6074__bF$buf1),
    .C(_6088_),
    .Y(_4569_)
);

OAI21X1 _16967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf1),
    .B(_6041__bF$buf7),
    .C(\datapath.registers.1226[14] [14]),
    .Y(_6089_)
);

OAI21X1 _16968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf2),
    .B(_6074__bF$buf0),
    .C(_6089_),
    .Y(_4570_)
);

OAI21X1 _16969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf0),
    .B(_6041__bF$buf6),
    .C(\datapath.registers.1226[14] [15]),
    .Y(_6090_)
);

OAI21X1 _16970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf2),
    .B(_6074__bF$buf4),
    .C(_6090_),
    .Y(_4571_)
);

OAI21X1 _16971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf15),
    .B(_6041__bF$buf5),
    .C(\datapath.registers.1226[14] [16]),
    .Y(_6091_)
);

OAI21X1 _16972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf4),
    .B(_6074__bF$buf3),
    .C(_6091_),
    .Y(_4572_)
);

OAI21X1 _16973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf14),
    .B(_6041__bF$buf4),
    .C(\datapath.registers.1226[14] [17]),
    .Y(_6092_)
);

OAI21X1 _16974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf3),
    .B(_6074__bF$buf2),
    .C(_6092_),
    .Y(_4573_)
);

OAI21X1 _16975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf13),
    .B(_6041__bF$buf3),
    .C(\datapath.registers.1226[14] [18]),
    .Y(_6093_)
);

OAI21X1 _16976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf2),
    .B(_6074__bF$buf1),
    .C(_6093_),
    .Y(_4574_)
);

OAI21X1 _16977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf12),
    .B(_6041__bF$buf2),
    .C(\datapath.registers.1226[14] [19]),
    .Y(_6094_)
);

OAI21X1 _16978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf2),
    .B(_6074__bF$buf0),
    .C(_6094_),
    .Y(_4575_)
);

OAI21X1 _16979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf11),
    .B(_6041__bF$buf1),
    .C(\datapath.registers.1226[14] [20]),
    .Y(_6095_)
);

OAI21X1 _16980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf3),
    .B(_6074__bF$buf4),
    .C(_6095_),
    .Y(_4577_)
);

OAI21X1 _16981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf10),
    .B(_6041__bF$buf0),
    .C(\datapath.registers.1226[14] [21]),
    .Y(_6096_)
);

OAI21X1 _16982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf4),
    .B(_6074__bF$buf3),
    .C(_6096_),
    .Y(_4578_)
);

OAI21X1 _16983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf9),
    .B(_6041__bF$buf8),
    .C(\datapath.registers.1226[14] [22]),
    .Y(_6097_)
);

OAI21X1 _16984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf3),
    .B(_6074__bF$buf2),
    .C(_6097_),
    .Y(_4579_)
);

OAI21X1 _16985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf8),
    .B(_6041__bF$buf7),
    .C(\datapath.registers.1226[14] [23]),
    .Y(_6098_)
);

OAI21X1 _16986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf2),
    .B(_6074__bF$buf1),
    .C(_6098_),
    .Y(_4580_)
);

OAI21X1 _16987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf7),
    .B(_6041__bF$buf6),
    .C(\datapath.registers.1226[14] [24]),
    .Y(_6099_)
);

OAI21X1 _16988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf2),
    .B(_6074__bF$buf0),
    .C(_6099_),
    .Y(_4581_)
);

OAI21X1 _16989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf6),
    .B(_6041__bF$buf5),
    .C(\datapath.registers.1226[14] [25]),
    .Y(_6100_)
);

OAI21X1 _16990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486__bF$buf3),
    .B(_6074__bF$buf4),
    .C(_6100_),
    .Y(_4582_)
);

OAI21X1 _16991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf5),
    .B(_6041__bF$buf4),
    .C(\datapath.registers.1226[14] [26]),
    .Y(_6101_)
);

OAI21X1 _16992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf2),
    .B(_6074__bF$buf3),
    .C(_6101_),
    .Y(_4583_)
);

OAI21X1 _16993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf4),
    .B(_6041__bF$buf3),
    .C(\datapath.registers.1226[14] [27]),
    .Y(_6102_)
);

OAI21X1 _16994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf3),
    .B(_6074__bF$buf2),
    .C(_6102_),
    .Y(_4584_)
);

OAI21X1 _16995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf3),
    .B(_6041__bF$buf2),
    .C(\datapath.registers.1226[14] [28]),
    .Y(_6103_)
);

OAI21X1 _16996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf3),
    .B(_6074__bF$buf1),
    .C(_6103_),
    .Y(_4585_)
);

OAI21X1 _16997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf2),
    .B(_6041__bF$buf1),
    .C(\datapath.registers.1226[14] [29]),
    .Y(_6104_)
);

OAI21X1 _16998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf2),
    .B(_6074__bF$buf0),
    .C(_6104_),
    .Y(_4586_)
);

OAI21X1 _16999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf1),
    .B(_6041__bF$buf0),
    .C(\datapath.registers.1226[14] [30]),
    .Y(_6105_)
);

OAI21X1 _17000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf2),
    .B(_6074__bF$buf4),
    .C(_6105_),
    .Y(_4588_)
);

OAI21X1 _17001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf0),
    .B(_6041__bF$buf8),
    .C(\datapath.registers.1226[14] [31]),
    .Y(_6106_)
);

OAI21X1 _17002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf3),
    .B(_6074__bF$buf3),
    .C(_6106_),
    .Y(_4589_)
);

NAND2X1 _17003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6039_),
    .B(_5544_),
    .Y(_6107_)
);

OAI21X1 _17004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf15),
    .B(_6041__bF$buf7),
    .C(\datapath.registers.1226[13] [0]),
    .Y(_6108_)
);

OAI21X1 _17005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf2),
    .B(_6107__bF$buf4),
    .C(_6108_),
    .Y(_4533_)
);

OAI21X1 _17006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf14),
    .B(_6041__bF$buf6),
    .C(\datapath.registers.1226[13] [1]),
    .Y(_6109_)
);

OAI21X1 _17007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf2),
    .B(_6107__bF$buf3),
    .C(_6109_),
    .Y(_4544_)
);

OAI21X1 _17008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf13),
    .B(_6041__bF$buf5),
    .C(\datapath.registers.1226[13] [2]),
    .Y(_6110_)
);

OAI21X1 _17009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf1),
    .B(_6107__bF$buf2),
    .C(_6110_),
    .Y(_4555_)
);

OAI21X1 _17010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf12),
    .B(_6041__bF$buf4),
    .C(\datapath.registers.1226[13] [3]),
    .Y(_6111_)
);

OAI21X1 _17011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf3),
    .B(_6107__bF$buf1),
    .C(_6111_),
    .Y(_4558_)
);

OAI21X1 _17012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf11),
    .B(_6041__bF$buf3),
    .C(\datapath.registers.1226[13] [4]),
    .Y(_6112_)
);

OAI21X1 _17013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf1),
    .B(_6107__bF$buf0),
    .C(_6112_),
    .Y(_4559_)
);

OAI21X1 _17014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf10),
    .B(_6041__bF$buf2),
    .C(\datapath.registers.1226[13] [5]),
    .Y(_6113_)
);

OAI21X1 _17015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf1),
    .B(_6107__bF$buf4),
    .C(_6113_),
    .Y(_4560_)
);

OAI21X1 _17016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf9),
    .B(_6041__bF$buf1),
    .C(\datapath.registers.1226[13] [6]),
    .Y(_6114_)
);

OAI21X1 _17017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf2),
    .B(_6107__bF$buf3),
    .C(_6114_),
    .Y(_4561_)
);

OAI21X1 _17018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf8),
    .B(_6041__bF$buf0),
    .C(\datapath.registers.1226[13] [7]),
    .Y(_6115_)
);

OAI21X1 _17019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf2),
    .B(_6107__bF$buf2),
    .C(_6115_),
    .Y(_4562_)
);

OAI21X1 _17020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf7),
    .B(_6041__bF$buf8),
    .C(\datapath.registers.1226[13] [8]),
    .Y(_6116_)
);

OAI21X1 _17021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf2),
    .B(_6107__bF$buf1),
    .C(_6116_),
    .Y(_4563_)
);

OAI21X1 _17022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf6),
    .B(_6041__bF$buf7),
    .C(\datapath.registers.1226[13] [9]),
    .Y(_6117_)
);

OAI21X1 _17023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf1),
    .B(_6107__bF$buf0),
    .C(_6117_),
    .Y(_4564_)
);

OAI21X1 _17024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf5),
    .B(_6041__bF$buf6),
    .C(\datapath.registers.1226[13] [10]),
    .Y(_6118_)
);

OAI21X1 _17025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf3),
    .B(_6107__bF$buf4),
    .C(_6118_),
    .Y(_4534_)
);

OAI21X1 _17026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf4),
    .B(_6041__bF$buf5),
    .C(\datapath.registers.1226[13] [11]),
    .Y(_6119_)
);

OAI21X1 _17027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf1),
    .B(_6107__bF$buf3),
    .C(_6119_),
    .Y(_4535_)
);

OAI21X1 _17028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf3),
    .B(_6041__bF$buf4),
    .C(\datapath.registers.1226[13] [12]),
    .Y(_6120_)
);

OAI21X1 _17029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf2),
    .B(_6107__bF$buf2),
    .C(_6120_),
    .Y(_4536_)
);

OAI21X1 _17030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf2),
    .B(_6041__bF$buf3),
    .C(\datapath.registers.1226[13] [13]),
    .Y(_6121_)
);

OAI21X1 _17031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf2),
    .B(_6107__bF$buf1),
    .C(_6121_),
    .Y(_4537_)
);

OAI21X1 _17032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf1),
    .B(_6041__bF$buf2),
    .C(\datapath.registers.1226[13] [14]),
    .Y(_6122_)
);

OAI21X1 _17033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf1),
    .B(_6107__bF$buf0),
    .C(_6122_),
    .Y(_4538_)
);

OAI21X1 _17034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf0),
    .B(_6041__bF$buf1),
    .C(\datapath.registers.1226[13] [15]),
    .Y(_6123_)
);

OAI21X1 _17035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf1),
    .B(_6107__bF$buf4),
    .C(_6123_),
    .Y(_4539_)
);

OAI21X1 _17036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf15),
    .B(_6041__bF$buf0),
    .C(\datapath.registers.1226[13] [16]),
    .Y(_6124_)
);

OAI21X1 _17037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf3),
    .B(_6107__bF$buf3),
    .C(_6124_),
    .Y(_4540_)
);

OAI21X1 _17038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf14),
    .B(_6041__bF$buf8),
    .C(\datapath.registers.1226[13] [17]),
    .Y(_6125_)
);

OAI21X1 _17039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf2),
    .B(_6107__bF$buf2),
    .C(_6125_),
    .Y(_4541_)
);

OAI21X1 _17040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf13),
    .B(_6041__bF$buf7),
    .C(\datapath.registers.1226[13] [18]),
    .Y(_6126_)
);

OAI21X1 _17041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf1),
    .B(_6107__bF$buf1),
    .C(_6126_),
    .Y(_4542_)
);

OAI21X1 _17042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf12),
    .B(_6041__bF$buf6),
    .C(\datapath.registers.1226[13] [19]),
    .Y(_6127_)
);

OAI21X1 _17043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf1),
    .B(_6107__bF$buf0),
    .C(_6127_),
    .Y(_4543_)
);

OAI21X1 _17044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf11),
    .B(_6041__bF$buf5),
    .C(\datapath.registers.1226[13] [20]),
    .Y(_6128_)
);

OAI21X1 _17045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf2),
    .B(_6107__bF$buf4),
    .C(_6128_),
    .Y(_4545_)
);

OAI21X1 _17046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf10),
    .B(_6041__bF$buf4),
    .C(\datapath.registers.1226[13] [21]),
    .Y(_6129_)
);

OAI21X1 _17047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf3),
    .B(_6107__bF$buf3),
    .C(_6129_),
    .Y(_4546_)
);

OAI21X1 _17048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf9),
    .B(_6041__bF$buf3),
    .C(\datapath.registers.1226[13] [22]),
    .Y(_6130_)
);

OAI21X1 _17049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf2),
    .B(_6107__bF$buf2),
    .C(_6130_),
    .Y(_4547_)
);

OAI21X1 _17050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf8),
    .B(_6041__bF$buf2),
    .C(\datapath.registers.1226[13] [23]),
    .Y(_6131_)
);

OAI21X1 _17051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf1),
    .B(_6107__bF$buf1),
    .C(_6131_),
    .Y(_4548_)
);

OAI21X1 _17052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf7),
    .B(_6041__bF$buf1),
    .C(\datapath.registers.1226[13] [24]),
    .Y(_6132_)
);

OAI21X1 _17053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf1),
    .B(_6107__bF$buf0),
    .C(_6132_),
    .Y(_4549_)
);

OAI21X1 _17054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf6),
    .B(_6041__bF$buf0),
    .C(\datapath.registers.1226[13] [25]),
    .Y(_6133_)
);

OAI21X1 _17055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486__bF$buf2),
    .B(_6107__bF$buf4),
    .C(_6133_),
    .Y(_4550_)
);

OAI21X1 _17056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf5),
    .B(_6041__bF$buf8),
    .C(\datapath.registers.1226[13] [26]),
    .Y(_6134_)
);

OAI21X1 _17057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf1),
    .B(_6107__bF$buf3),
    .C(_6134_),
    .Y(_4551_)
);

OAI21X1 _17058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf4),
    .B(_6041__bF$buf7),
    .C(\datapath.registers.1226[13] [27]),
    .Y(_6135_)
);

OAI21X1 _17059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf2),
    .B(_6107__bF$buf2),
    .C(_6135_),
    .Y(_4552_)
);

OAI21X1 _17060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf3),
    .B(_6041__bF$buf6),
    .C(\datapath.registers.1226[13] [28]),
    .Y(_6136_)
);

OAI21X1 _17061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf2),
    .B(_6107__bF$buf1),
    .C(_6136_),
    .Y(_4553_)
);

OAI21X1 _17062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf2),
    .B(_6041__bF$buf5),
    .C(\datapath.registers.1226[13] [29]),
    .Y(_6137_)
);

OAI21X1 _17063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf1),
    .B(_6107__bF$buf0),
    .C(_6137_),
    .Y(_4554_)
);

OAI21X1 _17064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf1),
    .B(_6041__bF$buf4),
    .C(\datapath.registers.1226[13] [30]),
    .Y(_6138_)
);

OAI21X1 _17065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf1),
    .B(_6107__bF$buf4),
    .C(_6138_),
    .Y(_4556_)
);

OAI21X1 _17066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf0),
    .B(_6041__bF$buf3),
    .C(\datapath.registers.1226[13] [31]),
    .Y(_6139_)
);

OAI21X1 _17067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf2),
    .B(_6107__bF$buf3),
    .C(_6139_),
    .Y(_4557_)
);

INVX8 _17068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_19_bF$buf2 ),
    .Y(_6140_)
);

INVX8 _17069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf50 ),
    .Y(_6141_)
);

NAND2X1 _17070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6140__bF$buf4),
    .B(_6141__bF$buf10),
    .Y(_6142_)
);

INVX8 _17071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_bF$buf42 ),
    .Y(_6143_)
);

INVX8 _17072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf38 ),
    .Y(_6144_)
);

INVX8 _17073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_18_bF$buf4 ),
    .Y(_6145_)
);

NAND3X1 _17074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf4),
    .B(_6144__bF$buf10),
    .C(_6145__bF$buf7),
    .Y(_6146_)
);

NOR2X1 _17075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6142_),
    .B(_6146_),
    .Y(_6147_)
);

INVX1 _17076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [0]),
    .Y(_6148_)
);

AOI21X1 _17077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [0]),
    .B(\datapath.idinstr_17_bF$buf37 ),
    .C(_6141__bF$buf9),
    .Y(_6149_)
);

OAI21X1 _17078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6148_),
    .B(\datapath.idinstr_17_bF$buf36 ),
    .C(_6149_),
    .Y(_6150_)
);

INVX1 _17079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [0]),
    .Y(_6151_)
);

AOI21X1 _17080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [0]),
    .B(\datapath.idinstr_17_bF$buf35 ),
    .C(\datapath.idinstr_15_bF$buf49 ),
    .Y(_6152_)
);

OAI21X1 _17081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6151_),
    .B(\datapath.idinstr_17_bF$buf34 ),
    .C(_6152_),
    .Y(_6153_)
);

NAND3X1 _17082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf3),
    .B(_6153_),
    .C(_6150_),
    .Y(_6154_)
);

INVX2 _17083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [0]),
    .Y(_6155_)
);

AOI21X1 _17084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [0]),
    .B(\datapath.idinstr_17_bF$buf33 ),
    .C(_6141__bF$buf8),
    .Y(_6156_)
);

OAI21X1 _17085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6155_),
    .B(\datapath.idinstr_17_bF$buf32 ),
    .C(_6156_),
    .Y(_6157_)
);

INVX1 _17086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[2] [0]),
    .Y(_6158_)
);

AOI21X1 _17087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[6] [0]),
    .B(\datapath.idinstr_17_bF$buf31 ),
    .C(\datapath.idinstr_15_bF$buf48 ),
    .Y(_6159_)
);

OAI21X1 _17088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6158_),
    .B(\datapath.idinstr_17_bF$buf30 ),
    .C(_6159_),
    .Y(_6160_)
);

NAND3X1 _17089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_bF$buf41 ),
    .B(_6160_),
    .C(_6157_),
    .Y(_6161_)
);

AOI21X1 _17090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6154_),
    .B(_6161_),
    .C(\datapath.idinstr_18_bF$buf3 ),
    .Y(_6162_)
);

MUX2X1 _17091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [0]),
    .B(\datapath.registers.1226[8] [0]),
    .S(\datapath.idinstr_15_bF$buf47 ),
    .Y(_6163_)
);

MUX2X1 _17092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [0]),
    .B(\datapath.registers.1226[10] [0]),
    .S(\datapath.idinstr_15_bF$buf46 ),
    .Y(_6164_)
);

MUX2X1 _17093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6164_),
    .B(_6163_),
    .S(\datapath.idinstr_16_bF$buf40 ),
    .Y(_6165_)
);

NAND2X1 _17094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf9),
    .B(_6165_),
    .Y(_6166_)
);

MUX2X1 _17095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [0]),
    .B(\datapath.registers.1226[12] [0]),
    .S(\datapath.idinstr_15_bF$buf45 ),
    .Y(_6167_)
);

MUX2X1 _17096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [0]),
    .B(\datapath.registers.1226[14] [0]),
    .S(\datapath.idinstr_15_bF$buf44 ),
    .Y(_6168_)
);

MUX2X1 _17097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6168_),
    .B(_6167_),
    .S(\datapath.idinstr_16_bF$buf39 ),
    .Y(_6169_)
);

NAND2X1 _17098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf29 ),
    .B(_6169_),
    .Y(_6170_)
);

AOI21X1 _17099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6166_),
    .B(_6170_),
    .C(_6145__bF$buf6),
    .Y(_6171_)
);

OAI21X1 _17100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6171_),
    .B(_6162_),
    .C(_6140__bF$buf3),
    .Y(_6172_)
);

MUX2X1 _17101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [0]),
    .B(\datapath.registers.1226[16] [0]),
    .S(\datapath.idinstr_15_bF$buf43 ),
    .Y(_6173_)
);

MUX2X1 _17102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [0]),
    .B(\datapath.registers.1226[18] [0]),
    .S(\datapath.idinstr_15_bF$buf42 ),
    .Y(_6174_)
);

MUX2X1 _17103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6174_),
    .B(_6173_),
    .S(\datapath.idinstr_16_bF$buf38 ),
    .Y(_6175_)
);

NAND2X1 _17104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf8),
    .B(_6175_),
    .Y(_6176_)
);

MUX2X1 _17105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [0]),
    .B(\datapath.registers.1226[20] [0]),
    .S(\datapath.idinstr_15_bF$buf41 ),
    .Y(_6177_)
);

MUX2X1 _17106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [0]),
    .B(\datapath.registers.1226[22] [0]),
    .S(\datapath.idinstr_15_bF$buf40 ),
    .Y(_6178_)
);

MUX2X1 _17107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6178_),
    .B(_6177_),
    .S(\datapath.idinstr_16_bF$buf37 ),
    .Y(_6179_)
);

NAND2X1 _17108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf28 ),
    .B(_6179_),
    .Y(_6180_)
);

AOI21X1 _17109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6176_),
    .B(_6180_),
    .C(\datapath.idinstr_18_bF$buf2 ),
    .Y(_6181_)
);

INVX1 _17110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [0]),
    .Y(_6182_)
);

AOI21X1 _17111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [0]),
    .B(\datapath.idinstr_17_bF$buf27 ),
    .C(_6141__bF$buf7),
    .Y(_6183_)
);

OAI21X1 _17112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6182_),
    .B(\datapath.idinstr_17_bF$buf26 ),
    .C(_6183_),
    .Y(_6184_)
);

NAND2X1 _17113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [0]),
    .B(_6144__bF$buf7),
    .Y(_6185_)
);

AOI21X1 _17114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [0]),
    .B(\datapath.idinstr_17_bF$buf25 ),
    .C(\datapath.idinstr_15_bF$buf39 ),
    .Y(_6186_)
);

AOI21X1 _17115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6186_),
    .B(_6185_),
    .C(_6143__bF$buf2),
    .Y(_6187_)
);

NAND2X1 _17116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6184_),
    .B(_6187_),
    .Y(_6188_)
);

INVX1 _17117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [0]),
    .Y(_6189_)
);

AOI21X1 _17118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [0]),
    .B(\datapath.idinstr_17_bF$buf24 ),
    .C(_6141__bF$buf6),
    .Y(_6190_)
);

OAI21X1 _17119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6189_),
    .B(\datapath.idinstr_17_bF$buf23 ),
    .C(_6190_),
    .Y(_6191_)
);

AOI21X1 _17120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[28] [0]),
    .B(\datapath.idinstr_17_bF$buf22 ),
    .C(\datapath.idinstr_15_bF$buf38 ),
    .Y(_6192_)
);

OAI21X1 _17121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5714_),
    .B(\datapath.idinstr_17_bF$buf21 ),
    .C(_6192_),
    .Y(_6193_)
);

NAND3X1 _17122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf1),
    .B(_6193_),
    .C(_6191_),
    .Y(_6194_)
);

AOI21X1 _17123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6188_),
    .B(_6194_),
    .C(_6145__bF$buf5),
    .Y(_6195_)
);

OAI21X1 _17124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6181_),
    .B(_6195_),
    .C(\datapath.idinstr_19_bF$buf1 ),
    .Y(_6196_)
);

AOI21X1 _17125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6196_),
    .B(_6172_),
    .C(_6147__bF$buf4),
    .Y(\datapath.registers.rega_data [0])
);

MUX2X1 _17126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [1]),
    .B(\datapath.registers.1226[8] [1]),
    .S(\datapath.idinstr_15_bF$buf37 ),
    .Y(_6197_)
);

MUX2X1 _17127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [1]),
    .B(\datapath.registers.1226[10] [1]),
    .S(\datapath.idinstr_15_bF$buf36 ),
    .Y(_6198_)
);

MUX2X1 _17128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6198_),
    .B(_6197_),
    .S(\datapath.idinstr_16_bF$buf36 ),
    .Y(_6199_)
);

NAND2X1 _17129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf6),
    .B(_6199_),
    .Y(_6200_)
);

MUX2X1 _17130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [1]),
    .B(\datapath.registers.1226[12] [1]),
    .S(\datapath.idinstr_15_bF$buf35 ),
    .Y(_6201_)
);

MUX2X1 _17131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [1]),
    .B(\datapath.registers.1226[14] [1]),
    .S(\datapath.idinstr_15_bF$buf34 ),
    .Y(_6202_)
);

MUX2X1 _17132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6202_),
    .B(_6201_),
    .S(\datapath.idinstr_16_bF$buf35 ),
    .Y(_6203_)
);

NAND2X1 _17133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf20 ),
    .B(_6203_),
    .Y(_6204_)
);

AOI21X1 _17134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6200_),
    .B(_6204_),
    .C(_6145__bF$buf4),
    .Y(_6205_)
);

INVX1 _17135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [1]),
    .Y(_6206_)
);

AOI21X1 _17136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf19 ),
    .B(\datapath.registers.1226[5] [1]),
    .C(_6141__bF$buf5),
    .Y(_6207_)
);

OAI21X1 _17137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf18 ),
    .B(_6206_),
    .C(_6207_),
    .Y(_6208_)
);

NAND2X1 _17138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [1]),
    .B(_6144__bF$buf5),
    .Y(_6209_)
);

AOI21X1 _17139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf17 ),
    .B(\datapath.registers.1226[4] [1]),
    .C(\datapath.idinstr_15_bF$buf33 ),
    .Y(_6210_)
);

AOI21X1 _17140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6210_),
    .B(_6209_),
    .C(\datapath.idinstr_16_bF$buf34 ),
    .Y(_6211_)
);

NAND2X1 _17141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6208_),
    .B(_6211_),
    .Y(_6212_)
);

INVX2 _17142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [1]),
    .Y(_6213_)
);

AOI21X1 _17143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf16 ),
    .B(\datapath.registers.1226[7] [1]),
    .C(_6141__bF$buf4),
    .Y(_6214_)
);

OAI21X1 _17144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf15 ),
    .B(_6213_),
    .C(_6214_),
    .Y(_6215_)
);

INVX1 _17145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[2] [1]),
    .Y(_6216_)
);

AOI21X1 _17146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf14 ),
    .B(\datapath.registers.1226[6] [1]),
    .C(\datapath.idinstr_15_bF$buf32 ),
    .Y(_6217_)
);

OAI21X1 _17147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf13 ),
    .B(_6216_),
    .C(_6217_),
    .Y(_6218_)
);

NAND3X1 _17148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_bF$buf33 ),
    .B(_6218_),
    .C(_6215_),
    .Y(_6219_)
);

AOI21X1 _17149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6212_),
    .B(_6219_),
    .C(\datapath.idinstr_18_bF$buf1 ),
    .Y(_6220_)
);

OAI21X1 _17150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6205_),
    .B(_6220_),
    .C(_6140__bF$buf2),
    .Y(_6221_)
);

MUX2X1 _17151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [1]),
    .B(\datapath.registers.1226[29] [1]),
    .S(\datapath.idinstr_16_bF$buf32 ),
    .Y(_6222_)
);

MUX2X1 _17152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [1]),
    .B(\datapath.registers.1226[28] [1]),
    .S(\datapath.idinstr_16_bF$buf31 ),
    .Y(_6223_)
);

MUX2X1 _17153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6223_),
    .B(_6222_),
    .S(_6141__bF$buf3),
    .Y(_6224_)
);

NAND2X1 _17154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf12 ),
    .B(_6224_),
    .Y(_6225_)
);

MUX2X1 _17155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [1]),
    .B(\datapath.registers.1226[25] [1]),
    .S(\datapath.idinstr_16_bF$buf30 ),
    .Y(_6226_)
);

MUX2X1 _17156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [1]),
    .B(\datapath.registers.1226[24] [1]),
    .S(\datapath.idinstr_16_bF$buf29 ),
    .Y(_6227_)
);

MUX2X1 _17157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6227_),
    .B(_6226_),
    .S(_6141__bF$buf2),
    .Y(_6228_)
);

NAND2X1 _17158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf4),
    .B(_6228_),
    .Y(_6229_)
);

AOI21X1 _17159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6225_),
    .B(_6229_),
    .C(_6145__bF$buf3),
    .Y(_6230_)
);

INVX1 _17160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [1]),
    .Y(_6231_)
);

AOI21X1 _17161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [1]),
    .B(\datapath.idinstr_17_bF$buf11 ),
    .C(_6141__bF$buf1),
    .Y(_6232_)
);

OAI21X1 _17162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6231_),
    .B(\datapath.idinstr_17_bF$buf10 ),
    .C(_6232_),
    .Y(_6233_)
);

INVX1 _17163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [1]),
    .Y(_6234_)
);

AOI21X1 _17164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [1]),
    .B(\datapath.idinstr_17_bF$buf9 ),
    .C(\datapath.idinstr_15_bF$buf31 ),
    .Y(_6235_)
);

OAI21X1 _17165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6234_),
    .B(\datapath.idinstr_17_bF$buf8 ),
    .C(_6235_),
    .Y(_6236_)
);

NAND3X1 _17166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_bF$buf28 ),
    .B(_6236_),
    .C(_6233_),
    .Y(_6237_)
);

INVX1 _17167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [1]),
    .Y(_6238_)
);

AOI21X1 _17168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [1]),
    .B(\datapath.idinstr_17_bF$buf7 ),
    .C(_6141__bF$buf0),
    .Y(_6239_)
);

OAI21X1 _17169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6238_),
    .B(\datapath.idinstr_17_bF$buf6 ),
    .C(_6239_),
    .Y(_6240_)
);

AOI21X1 _17170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [1]),
    .B(\datapath.idinstr_17_bF$buf5 ),
    .C(\datapath.idinstr_15_bF$buf30 ),
    .Y(_6241_)
);

OAI21X1 _17171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5995_),
    .B(\datapath.idinstr_17_bF$buf4 ),
    .C(_6241_),
    .Y(_6242_)
);

NAND3X1 _17172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf0),
    .B(_6242_),
    .C(_6240_),
    .Y(_6243_)
);

AOI21X1 _17173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6237_),
    .B(_6243_),
    .C(\datapath.idinstr_18_bF$buf0 ),
    .Y(_6244_)
);

OAI21X1 _17174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6230_),
    .B(_6244_),
    .C(\datapath.idinstr_19_bF$buf0 ),
    .Y(_6245_)
);

AOI21X1 _17175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6221_),
    .B(_6245_),
    .C(_6147__bF$buf3),
    .Y(\datapath.registers.rega_data [1])
);

MUX2X1 _17176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [2]),
    .B(\datapath.registers.1226[24] [2]),
    .S(\datapath.idinstr_15_bF$buf29 ),
    .Y(_6246_)
);

MUX2X1 _17177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [2]),
    .B(\datapath.registers.1226[26] [2]),
    .S(\datapath.idinstr_15_bF$buf28 ),
    .Y(_6247_)
);

MUX2X1 _17178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6247_),
    .B(_6246_),
    .S(\datapath.idinstr_16_bF$buf27 ),
    .Y(_6248_)
);

NAND2X1 _17179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf3),
    .B(_6248_),
    .Y(_6249_)
);

MUX2X1 _17180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [2]),
    .B(\datapath.registers.1226[28] [2]),
    .S(\datapath.idinstr_15_bF$buf27 ),
    .Y(_6250_)
);

MUX2X1 _17181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [2]),
    .B(\datapath.registers.1226[30] [2]),
    .S(\datapath.idinstr_15_bF$buf26 ),
    .Y(_6251_)
);

MUX2X1 _17182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6251_),
    .B(_6250_),
    .S(\datapath.idinstr_16_bF$buf26 ),
    .Y(_6252_)
);

NAND2X1 _17183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf3 ),
    .B(_6252_),
    .Y(_6253_)
);

AOI21X1 _17184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6249_),
    .B(_6253_),
    .C(_6145__bF$buf2),
    .Y(_6254_)
);

MUX2X1 _17185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [2]),
    .B(\datapath.registers.1226[16] [2]),
    .S(\datapath.idinstr_16_bF$buf25 ),
    .Y(_6255_)
);

NAND2X1 _17186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf10),
    .B(_6255_),
    .Y(_6256_)
);

MUX2X1 _17187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [2]),
    .B(\datapath.registers.1226[17] [2]),
    .S(\datapath.idinstr_16_bF$buf24 ),
    .Y(_6257_)
);

AOI21X1 _17188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf25 ),
    .B(_6257_),
    .C(\datapath.idinstr_17_bF$buf2 ),
    .Y(_6258_)
);

NAND2X1 _17189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6256_),
    .B(_6258_),
    .Y(_6259_)
);

MUX2X1 _17190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [2]),
    .B(\datapath.registers.1226[20] [2]),
    .S(\datapath.idinstr_16_bF$buf23 ),
    .Y(_6260_)
);

NAND2X1 _17191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf9),
    .B(_6260_),
    .Y(_6261_)
);

MUX2X1 _17192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [2]),
    .B(\datapath.registers.1226[21] [2]),
    .S(\datapath.idinstr_16_bF$buf22 ),
    .Y(_6262_)
);

AOI21X1 _17193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf24 ),
    .B(_6262_),
    .C(_6144__bF$buf2),
    .Y(_6263_)
);

NAND2X1 _17194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6261_),
    .B(_6263_),
    .Y(_6264_)
);

AOI21X1 _17195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6259_),
    .B(_6264_),
    .C(\datapath.idinstr_18_bF$buf7 ),
    .Y(_6265_)
);

OAI21X1 _17196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6254_),
    .B(_6265_),
    .C(\datapath.idinstr_19_bF$buf5 ),
    .Y(_6266_)
);

MUX2X1 _17197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [2]),
    .B(\datapath.registers.1226[8] [2]),
    .S(\datapath.idinstr_15_bF$buf23 ),
    .Y(_6267_)
);

MUX2X1 _17198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [2]),
    .B(\datapath.registers.1226[10] [2]),
    .S(\datapath.idinstr_15_bF$buf22 ),
    .Y(_6268_)
);

MUX2X1 _17199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6268_),
    .B(_6267_),
    .S(\datapath.idinstr_16_bF$buf21 ),
    .Y(_6269_)
);

NAND2X1 _17200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf1),
    .B(_6269_),
    .Y(_6270_)
);

MUX2X1 _17201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [2]),
    .B(\datapath.registers.1226[12] [2]),
    .S(\datapath.idinstr_15_bF$buf21 ),
    .Y(_6271_)
);

MUX2X1 _17202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [2]),
    .B(\datapath.registers.1226[14] [2]),
    .S(\datapath.idinstr_15_bF$buf20 ),
    .Y(_6272_)
);

MUX2X1 _17203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6272_),
    .B(_6271_),
    .S(\datapath.idinstr_16_bF$buf20 ),
    .Y(_6273_)
);

NAND2X1 _17204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf1 ),
    .B(_6273_),
    .Y(_6274_)
);

AOI21X1 _17205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6270_),
    .B(_6274_),
    .C(_6145__bF$buf1),
    .Y(_6275_)
);

INVX1 _17206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [2]),
    .Y(_6276_)
);

AOI21X1 _17207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf0 ),
    .B(\datapath.registers.1226[5] [2]),
    .C(_6141__bF$buf8),
    .Y(_6277_)
);

OAI21X1 _17208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf41 ),
    .B(_6276_),
    .C(_6277_),
    .Y(_6278_)
);

INVX1 _17209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [2]),
    .Y(_6279_)
);

AOI21X1 _17210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf40 ),
    .B(\datapath.registers.1226[4] [2]),
    .C(\datapath.idinstr_15_bF$buf19 ),
    .Y(_6280_)
);

OAI21X1 _17211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6279_),
    .B(\datapath.idinstr_17_bF$buf39 ),
    .C(_6280_),
    .Y(_6281_)
);

NAND3X1 _17212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf4),
    .B(_6281_),
    .C(_6278_),
    .Y(_6282_)
);

INVX1 _17213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [2]),
    .Y(_6283_)
);

AOI21X1 _17214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf38 ),
    .B(\datapath.registers.1226[7] [2]),
    .C(_6141__bF$buf7),
    .Y(_6284_)
);

OAI21X1 _17215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf37 ),
    .B(_6283_),
    .C(_6284_),
    .Y(_6285_)
);

INVX1 _17216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[2] [2]),
    .Y(_6286_)
);

AOI21X1 _17217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf36 ),
    .B(\datapath.registers.1226[6] [2]),
    .C(\datapath.idinstr_15_bF$buf18 ),
    .Y(_6287_)
);

OAI21X1 _17218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf35 ),
    .B(_6286_),
    .C(_6287_),
    .Y(_6288_)
);

NAND3X1 _17219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_bF$buf19 ),
    .B(_6288_),
    .C(_6285_),
    .Y(_6289_)
);

AOI21X1 _17220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6282_),
    .B(_6289_),
    .C(\datapath.idinstr_18_bF$buf6 ),
    .Y(_6290_)
);

OAI21X1 _17221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6275_),
    .B(_6290_),
    .C(_6140__bF$buf1),
    .Y(_6291_)
);

AOI21X1 _17222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6266_),
    .B(_6291_),
    .C(_6147__bF$buf2),
    .Y(\datapath.registers.rega_data [2])
);

MUX2X1 _17223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [3]),
    .B(\datapath.registers.1226[8] [3]),
    .S(\datapath.idinstr_15_bF$buf17 ),
    .Y(_6292_)
);

MUX2X1 _17224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [3]),
    .B(\datapath.registers.1226[10] [3]),
    .S(\datapath.idinstr_15_bF$buf16 ),
    .Y(_6293_)
);

MUX2X1 _17225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6293_),
    .B(_6292_),
    .S(\datapath.idinstr_16_bF$buf18 ),
    .Y(_6294_)
);

NAND2X1 _17226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf0),
    .B(_6294_),
    .Y(_6295_)
);

AND2X2 _17227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [3]),
    .B(\datapath.idinstr_15_bF$buf15 ),
    .Y(_6296_)
);

INVX1 _17228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [3]),
    .Y(_6297_)
);

OAI21X1 _17229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6297_),
    .B(\datapath.idinstr_15_bF$buf14 ),
    .C(\datapath.idinstr_16_bF$buf17 ),
    .Y(_6298_)
);

NAND2X1 _17230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [3]),
    .B(_6141__bF$buf6),
    .Y(_6299_)
);

AOI21X1 _17231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [3]),
    .B(\datapath.idinstr_15_bF$buf13 ),
    .C(\datapath.idinstr_16_bF$buf16 ),
    .Y(_6300_)
);

AOI21X1 _17232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6300_),
    .B(_6299_),
    .C(_6144__bF$buf10),
    .Y(_6301_)
);

OAI21X1 _17233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6296_),
    .B(_6298_),
    .C(_6301_),
    .Y(_6302_)
);

AOI21X1 _17234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6302_),
    .B(_6295_),
    .C(_6145__bF$buf0),
    .Y(_6303_)
);

MUX2X1 _17235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [3]),
    .B(\datapath.registers.1226[4] [3]),
    .S(\datapath.idinstr_15_bF$buf12 ),
    .Y(_6304_)
);

MUX2X1 _17236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [3]),
    .B(\datapath.registers.1226[6] [3]),
    .S(\datapath.idinstr_15_bF$buf11 ),
    .Y(_6305_)
);

MUX2X1 _17237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6305_),
    .B(_6304_),
    .S(\datapath.idinstr_16_bF$buf15 ),
    .Y(_6306_)
);

NAND2X1 _17238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf34 ),
    .B(_6306_),
    .Y(_6307_)
);

MUX2X1 _17239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [3]),
    .B(\datapath.registers.1226[0] [3]),
    .S(\datapath.idinstr_15_bF$buf10 ),
    .Y(_6308_)
);

MUX2X1 _17240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [3]),
    .B(\datapath.registers.1226[2] [3]),
    .S(\datapath.idinstr_15_bF$buf9 ),
    .Y(_6309_)
);

MUX2X1 _17241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6309_),
    .B(_6308_),
    .S(\datapath.idinstr_16_bF$buf14 ),
    .Y(_6310_)
);

NAND2X1 _17242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf9),
    .B(_6310_),
    .Y(_6311_)
);

AOI21X1 _17243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6307_),
    .B(_6311_),
    .C(\datapath.idinstr_18_bF$buf5 ),
    .Y(_6312_)
);

OAI21X1 _17244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6312_),
    .B(_6303_),
    .C(_6140__bF$buf0),
    .Y(_6313_)
);

INVX1 _17245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [3]),
    .Y(_6314_)
);

AOI21X1 _17246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [3]),
    .B(\datapath.idinstr_17_bF$buf33 ),
    .C(_6141__bF$buf5),
    .Y(_6315_)
);

OAI21X1 _17247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6314_),
    .B(\datapath.idinstr_17_bF$buf32 ),
    .C(_6315_),
    .Y(_6316_)
);

NAND2X1 _17248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [3]),
    .B(_6144__bF$buf8),
    .Y(_6317_)
);

AOI21X1 _17249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [3]),
    .B(\datapath.idinstr_17_bF$buf31 ),
    .C(\datapath.idinstr_15_bF$buf8 ),
    .Y(_6318_)
);

AOI21X1 _17250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6318_),
    .B(_6317_),
    .C(_6143__bF$buf3),
    .Y(_6319_)
);

NAND2X1 _17251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6316_),
    .B(_6319_),
    .Y(_6320_)
);

INVX1 _17252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [3]),
    .Y(_6321_)
);

AOI21X1 _17253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [3]),
    .B(\datapath.idinstr_17_bF$buf30 ),
    .C(_6141__bF$buf4),
    .Y(_6322_)
);

OAI21X1 _17254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6321_),
    .B(\datapath.idinstr_17_bF$buf29 ),
    .C(_6322_),
    .Y(_6323_)
);

AOI21X1 _17255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [3]),
    .B(\datapath.idinstr_17_bF$buf28 ),
    .C(\datapath.idinstr_15_bF$buf7 ),
    .Y(_6324_)
);

OAI21X1 _17256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5998_),
    .B(\datapath.idinstr_17_bF$buf27 ),
    .C(_6324_),
    .Y(_6325_)
);

NAND3X1 _17257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf2),
    .B(_6325_),
    .C(_6323_),
    .Y(_6326_)
);

AOI21X1 _17258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6320_),
    .B(_6326_),
    .C(\datapath.idinstr_18_bF$buf4 ),
    .Y(_6327_)
);

MUX2X1 _17259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [3]),
    .B(\datapath.registers.1226[29] [3]),
    .S(\datapath.idinstr_16_bF$buf13 ),
    .Y(_6328_)
);

MUX2X1 _17260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [3]),
    .B(\datapath.registers.1226[28] [3]),
    .S(\datapath.idinstr_16_bF$buf12 ),
    .Y(_6329_)
);

MUX2X1 _17261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6329_),
    .B(_6328_),
    .S(_6141__bF$buf3),
    .Y(_6330_)
);

NAND2X1 _17262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf26 ),
    .B(_6330_),
    .Y(_6331_)
);

MUX2X1 _17263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [3]),
    .B(\datapath.registers.1226[25] [3]),
    .S(\datapath.idinstr_16_bF$buf11 ),
    .Y(_6332_)
);

MUX2X1 _17264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [3]),
    .B(\datapath.registers.1226[24] [3]),
    .S(\datapath.idinstr_16_bF$buf10 ),
    .Y(_6333_)
);

MUX2X1 _17265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6333_),
    .B(_6332_),
    .S(_6141__bF$buf2),
    .Y(_6334_)
);

NAND2X1 _17266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf7),
    .B(_6334_),
    .Y(_6335_)
);

AOI21X1 _17267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6331_),
    .B(_6335_),
    .C(_6145__bF$buf7),
    .Y(_6336_)
);

OAI21X1 _17268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6336_),
    .B(_6327_),
    .C(\datapath.idinstr_19_bF$buf4 ),
    .Y(_6337_)
);

AOI21X1 _17269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6337_),
    .B(_6313_),
    .C(_6147__bF$buf1),
    .Y(\datapath.registers.rega_data [3])
);

MUX2X1 _17270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [4]),
    .B(\datapath.registers.1226[24] [4]),
    .S(\datapath.idinstr_15_bF$buf6 ),
    .Y(_6338_)
);

MUX2X1 _17271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [4]),
    .B(\datapath.registers.1226[26] [4]),
    .S(\datapath.idinstr_15_bF$buf5 ),
    .Y(_6339_)
);

MUX2X1 _17272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6339_),
    .B(_6338_),
    .S(\datapath.idinstr_16_bF$buf9 ),
    .Y(_6340_)
);

NAND2X1 _17273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf6),
    .B(_6340_),
    .Y(_6341_)
);

MUX2X1 _17274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [4]),
    .B(\datapath.registers.1226[28] [4]),
    .S(\datapath.idinstr_15_bF$buf4 ),
    .Y(_6342_)
);

MUX2X1 _17275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [4]),
    .B(\datapath.registers.1226[30] [4]),
    .S(\datapath.idinstr_15_bF$buf3 ),
    .Y(_6343_)
);

MUX2X1 _17276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6343_),
    .B(_6342_),
    .S(\datapath.idinstr_16_bF$buf8 ),
    .Y(_6344_)
);

NAND2X1 _17277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf25 ),
    .B(_6344_),
    .Y(_6345_)
);

AOI21X1 _17278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6341_),
    .B(_6345_),
    .C(_6145__bF$buf6),
    .Y(_6346_)
);

MUX2X1 _17279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [4]),
    .B(\datapath.registers.1226[16] [4]),
    .S(\datapath.idinstr_16_bF$buf7 ),
    .Y(_6347_)
);

NAND2X1 _17280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf1),
    .B(_6347_),
    .Y(_6348_)
);

MUX2X1 _17281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [4]),
    .B(\datapath.registers.1226[17] [4]),
    .S(\datapath.idinstr_16_bF$buf6 ),
    .Y(_6349_)
);

AOI21X1 _17282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf2 ),
    .B(_6349_),
    .C(\datapath.idinstr_17_bF$buf24 ),
    .Y(_6350_)
);

NAND2X1 _17283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6348_),
    .B(_6350_),
    .Y(_6351_)
);

MUX2X1 _17284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [4]),
    .B(\datapath.registers.1226[20] [4]),
    .S(\datapath.idinstr_16_bF$buf5 ),
    .Y(_6352_)
);

NAND2X1 _17285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf0),
    .B(_6352_),
    .Y(_6353_)
);

MUX2X1 _17286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [4]),
    .B(\datapath.registers.1226[21] [4]),
    .S(\datapath.idinstr_16_bF$buf4 ),
    .Y(_6354_)
);

AOI21X1 _17287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf1 ),
    .B(_6354_),
    .C(_6144__bF$buf5),
    .Y(_6355_)
);

NAND2X1 _17288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6353_),
    .B(_6355_),
    .Y(_6356_)
);

AOI21X1 _17289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6351_),
    .B(_6356_),
    .C(\datapath.idinstr_18_bF$buf3 ),
    .Y(_6357_)
);

OAI21X1 _17290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6346_),
    .B(_6357_),
    .C(\datapath.idinstr_19_bF$buf3 ),
    .Y(_6358_)
);

MUX2X1 _17291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [4]),
    .B(\datapath.registers.1226[8] [4]),
    .S(\datapath.idinstr_15_bF$buf0 ),
    .Y(_6359_)
);

MUX2X1 _17292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [4]),
    .B(\datapath.registers.1226[10] [4]),
    .S(\datapath.idinstr_15_bF$buf53 ),
    .Y(_6360_)
);

MUX2X1 _17293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6360_),
    .B(_6359_),
    .S(\datapath.idinstr_16_bF$buf3 ),
    .Y(_6361_)
);

NAND2X1 _17294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf4),
    .B(_6361_),
    .Y(_6362_)
);

INVX1 _17295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [4]),
    .Y(_6363_)
);

NOR2X1 _17296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6363_),
    .B(_6141__bF$buf10),
    .Y(_6364_)
);

INVX1 _17297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [4]),
    .Y(_6365_)
);

OAI21X1 _17298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6365_),
    .B(\datapath.idinstr_15_bF$buf52 ),
    .C(\datapath.idinstr_16_bF$buf2 ),
    .Y(_6366_)
);

NAND2X1 _17299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [4]),
    .B(_6141__bF$buf9),
    .Y(_6367_)
);

AOI21X1 _17300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [4]),
    .B(\datapath.idinstr_15_bF$buf51 ),
    .C(\datapath.idinstr_16_bF$buf1 ),
    .Y(_6368_)
);

AOI21X1 _17301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6368_),
    .B(_6367_),
    .C(_6144__bF$buf3),
    .Y(_6369_)
);

OAI21X1 _17302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6364_),
    .B(_6366_),
    .C(_6369_),
    .Y(_6370_)
);

AOI21X1 _17303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6370_),
    .B(_6362_),
    .C(_6145__bF$buf5),
    .Y(_6371_)
);

MUX2X1 _17304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [4]),
    .B(\datapath.registers.1226[4] [4]),
    .S(\datapath.idinstr_15_bF$buf50 ),
    .Y(_6372_)
);

MUX2X1 _17305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [4]),
    .B(\datapath.registers.1226[6] [4]),
    .S(\datapath.idinstr_15_bF$buf49 ),
    .Y(_6373_)
);

MUX2X1 _17306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6373_),
    .B(_6372_),
    .S(\datapath.idinstr_16_bF$buf0 ),
    .Y(_6374_)
);

NAND2X1 _17307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf23 ),
    .B(_6374_),
    .Y(_6375_)
);

MUX2X1 _17308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [4]),
    .B(\datapath.registers.1226[0] [4]),
    .S(\datapath.idinstr_15_bF$buf48 ),
    .Y(_6376_)
);

MUX2X1 _17309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [4]),
    .B(\datapath.registers.1226[2] [4]),
    .S(\datapath.idinstr_15_bF$buf47 ),
    .Y(_6377_)
);

MUX2X1 _17310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6377_),
    .B(_6376_),
    .S(\datapath.idinstr_16_bF$buf45 ),
    .Y(_6378_)
);

NAND2X1 _17311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf2),
    .B(_6378_),
    .Y(_6379_)
);

AOI21X1 _17312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6375_),
    .B(_6379_),
    .C(\datapath.idinstr_18_bF$buf2 ),
    .Y(_6380_)
);

OAI21X1 _17313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6380_),
    .B(_6371_),
    .C(_6140__bF$buf4),
    .Y(_6381_)
);

AOI21X1 _17314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6358_),
    .B(_6381_),
    .C(_6147__bF$buf0),
    .Y(\datapath.registers.rega_data [4])
);

MUX2X1 _17315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [5]),
    .B(\datapath.registers.1226[24] [5]),
    .S(\datapath.idinstr_15_bF$buf46 ),
    .Y(_6382_)
);

MUX2X1 _17316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [5]),
    .B(\datapath.registers.1226[26] [5]),
    .S(\datapath.idinstr_15_bF$buf45 ),
    .Y(_6383_)
);

MUX2X1 _17317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6383_),
    .B(_6382_),
    .S(\datapath.idinstr_16_bF$buf44 ),
    .Y(_6384_)
);

NAND2X1 _17318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf1),
    .B(_6384_),
    .Y(_6385_)
);

MUX2X1 _17319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [5]),
    .B(\datapath.registers.1226[28] [5]),
    .S(\datapath.idinstr_15_bF$buf44 ),
    .Y(_6386_)
);

MUX2X1 _17320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [5]),
    .B(\datapath.registers.1226[30] [5]),
    .S(\datapath.idinstr_15_bF$buf43 ),
    .Y(_6387_)
);

MUX2X1 _17321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6387_),
    .B(_6386_),
    .S(\datapath.idinstr_16_bF$buf43 ),
    .Y(_6388_)
);

NAND2X1 _17322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf22 ),
    .B(_6388_),
    .Y(_6389_)
);

AOI21X1 _17323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6385_),
    .B(_6389_),
    .C(_6145__bF$buf4),
    .Y(_6390_)
);

MUX2X1 _17324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [5]),
    .B(\datapath.registers.1226[16] [5]),
    .S(\datapath.idinstr_16_bF$buf42 ),
    .Y(_6391_)
);

NAND2X1 _17325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf8),
    .B(_6391_),
    .Y(_6392_)
);

MUX2X1 _17326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [5]),
    .B(\datapath.registers.1226[17] [5]),
    .S(\datapath.idinstr_16_bF$buf41 ),
    .Y(_6393_)
);

AOI21X1 _17327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf42 ),
    .B(_6393_),
    .C(\datapath.idinstr_17_bF$buf21 ),
    .Y(_6394_)
);

NAND2X1 _17328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6392_),
    .B(_6394_),
    .Y(_6395_)
);

MUX2X1 _17329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [5]),
    .B(\datapath.registers.1226[20] [5]),
    .S(\datapath.idinstr_16_bF$buf40 ),
    .Y(_6396_)
);

NAND2X1 _17330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf7),
    .B(_6396_),
    .Y(_6397_)
);

MUX2X1 _17331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [5]),
    .B(\datapath.registers.1226[21] [5]),
    .S(\datapath.idinstr_16_bF$buf39 ),
    .Y(_6398_)
);

AOI21X1 _17332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf41 ),
    .B(_6398_),
    .C(_6144__bF$buf0),
    .Y(_6399_)
);

NAND2X1 _17333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6397_),
    .B(_6399_),
    .Y(_6400_)
);

AOI21X1 _17334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6395_),
    .B(_6400_),
    .C(\datapath.idinstr_18_bF$buf1 ),
    .Y(_6401_)
);

OAI21X1 _17335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6390_),
    .B(_6401_),
    .C(\datapath.idinstr_19_bF$buf2 ),
    .Y(_6402_)
);

INVX1 _17336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [5]),
    .Y(_6403_)
);

AOI21X1 _17337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [5]),
    .B(\datapath.idinstr_17_bF$buf20 ),
    .C(_6141__bF$buf6),
    .Y(_6404_)
);

OAI21X1 _17338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf19 ),
    .B(_6403_),
    .C(_6404_),
    .Y(_6405_)
);

INVX1 _17339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [5]),
    .Y(_6406_)
);

AOI21X1 _17340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf18 ),
    .B(\datapath.registers.1226[12] [5]),
    .C(\datapath.idinstr_15_bF$buf40 ),
    .Y(_6407_)
);

OAI21X1 _17341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf17 ),
    .B(_6406_),
    .C(_6407_),
    .Y(_6408_)
);

NAND3X1 _17342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf1),
    .B(_6408_),
    .C(_6405_),
    .Y(_6409_)
);

INVX1 _17343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [5]),
    .Y(_6410_)
);

AOI21X1 _17344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [5]),
    .B(\datapath.idinstr_17_bF$buf16 ),
    .C(_6141__bF$buf5),
    .Y(_6411_)
);

OAI21X1 _17345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf15 ),
    .B(_6410_),
    .C(_6411_),
    .Y(_6412_)
);

INVX1 _17346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[10] [5]),
    .Y(_6413_)
);

AOI21X1 _17347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [5]),
    .B(\datapath.idinstr_17_bF$buf14 ),
    .C(\datapath.idinstr_15_bF$buf39 ),
    .Y(_6414_)
);

OAI21X1 _17348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf13 ),
    .B(_6413_),
    .C(_6414_),
    .Y(_6415_)
);

NAND3X1 _17349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_bF$buf38 ),
    .B(_6415_),
    .C(_6412_),
    .Y(_6416_)
);

AOI21X1 _17350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6409_),
    .B(_6416_),
    .C(_6145__bF$buf3),
    .Y(_6417_)
);

MUX2X1 _17351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [5]),
    .B(\datapath.registers.1226[0] [5]),
    .S(\datapath.idinstr_15_bF$buf38 ),
    .Y(_6418_)
);

MUX2X1 _17352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [5]),
    .B(\datapath.registers.1226[2] [5]),
    .S(\datapath.idinstr_15_bF$buf37 ),
    .Y(_6419_)
);

MUX2X1 _17353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6419_),
    .B(_6418_),
    .S(\datapath.idinstr_16_bF$buf37 ),
    .Y(_6420_)
);

NAND2X1 _17354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf10),
    .B(_6420_),
    .Y(_6421_)
);

MUX2X1 _17355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [5]),
    .B(\datapath.registers.1226[4] [5]),
    .S(\datapath.idinstr_15_bF$buf36 ),
    .Y(_6422_)
);

MUX2X1 _17356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [5]),
    .B(\datapath.registers.1226[6] [5]),
    .S(\datapath.idinstr_15_bF$buf35 ),
    .Y(_6423_)
);

MUX2X1 _17357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6423_),
    .B(_6422_),
    .S(\datapath.idinstr_16_bF$buf36 ),
    .Y(_6424_)
);

NAND2X1 _17358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf12 ),
    .B(_6424_),
    .Y(_6425_)
);

AOI21X1 _17359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6421_),
    .B(_6425_),
    .C(\datapath.idinstr_18_bF$buf0 ),
    .Y(_6426_)
);

OAI21X1 _17360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6426_),
    .B(_6417_),
    .C(_6140__bF$buf3),
    .Y(_6427_)
);

AOI21X1 _17361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6402_),
    .B(_6427_),
    .C(_6147__bF$buf4),
    .Y(\datapath.registers.rega_data [5])
);

MUX2X1 _17362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [6]),
    .B(\datapath.registers.1226[0] [6]),
    .S(\datapath.idinstr_15_bF$buf34 ),
    .Y(_6428_)
);

MUX2X1 _17363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [6]),
    .B(\datapath.registers.1226[2] [6]),
    .S(\datapath.idinstr_15_bF$buf33 ),
    .Y(_6429_)
);

MUX2X1 _17364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6429_),
    .B(_6428_),
    .S(\datapath.idinstr_16_bF$buf35 ),
    .Y(_6430_)
);

NAND2X1 _17365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf9),
    .B(_6430_),
    .Y(_6431_)
);

MUX2X1 _17366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [6]),
    .B(\datapath.registers.1226[4] [6]),
    .S(\datapath.idinstr_15_bF$buf32 ),
    .Y(_6432_)
);

MUX2X1 _17367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [6]),
    .B(\datapath.registers.1226[6] [6]),
    .S(\datapath.idinstr_15_bF$buf31 ),
    .Y(_6433_)
);

MUX2X1 _17368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6433_),
    .B(_6432_),
    .S(\datapath.idinstr_16_bF$buf34 ),
    .Y(_6434_)
);

NAND2X1 _17369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf11 ),
    .B(_6434_),
    .Y(_6435_)
);

AOI21X1 _17370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6431_),
    .B(_6435_),
    .C(\datapath.idinstr_18_bF$buf7 ),
    .Y(_6436_)
);

INVX1 _17371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [6]),
    .Y(_6437_)
);

AOI21X1 _17372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [6]),
    .B(\datapath.idinstr_17_bF$buf10 ),
    .C(_6141__bF$buf4),
    .Y(_6438_)
);

OAI21X1 _17373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf9 ),
    .B(_6437_),
    .C(_6438_),
    .Y(_6439_)
);

NAND2X1 _17374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [6]),
    .B(_6144__bF$buf8),
    .Y(_6440_)
);

AOI21X1 _17375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf8 ),
    .B(\datapath.registers.1226[12] [6]),
    .C(\datapath.idinstr_15_bF$buf30 ),
    .Y(_6441_)
);

AOI21X1 _17376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6441_),
    .B(_6440_),
    .C(\datapath.idinstr_16_bF$buf33 ),
    .Y(_6442_)
);

NAND2X1 _17377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6439_),
    .B(_6442_),
    .Y(_6443_)
);

INVX1 _17378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [6]),
    .Y(_6444_)
);

AOI21X1 _17379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [6]),
    .B(\datapath.idinstr_17_bF$buf7 ),
    .C(_6141__bF$buf3),
    .Y(_6445_)
);

OAI21X1 _17380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf6 ),
    .B(_6444_),
    .C(_6445_),
    .Y(_6446_)
);

INVX1 _17381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[10] [6]),
    .Y(_6447_)
);

AOI21X1 _17382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [6]),
    .B(\datapath.idinstr_17_bF$buf5 ),
    .C(\datapath.idinstr_15_bF$buf29 ),
    .Y(_6448_)
);

OAI21X1 _17383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf4 ),
    .B(_6447_),
    .C(_6448_),
    .Y(_6449_)
);

NAND3X1 _17384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_bF$buf32 ),
    .B(_6449_),
    .C(_6446_),
    .Y(_6450_)
);

AOI21X1 _17385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6443_),
    .B(_6450_),
    .C(_6145__bF$buf2),
    .Y(_6451_)
);

OAI21X1 _17386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6436_),
    .B(_6451_),
    .C(_6140__bF$buf2),
    .Y(_6452_)
);

MUX2X1 _17387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [6]),
    .B(\datapath.registers.1226[29] [6]),
    .S(\datapath.idinstr_16_bF$buf31 ),
    .Y(_6453_)
);

MUX2X1 _17388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [6]),
    .B(\datapath.registers.1226[28] [6]),
    .S(\datapath.idinstr_16_bF$buf30 ),
    .Y(_6454_)
);

MUX2X1 _17389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6454_),
    .B(_6453_),
    .S(_6141__bF$buf2),
    .Y(_6455_)
);

NAND2X1 _17390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf3 ),
    .B(_6455_),
    .Y(_6456_)
);

MUX2X1 _17391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [6]),
    .B(\datapath.registers.1226[25] [6]),
    .S(\datapath.idinstr_16_bF$buf29 ),
    .Y(_6457_)
);

MUX2X1 _17392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [6]),
    .B(\datapath.registers.1226[24] [6]),
    .S(\datapath.idinstr_16_bF$buf28 ),
    .Y(_6458_)
);

MUX2X1 _17393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6458_),
    .B(_6457_),
    .S(_6141__bF$buf1),
    .Y(_6459_)
);

NAND2X1 _17394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf7),
    .B(_6459_),
    .Y(_6460_)
);

AOI21X1 _17395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6456_),
    .B(_6460_),
    .C(_6145__bF$buf1),
    .Y(_6461_)
);

INVX1 _17396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [6]),
    .Y(_6462_)
);

AOI21X1 _17397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [6]),
    .B(\datapath.idinstr_17_bF$buf2 ),
    .C(_6141__bF$buf0),
    .Y(_6463_)
);

OAI21X1 _17398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6462_),
    .B(\datapath.idinstr_17_bF$buf1 ),
    .C(_6463_),
    .Y(_6464_)
);

INVX1 _17399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [6]),
    .Y(_6465_)
);

AOI21X1 _17400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [6]),
    .B(\datapath.idinstr_17_bF$buf0 ),
    .C(\datapath.idinstr_15_bF$buf28 ),
    .Y(_6466_)
);

OAI21X1 _17401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6465_),
    .B(\datapath.idinstr_17_bF$buf41 ),
    .C(_6466_),
    .Y(_6467_)
);

NAND3X1 _17402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_bF$buf27 ),
    .B(_6467_),
    .C(_6464_),
    .Y(_6468_)
);

INVX1 _17403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [6]),
    .Y(_6469_)
);

AOI21X1 _17404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [6]),
    .B(\datapath.idinstr_17_bF$buf40 ),
    .C(_6141__bF$buf10),
    .Y(_6470_)
);

OAI21X1 _17405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6469_),
    .B(\datapath.idinstr_17_bF$buf39 ),
    .C(_6470_),
    .Y(_6471_)
);

AOI21X1 _17406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [6]),
    .B(\datapath.idinstr_17_bF$buf38 ),
    .C(\datapath.idinstr_15_bF$buf27 ),
    .Y(_6472_)
);

OAI21X1 _17407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6002_),
    .B(\datapath.idinstr_17_bF$buf37 ),
    .C(_6472_),
    .Y(_6473_)
);

NAND3X1 _17408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf0),
    .B(_6473_),
    .C(_6471_),
    .Y(_6474_)
);

AOI21X1 _17409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6468_),
    .B(_6474_),
    .C(\datapath.idinstr_18_bF$buf6 ),
    .Y(_6475_)
);

OAI21X1 _17410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6461_),
    .B(_6475_),
    .C(\datapath.idinstr_19_bF$buf1 ),
    .Y(_6476_)
);

AOI21X1 _17411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6452_),
    .B(_6476_),
    .C(_6147__bF$buf3),
    .Y(\datapath.registers.rega_data [6])
);

MUX2X1 _17412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [7]),
    .B(\datapath.registers.1226[24] [7]),
    .S(\datapath.idinstr_15_bF$buf26 ),
    .Y(_6477_)
);

MUX2X1 _17413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [7]),
    .B(\datapath.registers.1226[26] [7]),
    .S(\datapath.idinstr_15_bF$buf25 ),
    .Y(_6478_)
);

MUX2X1 _17414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6478_),
    .B(_6477_),
    .S(\datapath.idinstr_16_bF$buf26 ),
    .Y(_6479_)
);

NAND2X1 _17415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf6),
    .B(_6479_),
    .Y(_6480_)
);

MUX2X1 _17416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [7]),
    .B(\datapath.registers.1226[28] [7]),
    .S(\datapath.idinstr_15_bF$buf24 ),
    .Y(_6481_)
);

MUX2X1 _17417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [7]),
    .B(\datapath.registers.1226[30] [7]),
    .S(\datapath.idinstr_15_bF$buf23 ),
    .Y(_6482_)
);

MUX2X1 _17418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6482_),
    .B(_6481_),
    .S(\datapath.idinstr_16_bF$buf25 ),
    .Y(_6483_)
);

NAND2X1 _17419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf36 ),
    .B(_6483_),
    .Y(_6484_)
);

AOI21X1 _17420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6480_),
    .B(_6484_),
    .C(_6145__bF$buf0),
    .Y(_6485_)
);

MUX2X1 _17421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [7]),
    .B(\datapath.registers.1226[16] [7]),
    .S(\datapath.idinstr_16_bF$buf24 ),
    .Y(_6486_)
);

NAND2X1 _17422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf9),
    .B(_6486_),
    .Y(_6487_)
);

MUX2X1 _17423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [7]),
    .B(\datapath.registers.1226[17] [7]),
    .S(\datapath.idinstr_16_bF$buf23 ),
    .Y(_6488_)
);

AOI21X1 _17424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf22 ),
    .B(_6488_),
    .C(\datapath.idinstr_17_bF$buf35 ),
    .Y(_6489_)
);

NAND2X1 _17425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6487_),
    .B(_6489_),
    .Y(_6490_)
);

MUX2X1 _17426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [7]),
    .B(\datapath.registers.1226[20] [7]),
    .S(\datapath.idinstr_16_bF$buf22 ),
    .Y(_6491_)
);

NAND2X1 _17427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf8),
    .B(_6491_),
    .Y(_6492_)
);

MUX2X1 _17428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [7]),
    .B(\datapath.registers.1226[21] [7]),
    .S(\datapath.idinstr_16_bF$buf21 ),
    .Y(_6493_)
);

AOI21X1 _17429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf21 ),
    .B(_6493_),
    .C(_6144__bF$buf5),
    .Y(_6494_)
);

NAND2X1 _17430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6492_),
    .B(_6494_),
    .Y(_6495_)
);

AOI21X1 _17431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6490_),
    .B(_6495_),
    .C(\datapath.idinstr_18_bF$buf5 ),
    .Y(_6496_)
);

OAI21X1 _17432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6485_),
    .B(_6496_),
    .C(\datapath.idinstr_19_bF$buf0 ),
    .Y(_6497_)
);

MUX2X1 _17433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [7]),
    .B(\datapath.registers.1226[8] [7]),
    .S(\datapath.idinstr_15_bF$buf20 ),
    .Y(_6498_)
);

MUX2X1 _17434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [7]),
    .B(\datapath.registers.1226[10] [7]),
    .S(\datapath.idinstr_15_bF$buf19 ),
    .Y(_6499_)
);

MUX2X1 _17435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6499_),
    .B(_6498_),
    .S(\datapath.idinstr_16_bF$buf20 ),
    .Y(_6500_)
);

NAND2X1 _17436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf4),
    .B(_6500_),
    .Y(_6501_)
);

AND2X2 _17437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [7]),
    .B(\datapath.idinstr_15_bF$buf18 ),
    .Y(_6502_)
);

INVX1 _17438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [7]),
    .Y(_6503_)
);

OAI21X1 _17439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6503_),
    .B(\datapath.idinstr_15_bF$buf17 ),
    .C(\datapath.idinstr_16_bF$buf19 ),
    .Y(_6504_)
);

NAND2X1 _17440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [7]),
    .B(_6141__bF$buf7),
    .Y(_6505_)
);

AOI21X1 _17441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [7]),
    .B(\datapath.idinstr_15_bF$buf16 ),
    .C(\datapath.idinstr_16_bF$buf18 ),
    .Y(_6506_)
);

AOI21X1 _17442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6506_),
    .B(_6505_),
    .C(_6144__bF$buf3),
    .Y(_6507_)
);

OAI21X1 _17443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6502_),
    .B(_6504_),
    .C(_6507_),
    .Y(_6508_)
);

AOI21X1 _17444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6508_),
    .B(_6501_),
    .C(_6145__bF$buf7),
    .Y(_6509_)
);

MUX2X1 _17445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [7]),
    .B(\datapath.registers.1226[4] [7]),
    .S(\datapath.idinstr_15_bF$buf15 ),
    .Y(_6510_)
);

MUX2X1 _17446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [7]),
    .B(\datapath.registers.1226[6] [7]),
    .S(\datapath.idinstr_15_bF$buf14 ),
    .Y(_6511_)
);

MUX2X1 _17447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6511_),
    .B(_6510_),
    .S(\datapath.idinstr_16_bF$buf17 ),
    .Y(_6512_)
);

NAND2X1 _17448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf34 ),
    .B(_6512_),
    .Y(_6513_)
);

MUX2X1 _17449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [7]),
    .B(\datapath.registers.1226[0] [7]),
    .S(\datapath.idinstr_15_bF$buf13 ),
    .Y(_6514_)
);

MUX2X1 _17450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [7]),
    .B(\datapath.registers.1226[2] [7]),
    .S(\datapath.idinstr_15_bF$buf12 ),
    .Y(_6515_)
);

MUX2X1 _17451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6515_),
    .B(_6514_),
    .S(\datapath.idinstr_16_bF$buf16 ),
    .Y(_6516_)
);

NAND2X1 _17452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf2),
    .B(_6516_),
    .Y(_6517_)
);

AOI21X1 _17453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6513_),
    .B(_6517_),
    .C(\datapath.idinstr_18_bF$buf4 ),
    .Y(_6518_)
);

OAI21X1 _17454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6518_),
    .B(_6509_),
    .C(_6140__bF$buf1),
    .Y(_6519_)
);

AOI21X1 _17455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6497_),
    .B(_6519_),
    .C(_6147__bF$buf2),
    .Y(\datapath.registers.rega_data [7])
);

MUX2X1 _17456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [8]),
    .B(\datapath.registers.1226[8] [8]),
    .S(\datapath.idinstr_15_bF$buf11 ),
    .Y(_6520_)
);

MUX2X1 _17457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [8]),
    .B(\datapath.registers.1226[10] [8]),
    .S(\datapath.idinstr_15_bF$buf10 ),
    .Y(_6521_)
);

MUX2X1 _17458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6521_),
    .B(_6520_),
    .S(\datapath.idinstr_16_bF$buf15 ),
    .Y(_6522_)
);

NAND2X1 _17459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf1),
    .B(_6522_),
    .Y(_6523_)
);

AND2X2 _17460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [8]),
    .B(\datapath.idinstr_15_bF$buf9 ),
    .Y(_6524_)
);

INVX1 _17461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [8]),
    .Y(_6525_)
);

OAI21X1 _17462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6525_),
    .B(\datapath.idinstr_15_bF$buf8 ),
    .C(\datapath.idinstr_16_bF$buf14 ),
    .Y(_6526_)
);

NAND2X1 _17463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [8]),
    .B(_6141__bF$buf6),
    .Y(_6527_)
);

AOI21X1 _17464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [8]),
    .B(\datapath.idinstr_15_bF$buf7 ),
    .C(\datapath.idinstr_16_bF$buf13 ),
    .Y(_6528_)
);

AOI21X1 _17465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6528_),
    .B(_6527_),
    .C(_6144__bF$buf0),
    .Y(_6529_)
);

OAI21X1 _17466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6524_),
    .B(_6526_),
    .C(_6529_),
    .Y(_6530_)
);

AOI21X1 _17467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6530_),
    .B(_6523_),
    .C(_6145__bF$buf6),
    .Y(_6531_)
);

MUX2X1 _17468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [8]),
    .B(\datapath.registers.1226[4] [8]),
    .S(\datapath.idinstr_15_bF$buf6 ),
    .Y(_6532_)
);

MUX2X1 _17469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [8]),
    .B(\datapath.registers.1226[6] [8]),
    .S(\datapath.idinstr_15_bF$buf5 ),
    .Y(_6533_)
);

MUX2X1 _17470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6533_),
    .B(_6532_),
    .S(\datapath.idinstr_16_bF$buf12 ),
    .Y(_6534_)
);

NAND2X1 _17471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf33 ),
    .B(_6534_),
    .Y(_6535_)
);

MUX2X1 _17472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [8]),
    .B(\datapath.registers.1226[0] [8]),
    .S(\datapath.idinstr_15_bF$buf4 ),
    .Y(_6536_)
);

MUX2X1 _17473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [8]),
    .B(\datapath.registers.1226[2] [8]),
    .S(\datapath.idinstr_15_bF$buf3 ),
    .Y(_6537_)
);

MUX2X1 _17474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6537_),
    .B(_6536_),
    .S(\datapath.idinstr_16_bF$buf11 ),
    .Y(_6538_)
);

NAND2X1 _17475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf10),
    .B(_6538_),
    .Y(_6539_)
);

AOI21X1 _17476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6535_),
    .B(_6539_),
    .C(\datapath.idinstr_18_bF$buf3 ),
    .Y(_6540_)
);

OAI21X1 _17477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6540_),
    .B(_6531_),
    .C(_6140__bF$buf0),
    .Y(_6541_)
);

INVX1 _17478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [8]),
    .Y(_6542_)
);

AOI21X1 _17479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [8]),
    .B(\datapath.idinstr_17_bF$buf32 ),
    .C(_6141__bF$buf5),
    .Y(_6543_)
);

OAI21X1 _17480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6542_),
    .B(\datapath.idinstr_17_bF$buf31 ),
    .C(_6543_),
    .Y(_6544_)
);

NAND2X1 _17481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [8]),
    .B(_6144__bF$buf9),
    .Y(_6545_)
);

AOI21X1 _17482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [8]),
    .B(\datapath.idinstr_17_bF$buf30 ),
    .C(\datapath.idinstr_15_bF$buf2 ),
    .Y(_6546_)
);

AOI21X1 _17483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6546_),
    .B(_6545_),
    .C(_6143__bF$buf4),
    .Y(_6547_)
);

NAND2X1 _17484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6544_),
    .B(_6547_),
    .Y(_6548_)
);

INVX1 _17485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [8]),
    .Y(_6549_)
);

AOI21X1 _17486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [8]),
    .B(\datapath.idinstr_17_bF$buf29 ),
    .C(_6141__bF$buf4),
    .Y(_6550_)
);

OAI21X1 _17487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6549_),
    .B(\datapath.idinstr_17_bF$buf28 ),
    .C(_6550_),
    .Y(_6551_)
);

AOI21X1 _17488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [8]),
    .B(\datapath.idinstr_17_bF$buf27 ),
    .C(\datapath.idinstr_15_bF$buf1 ),
    .Y(_6552_)
);

OAI21X1 _17489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6006_),
    .B(\datapath.idinstr_17_bF$buf26 ),
    .C(_6552_),
    .Y(_6553_)
);

NAND3X1 _17490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf3),
    .B(_6553_),
    .C(_6551_),
    .Y(_6554_)
);

AOI21X1 _17491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6548_),
    .B(_6554_),
    .C(\datapath.idinstr_18_bF$buf2 ),
    .Y(_6555_)
);

MUX2X1 _17492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [8]),
    .B(\datapath.registers.1226[29] [8]),
    .S(\datapath.idinstr_16_bF$buf10 ),
    .Y(_6556_)
);

MUX2X1 _17493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [8]),
    .B(\datapath.registers.1226[28] [8]),
    .S(\datapath.idinstr_16_bF$buf9 ),
    .Y(_6557_)
);

MUX2X1 _17494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6557_),
    .B(_6556_),
    .S(_6141__bF$buf3),
    .Y(_6558_)
);

NAND2X1 _17495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf25 ),
    .B(_6558_),
    .Y(_6559_)
);

MUX2X1 _17496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [8]),
    .B(\datapath.registers.1226[25] [8]),
    .S(\datapath.idinstr_16_bF$buf8 ),
    .Y(_6560_)
);

MUX2X1 _17497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [8]),
    .B(\datapath.registers.1226[24] [8]),
    .S(\datapath.idinstr_16_bF$buf7 ),
    .Y(_6561_)
);

MUX2X1 _17498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6561_),
    .B(_6560_),
    .S(_6141__bF$buf2),
    .Y(_6562_)
);

NAND2X1 _17499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf8),
    .B(_6562_),
    .Y(_6563_)
);

AOI21X1 _17500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6559_),
    .B(_6563_),
    .C(_6145__bF$buf5),
    .Y(_6564_)
);

OAI21X1 _17501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6564_),
    .B(_6555_),
    .C(\datapath.idinstr_19_bF$buf5 ),
    .Y(_6565_)
);

AOI21X1 _17502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6565_),
    .B(_6541_),
    .C(_6147__bF$buf1),
    .Y(\datapath.registers.rega_data [8])
);

MUX2X1 _17503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [9]),
    .B(\datapath.registers.1226[24] [9]),
    .S(\datapath.idinstr_15_bF$buf0 ),
    .Y(_6566_)
);

MUX2X1 _17504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [9]),
    .B(\datapath.registers.1226[26] [9]),
    .S(\datapath.idinstr_15_bF$buf53 ),
    .Y(_6567_)
);

MUX2X1 _17505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6567_),
    .B(_6566_),
    .S(\datapath.idinstr_16_bF$buf6 ),
    .Y(_6568_)
);

NAND2X1 _17506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf7),
    .B(_6568_),
    .Y(_6569_)
);

MUX2X1 _17507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [9]),
    .B(\datapath.registers.1226[28] [9]),
    .S(\datapath.idinstr_15_bF$buf52 ),
    .Y(_6570_)
);

MUX2X1 _17508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [9]),
    .B(\datapath.registers.1226[30] [9]),
    .S(\datapath.idinstr_15_bF$buf51 ),
    .Y(_6571_)
);

MUX2X1 _17509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6571_),
    .B(_6570_),
    .S(\datapath.idinstr_16_bF$buf5 ),
    .Y(_6572_)
);

NAND2X1 _17510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf24 ),
    .B(_6572_),
    .Y(_6573_)
);

AOI21X1 _17511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6569_),
    .B(_6573_),
    .C(_6145__bF$buf4),
    .Y(_6574_)
);

MUX2X1 _17512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [9]),
    .B(\datapath.registers.1226[16] [9]),
    .S(\datapath.idinstr_16_bF$buf4 ),
    .Y(_6575_)
);

NAND2X1 _17513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf1),
    .B(_6575_),
    .Y(_6576_)
);

MUX2X1 _17514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [9]),
    .B(\datapath.registers.1226[17] [9]),
    .S(\datapath.idinstr_16_bF$buf3 ),
    .Y(_6577_)
);

AOI21X1 _17515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf50 ),
    .B(_6577_),
    .C(\datapath.idinstr_17_bF$buf23 ),
    .Y(_6578_)
);

NAND2X1 _17516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6576_),
    .B(_6578_),
    .Y(_6579_)
);

MUX2X1 _17517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [9]),
    .B(\datapath.registers.1226[20] [9]),
    .S(\datapath.idinstr_16_bF$buf2 ),
    .Y(_6580_)
);

NAND2X1 _17518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf0),
    .B(_6580_),
    .Y(_6581_)
);

MUX2X1 _17519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [9]),
    .B(\datapath.registers.1226[21] [9]),
    .S(\datapath.idinstr_16_bF$buf1 ),
    .Y(_6582_)
);

AOI21X1 _17520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf49 ),
    .B(_6582_),
    .C(_6144__bF$buf6),
    .Y(_6583_)
);

NAND2X1 _17521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6581_),
    .B(_6583_),
    .Y(_6584_)
);

AOI21X1 _17522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6579_),
    .B(_6584_),
    .C(\datapath.idinstr_18_bF$buf1 ),
    .Y(_6585_)
);

OAI21X1 _17523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6574_),
    .B(_6585_),
    .C(\datapath.idinstr_19_bF$buf4 ),
    .Y(_6586_)
);

MUX2X1 _17524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [9]),
    .B(\datapath.registers.1226[8] [9]),
    .S(\datapath.idinstr_15_bF$buf48 ),
    .Y(_6587_)
);

MUX2X1 _17525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [9]),
    .B(\datapath.registers.1226[10] [9]),
    .S(\datapath.idinstr_15_bF$buf47 ),
    .Y(_6588_)
);

MUX2X1 _17526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6588_),
    .B(_6587_),
    .S(\datapath.idinstr_16_bF$buf0 ),
    .Y(_6589_)
);

NAND2X1 _17527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf5),
    .B(_6589_),
    .Y(_6590_)
);

INVX1 _17528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [9]),
    .Y(_6591_)
);

NOR2X1 _17529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6591_),
    .B(_6141__bF$buf10),
    .Y(_6592_)
);

INVX1 _17530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [9]),
    .Y(_6593_)
);

OAI21X1 _17531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6593_),
    .B(\datapath.idinstr_15_bF$buf46 ),
    .C(\datapath.idinstr_16_bF$buf45 ),
    .Y(_6594_)
);

NAND2X1 _17532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [9]),
    .B(_6141__bF$buf9),
    .Y(_6595_)
);

AOI21X1 _17533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [9]),
    .B(\datapath.idinstr_15_bF$buf45 ),
    .C(\datapath.idinstr_16_bF$buf44 ),
    .Y(_6596_)
);

AOI21X1 _17534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6596_),
    .B(_6595_),
    .C(_6144__bF$buf4),
    .Y(_6597_)
);

OAI21X1 _17535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6592_),
    .B(_6594_),
    .C(_6597_),
    .Y(_6598_)
);

AOI21X1 _17536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6598_),
    .B(_6590_),
    .C(_6145__bF$buf3),
    .Y(_6599_)
);

MUX2X1 _17537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [9]),
    .B(\datapath.registers.1226[4] [9]),
    .S(\datapath.idinstr_15_bF$buf44 ),
    .Y(_6600_)
);

MUX2X1 _17538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [9]),
    .B(\datapath.registers.1226[6] [9]),
    .S(\datapath.idinstr_15_bF$buf43 ),
    .Y(_6601_)
);

MUX2X1 _17539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6601_),
    .B(_6600_),
    .S(\datapath.idinstr_16_bF$buf43 ),
    .Y(_6602_)
);

NAND2X1 _17540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf22 ),
    .B(_6602_),
    .Y(_6603_)
);

MUX2X1 _17541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [9]),
    .B(\datapath.registers.1226[0] [9]),
    .S(\datapath.idinstr_15_bF$buf42 ),
    .Y(_6604_)
);

MUX2X1 _17542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [9]),
    .B(\datapath.registers.1226[2] [9]),
    .S(\datapath.idinstr_15_bF$buf41 ),
    .Y(_6605_)
);

MUX2X1 _17543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6605_),
    .B(_6604_),
    .S(\datapath.idinstr_16_bF$buf42 ),
    .Y(_6606_)
);

NAND2X1 _17544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf3),
    .B(_6606_),
    .Y(_6607_)
);

AOI21X1 _17545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6603_),
    .B(_6607_),
    .C(\datapath.idinstr_18_bF$buf0 ),
    .Y(_6608_)
);

OAI21X1 _17546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6608_),
    .B(_6599_),
    .C(_6140__bF$buf4),
    .Y(_6609_)
);

AOI21X1 _17547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6586_),
    .B(_6609_),
    .C(_6147__bF$buf0),
    .Y(\datapath.registers.rega_data [9])
);

MUX2X1 _17548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [10]),
    .B(\datapath.registers.1226[8] [10]),
    .S(\datapath.idinstr_15_bF$buf40 ),
    .Y(_6610_)
);

MUX2X1 _17549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [10]),
    .B(\datapath.registers.1226[10] [10]),
    .S(\datapath.idinstr_15_bF$buf39 ),
    .Y(_6611_)
);

MUX2X1 _17550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6611_),
    .B(_6610_),
    .S(\datapath.idinstr_16_bF$buf41 ),
    .Y(_6612_)
);

NAND2X1 _17551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf2),
    .B(_6612_),
    .Y(_6613_)
);

INVX1 _17552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [10]),
    .Y(_6614_)
);

NOR2X1 _17553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6614_),
    .B(_6141__bF$buf8),
    .Y(_6615_)
);

INVX1 _17554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [10]),
    .Y(_6616_)
);

OAI21X1 _17555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6616_),
    .B(\datapath.idinstr_15_bF$buf38 ),
    .C(\datapath.idinstr_16_bF$buf40 ),
    .Y(_6617_)
);

NAND2X1 _17556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [10]),
    .B(_6141__bF$buf7),
    .Y(_6618_)
);

AOI21X1 _17557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [10]),
    .B(\datapath.idinstr_15_bF$buf37 ),
    .C(\datapath.idinstr_16_bF$buf39 ),
    .Y(_6619_)
);

AOI21X1 _17558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6619_),
    .B(_6618_),
    .C(_6144__bF$buf1),
    .Y(_6620_)
);

OAI21X1 _17559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6615_),
    .B(_6617_),
    .C(_6620_),
    .Y(_6621_)
);

AOI21X1 _17560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6621_),
    .B(_6613_),
    .C(_6145__bF$buf2),
    .Y(_6622_)
);

MUX2X1 _17561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [10]),
    .B(\datapath.registers.1226[4] [10]),
    .S(\datapath.idinstr_15_bF$buf36 ),
    .Y(_6623_)
);

MUX2X1 _17562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [10]),
    .B(\datapath.registers.1226[6] [10]),
    .S(\datapath.idinstr_15_bF$buf35 ),
    .Y(_6624_)
);

MUX2X1 _17563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6624_),
    .B(_6623_),
    .S(\datapath.idinstr_16_bF$buf38 ),
    .Y(_6625_)
);

NAND2X1 _17564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf21 ),
    .B(_6625_),
    .Y(_6626_)
);

MUX2X1 _17565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [10]),
    .B(\datapath.registers.1226[0] [10]),
    .S(\datapath.idinstr_15_bF$buf34 ),
    .Y(_6627_)
);

MUX2X1 _17566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [10]),
    .B(\datapath.registers.1226[2] [10]),
    .S(\datapath.idinstr_15_bF$buf33 ),
    .Y(_6628_)
);

MUX2X1 _17567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6628_),
    .B(_6627_),
    .S(\datapath.idinstr_16_bF$buf37 ),
    .Y(_6629_)
);

NAND2X1 _17568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf0),
    .B(_6629_),
    .Y(_6630_)
);

AOI21X1 _17569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6626_),
    .B(_6630_),
    .C(\datapath.idinstr_18_bF$buf7 ),
    .Y(_6631_)
);

OAI21X1 _17570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6631_),
    .B(_6622_),
    .C(_6140__bF$buf3),
    .Y(_6632_)
);

INVX1 _17571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [10]),
    .Y(_6633_)
);

AOI21X1 _17572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [10]),
    .B(\datapath.idinstr_17_bF$buf20 ),
    .C(_6141__bF$buf6),
    .Y(_6634_)
);

OAI21X1 _17573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6633_),
    .B(\datapath.idinstr_17_bF$buf19 ),
    .C(_6634_),
    .Y(_6635_)
);

NAND2X1 _17574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [10]),
    .B(_6144__bF$buf10),
    .Y(_6636_)
);

AOI21X1 _17575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [10]),
    .B(\datapath.idinstr_17_bF$buf18 ),
    .C(\datapath.idinstr_15_bF$buf32 ),
    .Y(_6637_)
);

AOI21X1 _17576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6637_),
    .B(_6636_),
    .C(_6143__bF$buf2),
    .Y(_6638_)
);

NAND2X1 _17577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6635_),
    .B(_6638_),
    .Y(_6639_)
);

INVX1 _17578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [10]),
    .Y(_6640_)
);

AOI21X1 _17579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [10]),
    .B(\datapath.idinstr_17_bF$buf17 ),
    .C(_6141__bF$buf5),
    .Y(_6641_)
);

OAI21X1 _17580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6640_),
    .B(\datapath.idinstr_17_bF$buf16 ),
    .C(_6641_),
    .Y(_6642_)
);

AOI21X1 _17581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [10]),
    .B(\datapath.idinstr_17_bF$buf15 ),
    .C(\datapath.idinstr_15_bF$buf31 ),
    .Y(_6643_)
);

OAI21X1 _17582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6009_),
    .B(\datapath.idinstr_17_bF$buf14 ),
    .C(_6643_),
    .Y(_6644_)
);

NAND3X1 _17583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf1),
    .B(_6644_),
    .C(_6642_),
    .Y(_6645_)
);

AOI21X1 _17584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6639_),
    .B(_6645_),
    .C(\datapath.idinstr_18_bF$buf6 ),
    .Y(_6646_)
);

MUX2X1 _17585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [10]),
    .B(\datapath.registers.1226[29] [10]),
    .S(\datapath.idinstr_16_bF$buf36 ),
    .Y(_6647_)
);

MUX2X1 _17586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [10]),
    .B(\datapath.registers.1226[28] [10]),
    .S(\datapath.idinstr_16_bF$buf35 ),
    .Y(_6648_)
);

MUX2X1 _17587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6648_),
    .B(_6647_),
    .S(_6141__bF$buf4),
    .Y(_6649_)
);

NAND2X1 _17588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf13 ),
    .B(_6649_),
    .Y(_6650_)
);

MUX2X1 _17589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [10]),
    .B(\datapath.registers.1226[25] [10]),
    .S(\datapath.idinstr_16_bF$buf34 ),
    .Y(_6651_)
);

MUX2X1 _17590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [10]),
    .B(\datapath.registers.1226[24] [10]),
    .S(\datapath.idinstr_16_bF$buf33 ),
    .Y(_6652_)
);

MUX2X1 _17591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6652_),
    .B(_6651_),
    .S(_6141__bF$buf3),
    .Y(_6653_)
);

NAND2X1 _17592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf9),
    .B(_6653_),
    .Y(_6654_)
);

AOI21X1 _17593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6650_),
    .B(_6654_),
    .C(_6145__bF$buf1),
    .Y(_6655_)
);

OAI21X1 _17594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6655_),
    .B(_6646_),
    .C(\datapath.idinstr_19_bF$buf3 ),
    .Y(_6656_)
);

AOI21X1 _17595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6656_),
    .B(_6632_),
    .C(_6147__bF$buf4),
    .Y(\datapath.registers.rega_data [10])
);

MUX2X1 _17596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [11]),
    .B(\datapath.registers.1226[24] [11]),
    .S(\datapath.idinstr_15_bF$buf30 ),
    .Y(_6657_)
);

MUX2X1 _17597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [11]),
    .B(\datapath.registers.1226[26] [11]),
    .S(\datapath.idinstr_15_bF$buf29 ),
    .Y(_6658_)
);

MUX2X1 _17598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6658_),
    .B(_6657_),
    .S(\datapath.idinstr_16_bF$buf32 ),
    .Y(_6659_)
);

NAND2X1 _17599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf8),
    .B(_6659_),
    .Y(_6660_)
);

MUX2X1 _17600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [11]),
    .B(\datapath.registers.1226[28] [11]),
    .S(\datapath.idinstr_15_bF$buf28 ),
    .Y(_6661_)
);

MUX2X1 _17601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [11]),
    .B(\datapath.registers.1226[30] [11]),
    .S(\datapath.idinstr_15_bF$buf27 ),
    .Y(_6662_)
);

MUX2X1 _17602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6662_),
    .B(_6661_),
    .S(\datapath.idinstr_16_bF$buf31 ),
    .Y(_6663_)
);

NAND2X1 _17603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf12 ),
    .B(_6663_),
    .Y(_6664_)
);

AOI21X1 _17604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6660_),
    .B(_6664_),
    .C(_6145__bF$buf0),
    .Y(_6665_)
);

MUX2X1 _17605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [11]),
    .B(\datapath.registers.1226[16] [11]),
    .S(\datapath.idinstr_16_bF$buf30 ),
    .Y(_6666_)
);

NAND2X1 _17606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf2),
    .B(_6666_),
    .Y(_6667_)
);

MUX2X1 _17607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [11]),
    .B(\datapath.registers.1226[17] [11]),
    .S(\datapath.idinstr_16_bF$buf29 ),
    .Y(_6668_)
);

AOI21X1 _17608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf26 ),
    .B(_6668_),
    .C(\datapath.idinstr_17_bF$buf11 ),
    .Y(_6669_)
);

NAND2X1 _17609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6667_),
    .B(_6669_),
    .Y(_6670_)
);

MUX2X1 _17610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [11]),
    .B(\datapath.registers.1226[20] [11]),
    .S(\datapath.idinstr_16_bF$buf28 ),
    .Y(_6671_)
);

NAND2X1 _17611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf1),
    .B(_6671_),
    .Y(_6672_)
);

MUX2X1 _17612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [11]),
    .B(\datapath.registers.1226[21] [11]),
    .S(\datapath.idinstr_16_bF$buf27 ),
    .Y(_6673_)
);

AOI21X1 _17613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf25 ),
    .B(_6673_),
    .C(_6144__bF$buf7),
    .Y(_6674_)
);

NAND2X1 _17614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6672_),
    .B(_6674_),
    .Y(_6675_)
);

AOI21X1 _17615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6670_),
    .B(_6675_),
    .C(\datapath.idinstr_18_bF$buf5 ),
    .Y(_6676_)
);

OAI21X1 _17616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6665_),
    .B(_6676_),
    .C(\datapath.idinstr_19_bF$buf2 ),
    .Y(_6677_)
);

MUX2X1 _17617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [11]),
    .B(\datapath.registers.1226[8] [11]),
    .S(\datapath.idinstr_15_bF$buf24 ),
    .Y(_6678_)
);

MUX2X1 _17618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [11]),
    .B(\datapath.registers.1226[10] [11]),
    .S(\datapath.idinstr_15_bF$buf23 ),
    .Y(_6679_)
);

MUX2X1 _17619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6679_),
    .B(_6678_),
    .S(\datapath.idinstr_16_bF$buf26 ),
    .Y(_6680_)
);

NAND2X1 _17620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf6),
    .B(_6680_),
    .Y(_6681_)
);

AND2X2 _17621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [11]),
    .B(\datapath.idinstr_15_bF$buf22 ),
    .Y(_6682_)
);

INVX1 _17622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [11]),
    .Y(_6683_)
);

OAI21X1 _17623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6683_),
    .B(\datapath.idinstr_15_bF$buf21 ),
    .C(\datapath.idinstr_16_bF$buf25 ),
    .Y(_6684_)
);

NAND2X1 _17624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [11]),
    .B(_6141__bF$buf0),
    .Y(_6685_)
);

AOI21X1 _17625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [11]),
    .B(\datapath.idinstr_15_bF$buf20 ),
    .C(\datapath.idinstr_16_bF$buf24 ),
    .Y(_6686_)
);

AOI21X1 _17626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6686_),
    .B(_6685_),
    .C(_6144__bF$buf5),
    .Y(_6687_)
);

OAI21X1 _17627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6682_),
    .B(_6684_),
    .C(_6687_),
    .Y(_6688_)
);

AOI21X1 _17628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6688_),
    .B(_6681_),
    .C(_6145__bF$buf7),
    .Y(_6689_)
);

MUX2X1 _17629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [11]),
    .B(\datapath.registers.1226[4] [11]),
    .S(\datapath.idinstr_15_bF$buf19 ),
    .Y(_6690_)
);

MUX2X1 _17630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [11]),
    .B(\datapath.registers.1226[6] [11]),
    .S(\datapath.idinstr_15_bF$buf18 ),
    .Y(_6691_)
);

MUX2X1 _17631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6691_),
    .B(_6690_),
    .S(\datapath.idinstr_16_bF$buf23 ),
    .Y(_6692_)
);

NAND2X1 _17632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf10 ),
    .B(_6692_),
    .Y(_6693_)
);

MUX2X1 _17633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [11]),
    .B(\datapath.registers.1226[0] [11]),
    .S(\datapath.idinstr_15_bF$buf17 ),
    .Y(_6694_)
);

MUX2X1 _17634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [11]),
    .B(\datapath.registers.1226[2] [11]),
    .S(\datapath.idinstr_15_bF$buf16 ),
    .Y(_6695_)
);

MUX2X1 _17635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6695_),
    .B(_6694_),
    .S(\datapath.idinstr_16_bF$buf22 ),
    .Y(_6696_)
);

NAND2X1 _17636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf4),
    .B(_6696_),
    .Y(_6697_)
);

AOI21X1 _17637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6693_),
    .B(_6697_),
    .C(\datapath.idinstr_18_bF$buf4 ),
    .Y(_6698_)
);

OAI21X1 _17638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6698_),
    .B(_6689_),
    .C(_6140__bF$buf2),
    .Y(_6699_)
);

AOI21X1 _17639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6677_),
    .B(_6699_),
    .C(_6147__bF$buf3),
    .Y(\datapath.registers.rega_data [11])
);

MUX2X1 _17640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [12]),
    .B(\datapath.registers.1226[24] [12]),
    .S(\datapath.idinstr_15_bF$buf15 ),
    .Y(_6700_)
);

MUX2X1 _17641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [12]),
    .B(\datapath.registers.1226[26] [12]),
    .S(\datapath.idinstr_15_bF$buf14 ),
    .Y(_6701_)
);

MUX2X1 _17642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6701_),
    .B(_6700_),
    .S(\datapath.idinstr_16_bF$buf21 ),
    .Y(_6702_)
);

NAND2X1 _17643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf3),
    .B(_6702_),
    .Y(_6703_)
);

MUX2X1 _17644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [12]),
    .B(\datapath.registers.1226[28] [12]),
    .S(\datapath.idinstr_15_bF$buf13 ),
    .Y(_6704_)
);

MUX2X1 _17645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [12]),
    .B(\datapath.registers.1226[30] [12]),
    .S(\datapath.idinstr_15_bF$buf12 ),
    .Y(_6705_)
);

MUX2X1 _17646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6705_),
    .B(_6704_),
    .S(\datapath.idinstr_16_bF$buf20 ),
    .Y(_6706_)
);

NAND2X1 _17647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf9 ),
    .B(_6706_),
    .Y(_6707_)
);

AOI21X1 _17648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6703_),
    .B(_6707_),
    .C(_6145__bF$buf6),
    .Y(_6708_)
);

MUX2X1 _17649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [12]),
    .B(\datapath.registers.1226[16] [12]),
    .S(\datapath.idinstr_16_bF$buf19 ),
    .Y(_6709_)
);

NAND2X1 _17650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf10),
    .B(_6709_),
    .Y(_6710_)
);

MUX2X1 _17651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [12]),
    .B(\datapath.registers.1226[17] [12]),
    .S(\datapath.idinstr_16_bF$buf18 ),
    .Y(_6711_)
);

AOI21X1 _17652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf11 ),
    .B(_6711_),
    .C(\datapath.idinstr_17_bF$buf8 ),
    .Y(_6712_)
);

NAND2X1 _17653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6710_),
    .B(_6712_),
    .Y(_6713_)
);

MUX2X1 _17654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [12]),
    .B(\datapath.registers.1226[20] [12]),
    .S(\datapath.idinstr_16_bF$buf17 ),
    .Y(_6714_)
);

NAND2X1 _17655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf9),
    .B(_6714_),
    .Y(_6715_)
);

MUX2X1 _17656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [12]),
    .B(\datapath.registers.1226[21] [12]),
    .S(\datapath.idinstr_16_bF$buf16 ),
    .Y(_6716_)
);

AOI21X1 _17657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf10 ),
    .B(_6716_),
    .C(_6144__bF$buf2),
    .Y(_6717_)
);

NAND2X1 _17658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6715_),
    .B(_6717_),
    .Y(_6718_)
);

AOI21X1 _17659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6713_),
    .B(_6718_),
    .C(\datapath.idinstr_18_bF$buf3 ),
    .Y(_6719_)
);

OAI21X1 _17660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6708_),
    .B(_6719_),
    .C(\datapath.idinstr_19_bF$buf1 ),
    .Y(_6720_)
);

INVX1 _17661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [12]),
    .Y(_6721_)
);

AOI21X1 _17662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [12]),
    .B(\datapath.idinstr_17_bF$buf7 ),
    .C(_6141__bF$buf8),
    .Y(_6722_)
);

OAI21X1 _17663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf6 ),
    .B(_6721_),
    .C(_6722_),
    .Y(_6723_)
);

INVX1 _17664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [12]),
    .Y(_6724_)
);

AOI21X1 _17665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf5 ),
    .B(\datapath.registers.1226[12] [12]),
    .C(\datapath.idinstr_15_bF$buf9 ),
    .Y(_6725_)
);

OAI21X1 _17666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf4 ),
    .B(_6724_),
    .C(_6725_),
    .Y(_6726_)
);

NAND3X1 _17667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf0),
    .B(_6726_),
    .C(_6723_),
    .Y(_6727_)
);

INVX1 _17668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [12]),
    .Y(_6728_)
);

AOI21X1 _17669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [12]),
    .B(\datapath.idinstr_17_bF$buf3 ),
    .C(_6141__bF$buf7),
    .Y(_6729_)
);

OAI21X1 _17670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf2 ),
    .B(_6728_),
    .C(_6729_),
    .Y(_6730_)
);

INVX1 _17671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[10] [12]),
    .Y(_6731_)
);

AOI21X1 _17672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [12]),
    .B(\datapath.idinstr_17_bF$buf1 ),
    .C(\datapath.idinstr_15_bF$buf8 ),
    .Y(_6732_)
);

OAI21X1 _17673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf0 ),
    .B(_6731_),
    .C(_6732_),
    .Y(_6733_)
);

NAND3X1 _17674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_bF$buf15 ),
    .B(_6733_),
    .C(_6730_),
    .Y(_6734_)
);

AOI21X1 _17675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6727_),
    .B(_6734_),
    .C(_6145__bF$buf5),
    .Y(_6735_)
);

MUX2X1 _17676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [12]),
    .B(\datapath.registers.1226[0] [12]),
    .S(\datapath.idinstr_15_bF$buf7 ),
    .Y(_6736_)
);

MUX2X1 _17677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [12]),
    .B(\datapath.registers.1226[2] [12]),
    .S(\datapath.idinstr_15_bF$buf6 ),
    .Y(_6737_)
);

MUX2X1 _17678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6737_),
    .B(_6736_),
    .S(\datapath.idinstr_16_bF$buf14 ),
    .Y(_6738_)
);

NAND2X1 _17679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf1),
    .B(_6738_),
    .Y(_6739_)
);

MUX2X1 _17680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [12]),
    .B(\datapath.registers.1226[4] [12]),
    .S(\datapath.idinstr_15_bF$buf5 ),
    .Y(_6740_)
);

MUX2X1 _17681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [12]),
    .B(\datapath.registers.1226[6] [12]),
    .S(\datapath.idinstr_15_bF$buf4 ),
    .Y(_6741_)
);

MUX2X1 _17682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6741_),
    .B(_6740_),
    .S(\datapath.idinstr_16_bF$buf13 ),
    .Y(_6742_)
);

NAND2X1 _17683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf41 ),
    .B(_6742_),
    .Y(_6743_)
);

AOI21X1 _17684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6739_),
    .B(_6743_),
    .C(\datapath.idinstr_18_bF$buf2 ),
    .Y(_6744_)
);

OAI21X1 _17685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6744_),
    .B(_6735_),
    .C(_6140__bF$buf1),
    .Y(_6745_)
);

AOI21X1 _17686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6720_),
    .B(_6745_),
    .C(_6147__bF$buf2),
    .Y(\datapath.registers.rega_data [12])
);

MUX2X1 _17687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [13]),
    .B(\datapath.registers.1226[24] [13]),
    .S(\datapath.idinstr_15_bF$buf3 ),
    .Y(_6746_)
);

MUX2X1 _17688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [13]),
    .B(\datapath.registers.1226[26] [13]),
    .S(\datapath.idinstr_15_bF$buf2 ),
    .Y(_6747_)
);

MUX2X1 _17689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6747_),
    .B(_6746_),
    .S(\datapath.idinstr_16_bF$buf12 ),
    .Y(_6748_)
);

NAND2X1 _17690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf0),
    .B(_6748_),
    .Y(_6749_)
);

MUX2X1 _17691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [13]),
    .B(\datapath.registers.1226[28] [13]),
    .S(\datapath.idinstr_15_bF$buf1 ),
    .Y(_6750_)
);

MUX2X1 _17692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [13]),
    .B(\datapath.registers.1226[30] [13]),
    .S(\datapath.idinstr_15_bF$buf0 ),
    .Y(_6751_)
);

MUX2X1 _17693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6751_),
    .B(_6750_),
    .S(\datapath.idinstr_16_bF$buf11 ),
    .Y(_6752_)
);

NAND2X1 _17694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf40 ),
    .B(_6752_),
    .Y(_6753_)
);

AOI21X1 _17695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6749_),
    .B(_6753_),
    .C(_6145__bF$buf4),
    .Y(_6754_)
);

MUX2X1 _17696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [13]),
    .B(\datapath.registers.1226[16] [13]),
    .S(\datapath.idinstr_16_bF$buf10 ),
    .Y(_6755_)
);

NAND2X1 _17697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf6),
    .B(_6755_),
    .Y(_6756_)
);

MUX2X1 _17698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [13]),
    .B(\datapath.registers.1226[17] [13]),
    .S(\datapath.idinstr_16_bF$buf9 ),
    .Y(_6757_)
);

AOI21X1 _17699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf53 ),
    .B(_6757_),
    .C(\datapath.idinstr_17_bF$buf39 ),
    .Y(_6758_)
);

NAND2X1 _17700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6756_),
    .B(_6758_),
    .Y(_6759_)
);

MUX2X1 _17701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [13]),
    .B(\datapath.registers.1226[20] [13]),
    .S(\datapath.idinstr_16_bF$buf8 ),
    .Y(_6760_)
);

NAND2X1 _17702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf5),
    .B(_6760_),
    .Y(_6761_)
);

MUX2X1 _17703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [13]),
    .B(\datapath.registers.1226[21] [13]),
    .S(\datapath.idinstr_16_bF$buf7 ),
    .Y(_6762_)
);

AOI21X1 _17704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf52 ),
    .B(_6762_),
    .C(_6144__bF$buf10),
    .Y(_6763_)
);

NAND2X1 _17705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6761_),
    .B(_6763_),
    .Y(_6764_)
);

AOI21X1 _17706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6759_),
    .B(_6764_),
    .C(\datapath.idinstr_18_bF$buf1 ),
    .Y(_6765_)
);

OAI21X1 _17707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6754_),
    .B(_6765_),
    .C(\datapath.idinstr_19_bF$buf0 ),
    .Y(_6766_)
);

INVX1 _17708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [13]),
    .Y(_6767_)
);

AOI21X1 _17709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [13]),
    .B(\datapath.idinstr_17_bF$buf38 ),
    .C(_6141__bF$buf4),
    .Y(_6768_)
);

OAI21X1 _17710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf37 ),
    .B(_6767_),
    .C(_6768_),
    .Y(_6769_)
);

INVX1 _17711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [13]),
    .Y(_6770_)
);

AOI21X1 _17712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf36 ),
    .B(\datapath.registers.1226[12] [13]),
    .C(\datapath.idinstr_15_bF$buf51 ),
    .Y(_6771_)
);

OAI21X1 _17713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf35 ),
    .B(_6770_),
    .C(_6771_),
    .Y(_6772_)
);

NAND3X1 _17714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf4),
    .B(_6772_),
    .C(_6769_),
    .Y(_6773_)
);

INVX1 _17715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [13]),
    .Y(_6774_)
);

AOI21X1 _17716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [13]),
    .B(\datapath.idinstr_17_bF$buf34 ),
    .C(_6141__bF$buf3),
    .Y(_6775_)
);

OAI21X1 _17717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf33 ),
    .B(_6774_),
    .C(_6775_),
    .Y(_6776_)
);

INVX1 _17718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[10] [13]),
    .Y(_6777_)
);

AOI21X1 _17719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [13]),
    .B(\datapath.idinstr_17_bF$buf32 ),
    .C(\datapath.idinstr_15_bF$buf50 ),
    .Y(_6778_)
);

OAI21X1 _17720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf31 ),
    .B(_6777_),
    .C(_6778_),
    .Y(_6779_)
);

NAND3X1 _17721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_bF$buf6 ),
    .B(_6779_),
    .C(_6776_),
    .Y(_6780_)
);

AOI21X1 _17722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6773_),
    .B(_6780_),
    .C(_6145__bF$buf3),
    .Y(_6781_)
);

MUX2X1 _17723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [13]),
    .B(\datapath.registers.1226[0] [13]),
    .S(\datapath.idinstr_15_bF$buf49 ),
    .Y(_6782_)
);

MUX2X1 _17724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [13]),
    .B(\datapath.registers.1226[2] [13]),
    .S(\datapath.idinstr_15_bF$buf48 ),
    .Y(_6783_)
);

MUX2X1 _17725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6783_),
    .B(_6782_),
    .S(\datapath.idinstr_16_bF$buf5 ),
    .Y(_6784_)
);

NAND2X1 _17726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf9),
    .B(_6784_),
    .Y(_6785_)
);

MUX2X1 _17727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [13]),
    .B(\datapath.registers.1226[4] [13]),
    .S(\datapath.idinstr_15_bF$buf47 ),
    .Y(_6786_)
);

MUX2X1 _17728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [13]),
    .B(\datapath.registers.1226[6] [13]),
    .S(\datapath.idinstr_15_bF$buf46 ),
    .Y(_6787_)
);

MUX2X1 _17729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6787_),
    .B(_6786_),
    .S(\datapath.idinstr_16_bF$buf4 ),
    .Y(_6788_)
);

NAND2X1 _17730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf30 ),
    .B(_6788_),
    .Y(_6789_)
);

AOI21X1 _17731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6785_),
    .B(_6789_),
    .C(\datapath.idinstr_18_bF$buf0 ),
    .Y(_6790_)
);

OAI21X1 _17732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6790_),
    .B(_6781_),
    .C(_6140__bF$buf0),
    .Y(_6791_)
);

AOI21X1 _17733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6766_),
    .B(_6791_),
    .C(_6147__bF$buf1),
    .Y(\datapath.registers.rega_data [13])
);

MUX2X1 _17734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [14]),
    .B(\datapath.registers.1226[24] [14]),
    .S(\datapath.idinstr_15_bF$buf45 ),
    .Y(_6792_)
);

MUX2X1 _17735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [14]),
    .B(\datapath.registers.1226[26] [14]),
    .S(\datapath.idinstr_15_bF$buf44 ),
    .Y(_6793_)
);

MUX2X1 _17736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6793_),
    .B(_6792_),
    .S(\datapath.idinstr_16_bF$buf3 ),
    .Y(_6794_)
);

NAND2X1 _17737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf8),
    .B(_6794_),
    .Y(_6795_)
);

MUX2X1 _17738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [14]),
    .B(\datapath.registers.1226[28] [14]),
    .S(\datapath.idinstr_15_bF$buf43 ),
    .Y(_6796_)
);

MUX2X1 _17739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [14]),
    .B(\datapath.registers.1226[30] [14]),
    .S(\datapath.idinstr_15_bF$buf42 ),
    .Y(_6797_)
);

MUX2X1 _17740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6797_),
    .B(_6796_),
    .S(\datapath.idinstr_16_bF$buf2 ),
    .Y(_6798_)
);

NAND2X1 _17741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf29 ),
    .B(_6798_),
    .Y(_6799_)
);

AOI21X1 _17742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6795_),
    .B(_6799_),
    .C(_6145__bF$buf2),
    .Y(_6800_)
);

MUX2X1 _17743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [14]),
    .B(\datapath.registers.1226[16] [14]),
    .S(\datapath.idinstr_16_bF$buf1 ),
    .Y(_6801_)
);

NAND2X1 _17744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf2),
    .B(_6801_),
    .Y(_6802_)
);

MUX2X1 _17745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [14]),
    .B(\datapath.registers.1226[17] [14]),
    .S(\datapath.idinstr_16_bF$buf0 ),
    .Y(_6803_)
);

AOI21X1 _17746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf41 ),
    .B(_6803_),
    .C(\datapath.idinstr_17_bF$buf28 ),
    .Y(_6804_)
);

NAND2X1 _17747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6802_),
    .B(_6804_),
    .Y(_6805_)
);

MUX2X1 _17748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [14]),
    .B(\datapath.registers.1226[20] [14]),
    .S(\datapath.idinstr_16_bF$buf45 ),
    .Y(_6806_)
);

NAND2X1 _17749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf1),
    .B(_6806_),
    .Y(_6807_)
);

MUX2X1 _17750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [14]),
    .B(\datapath.registers.1226[21] [14]),
    .S(\datapath.idinstr_16_bF$buf44 ),
    .Y(_6808_)
);

AOI21X1 _17751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf40 ),
    .B(_6808_),
    .C(_6144__bF$buf7),
    .Y(_6809_)
);

NAND2X1 _17752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6807_),
    .B(_6809_),
    .Y(_6810_)
);

AOI21X1 _17753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6805_),
    .B(_6810_),
    .C(\datapath.idinstr_18_bF$buf7 ),
    .Y(_6811_)
);

OAI21X1 _17754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6800_),
    .B(_6811_),
    .C(\datapath.idinstr_19_bF$buf5 ),
    .Y(_6812_)
);

MUX2X1 _17755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [14]),
    .B(\datapath.registers.1226[8] [14]),
    .S(\datapath.idinstr_15_bF$buf39 ),
    .Y(_6813_)
);

MUX2X1 _17756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [14]),
    .B(\datapath.registers.1226[10] [14]),
    .S(\datapath.idinstr_15_bF$buf38 ),
    .Y(_6814_)
);

MUX2X1 _17757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6814_),
    .B(_6813_),
    .S(\datapath.idinstr_16_bF$buf43 ),
    .Y(_6815_)
);

NAND2X1 _17758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf6),
    .B(_6815_),
    .Y(_6816_)
);

AND2X2 _17759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [14]),
    .B(\datapath.idinstr_15_bF$buf37 ),
    .Y(_6817_)
);

INVX1 _17760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [14]),
    .Y(_6818_)
);

OAI21X1 _17761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6818_),
    .B(\datapath.idinstr_15_bF$buf36 ),
    .C(\datapath.idinstr_16_bF$buf42 ),
    .Y(_6819_)
);

NAND2X1 _17762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [14]),
    .B(_6141__bF$buf0),
    .Y(_6820_)
);

AOI21X1 _17763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [14]),
    .B(\datapath.idinstr_15_bF$buf35 ),
    .C(\datapath.idinstr_16_bF$buf41 ),
    .Y(_6821_)
);

AOI21X1 _17764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6821_),
    .B(_6820_),
    .C(_6144__bF$buf5),
    .Y(_6822_)
);

OAI21X1 _17765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6817_),
    .B(_6819_),
    .C(_6822_),
    .Y(_6823_)
);

AOI21X1 _17766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6823_),
    .B(_6816_),
    .C(_6145__bF$buf1),
    .Y(_6824_)
);

MUX2X1 _17767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [14]),
    .B(\datapath.registers.1226[4] [14]),
    .S(\datapath.idinstr_15_bF$buf34 ),
    .Y(_6825_)
);

MUX2X1 _17768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [14]),
    .B(\datapath.registers.1226[6] [14]),
    .S(\datapath.idinstr_15_bF$buf33 ),
    .Y(_6826_)
);

MUX2X1 _17769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6826_),
    .B(_6825_),
    .S(\datapath.idinstr_16_bF$buf40 ),
    .Y(_6827_)
);

NAND2X1 _17770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf27 ),
    .B(_6827_),
    .Y(_6828_)
);

MUX2X1 _17771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [14]),
    .B(\datapath.registers.1226[0] [14]),
    .S(\datapath.idinstr_15_bF$buf32 ),
    .Y(_6829_)
);

MUX2X1 _17772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [14]),
    .B(\datapath.registers.1226[2] [14]),
    .S(\datapath.idinstr_15_bF$buf31 ),
    .Y(_6830_)
);

MUX2X1 _17773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6830_),
    .B(_6829_),
    .S(\datapath.idinstr_16_bF$buf39 ),
    .Y(_6831_)
);

NAND2X1 _17774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf4),
    .B(_6831_),
    .Y(_6832_)
);

AOI21X1 _17775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6828_),
    .B(_6832_),
    .C(\datapath.idinstr_18_bF$buf6 ),
    .Y(_6833_)
);

OAI21X1 _17776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6833_),
    .B(_6824_),
    .C(_6140__bF$buf4),
    .Y(_6834_)
);

AOI21X1 _17777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6812_),
    .B(_6834_),
    .C(_6147__bF$buf0),
    .Y(\datapath.registers.rega_data [14])
);

MUX2X1 _17778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [15]),
    .B(\datapath.registers.1226[24] [15]),
    .S(\datapath.idinstr_15_bF$buf30 ),
    .Y(_6835_)
);

MUX2X1 _17779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [15]),
    .B(\datapath.registers.1226[26] [15]),
    .S(\datapath.idinstr_15_bF$buf29 ),
    .Y(_6836_)
);

MUX2X1 _17780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6836_),
    .B(_6835_),
    .S(\datapath.idinstr_16_bF$buf38 ),
    .Y(_6837_)
);

NAND2X1 _17781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf3),
    .B(_6837_),
    .Y(_6838_)
);

MUX2X1 _17782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [15]),
    .B(\datapath.registers.1226[28] [15]),
    .S(\datapath.idinstr_15_bF$buf28 ),
    .Y(_6839_)
);

MUX2X1 _17783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [15]),
    .B(\datapath.registers.1226[30] [15]),
    .S(\datapath.idinstr_15_bF$buf27 ),
    .Y(_6840_)
);

MUX2X1 _17784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6840_),
    .B(_6839_),
    .S(\datapath.idinstr_16_bF$buf37 ),
    .Y(_6841_)
);

NAND2X1 _17785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf26 ),
    .B(_6841_),
    .Y(_6842_)
);

AOI21X1 _17786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6838_),
    .B(_6842_),
    .C(_6145__bF$buf0),
    .Y(_6843_)
);

MUX2X1 _17787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [15]),
    .B(\datapath.registers.1226[16] [15]),
    .S(\datapath.idinstr_16_bF$buf36 ),
    .Y(_6844_)
);

NAND2X1 _17788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf10),
    .B(_6844_),
    .Y(_6845_)
);

MUX2X1 _17789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [15]),
    .B(\datapath.registers.1226[17] [15]),
    .S(\datapath.idinstr_16_bF$buf35 ),
    .Y(_6846_)
);

AOI21X1 _17790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf26 ),
    .B(_6846_),
    .C(\datapath.idinstr_17_bF$buf25 ),
    .Y(_6847_)
);

NAND2X1 _17791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6845_),
    .B(_6847_),
    .Y(_6848_)
);

MUX2X1 _17792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [15]),
    .B(\datapath.registers.1226[20] [15]),
    .S(\datapath.idinstr_16_bF$buf34 ),
    .Y(_6849_)
);

NAND2X1 _17793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf9),
    .B(_6849_),
    .Y(_6850_)
);

MUX2X1 _17794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [15]),
    .B(\datapath.registers.1226[21] [15]),
    .S(\datapath.idinstr_16_bF$buf33 ),
    .Y(_6851_)
);

AOI21X1 _17795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf25 ),
    .B(_6851_),
    .C(_6144__bF$buf2),
    .Y(_6852_)
);

NAND2X1 _17796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6850_),
    .B(_6852_),
    .Y(_6853_)
);

AOI21X1 _17797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6848_),
    .B(_6853_),
    .C(\datapath.idinstr_18_bF$buf5 ),
    .Y(_6854_)
);

OAI21X1 _17798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6843_),
    .B(_6854_),
    .C(\datapath.idinstr_19_bF$buf4 ),
    .Y(_6855_)
);

MUX2X1 _17799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [15]),
    .B(\datapath.registers.1226[8] [15]),
    .S(\datapath.idinstr_15_bF$buf24 ),
    .Y(_6856_)
);

MUX2X1 _17800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [15]),
    .B(\datapath.registers.1226[10] [15]),
    .S(\datapath.idinstr_15_bF$buf23 ),
    .Y(_6857_)
);

MUX2X1 _17801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6857_),
    .B(_6856_),
    .S(\datapath.idinstr_16_bF$buf32 ),
    .Y(_6858_)
);

NAND2X1 _17802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf1),
    .B(_6858_),
    .Y(_6859_)
);

INVX1 _17803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [15]),
    .Y(_6860_)
);

NOR2X1 _17804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6860_),
    .B(_6141__bF$buf8),
    .Y(_6861_)
);

INVX1 _17805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [15]),
    .Y(_6862_)
);

OAI21X1 _17806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6862_),
    .B(\datapath.idinstr_15_bF$buf22 ),
    .C(\datapath.idinstr_16_bF$buf31 ),
    .Y(_6863_)
);

NAND2X1 _17807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [15]),
    .B(_6141__bF$buf7),
    .Y(_6864_)
);

AOI21X1 _17808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [15]),
    .B(\datapath.idinstr_15_bF$buf21 ),
    .C(\datapath.idinstr_16_bF$buf30 ),
    .Y(_6865_)
);

AOI21X1 _17809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6865_),
    .B(_6864_),
    .C(_6144__bF$buf0),
    .Y(_6866_)
);

OAI21X1 _17810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6861_),
    .B(_6863_),
    .C(_6866_),
    .Y(_6867_)
);

AOI21X1 _17811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6867_),
    .B(_6859_),
    .C(_6145__bF$buf7),
    .Y(_6868_)
);

MUX2X1 _17812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [15]),
    .B(\datapath.registers.1226[4] [15]),
    .S(\datapath.idinstr_15_bF$buf20 ),
    .Y(_6869_)
);

MUX2X1 _17813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [15]),
    .B(\datapath.registers.1226[6] [15]),
    .S(\datapath.idinstr_15_bF$buf19 ),
    .Y(_6870_)
);

MUX2X1 _17814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6870_),
    .B(_6869_),
    .S(\datapath.idinstr_16_bF$buf29 ),
    .Y(_6871_)
);

NAND2X1 _17815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf24 ),
    .B(_6871_),
    .Y(_6872_)
);

MUX2X1 _17816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [15]),
    .B(\datapath.registers.1226[0] [15]),
    .S(\datapath.idinstr_15_bF$buf18 ),
    .Y(_6873_)
);

MUX2X1 _17817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [15]),
    .B(\datapath.registers.1226[2] [15]),
    .S(\datapath.idinstr_15_bF$buf17 ),
    .Y(_6874_)
);

MUX2X1 _17818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6874_),
    .B(_6873_),
    .S(\datapath.idinstr_16_bF$buf28 ),
    .Y(_6875_)
);

NAND2X1 _17819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf10),
    .B(_6875_),
    .Y(_6876_)
);

AOI21X1 _17820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6872_),
    .B(_6876_),
    .C(\datapath.idinstr_18_bF$buf4 ),
    .Y(_6877_)
);

OAI21X1 _17821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6877_),
    .B(_6868_),
    .C(_6140__bF$buf3),
    .Y(_6878_)
);

AOI21X1 _17822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6855_),
    .B(_6878_),
    .C(_6147__bF$buf4),
    .Y(\datapath.registers.rega_data [15])
);

MUX2X1 _17823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [16]),
    .B(\datapath.registers.1226[8] [16]),
    .S(\datapath.idinstr_15_bF$buf16 ),
    .Y(_6879_)
);

MUX2X1 _17824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [16]),
    .B(\datapath.registers.1226[10] [16]),
    .S(\datapath.idinstr_15_bF$buf15 ),
    .Y(_6880_)
);

MUX2X1 _17825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6880_),
    .B(_6879_),
    .S(\datapath.idinstr_16_bF$buf27 ),
    .Y(_6881_)
);

NAND2X1 _17826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf9),
    .B(_6881_),
    .Y(_6882_)
);

INVX1 _17827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [16]),
    .Y(_6883_)
);

NOR2X1 _17828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6883_),
    .B(_6141__bF$buf6),
    .Y(_6884_)
);

INVX1 _17829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [16]),
    .Y(_6885_)
);

OAI21X1 _17830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6885_),
    .B(\datapath.idinstr_15_bF$buf14 ),
    .C(\datapath.idinstr_16_bF$buf26 ),
    .Y(_6886_)
);

NAND2X1 _17831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [16]),
    .B(_6141__bF$buf5),
    .Y(_6887_)
);

AOI21X1 _17832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [16]),
    .B(\datapath.idinstr_15_bF$buf13 ),
    .C(\datapath.idinstr_16_bF$buf25 ),
    .Y(_6888_)
);

AOI21X1 _17833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6888_),
    .B(_6887_),
    .C(_6144__bF$buf8),
    .Y(_6889_)
);

OAI21X1 _17834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6884_),
    .B(_6886_),
    .C(_6889_),
    .Y(_6890_)
);

AOI21X1 _17835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6890_),
    .B(_6882_),
    .C(_6145__bF$buf6),
    .Y(_6891_)
);

MUX2X1 _17836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [16]),
    .B(\datapath.registers.1226[4] [16]),
    .S(\datapath.idinstr_15_bF$buf12 ),
    .Y(_6892_)
);

MUX2X1 _17837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [16]),
    .B(\datapath.registers.1226[6] [16]),
    .S(\datapath.idinstr_15_bF$buf11 ),
    .Y(_6893_)
);

MUX2X1 _17838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6893_),
    .B(_6892_),
    .S(\datapath.idinstr_16_bF$buf24 ),
    .Y(_6894_)
);

NAND2X1 _17839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf23 ),
    .B(_6894_),
    .Y(_6895_)
);

MUX2X1 _17840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [16]),
    .B(\datapath.registers.1226[0] [16]),
    .S(\datapath.idinstr_15_bF$buf10 ),
    .Y(_6896_)
);

MUX2X1 _17841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [16]),
    .B(\datapath.registers.1226[2] [16]),
    .S(\datapath.idinstr_15_bF$buf9 ),
    .Y(_6897_)
);

MUX2X1 _17842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6897_),
    .B(_6896_),
    .S(\datapath.idinstr_16_bF$buf23 ),
    .Y(_6898_)
);

NAND2X1 _17843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf7),
    .B(_6898_),
    .Y(_6899_)
);

AOI21X1 _17844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6895_),
    .B(_6899_),
    .C(\datapath.idinstr_18_bF$buf3 ),
    .Y(_6900_)
);

OAI21X1 _17845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6900_),
    .B(_6891_),
    .C(_6140__bF$buf2),
    .Y(_6901_)
);

INVX1 _17846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [16]),
    .Y(_6902_)
);

AOI21X1 _17847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [16]),
    .B(\datapath.idinstr_17_bF$buf22 ),
    .C(_6141__bF$buf4),
    .Y(_6903_)
);

OAI21X1 _17848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6902_),
    .B(\datapath.idinstr_17_bF$buf21 ),
    .C(_6903_),
    .Y(_6904_)
);

NAND2X1 _17849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [16]),
    .B(_6144__bF$buf6),
    .Y(_6905_)
);

AOI21X1 _17850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [16]),
    .B(\datapath.idinstr_17_bF$buf20 ),
    .C(\datapath.idinstr_15_bF$buf8 ),
    .Y(_6906_)
);

AOI21X1 _17851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6906_),
    .B(_6905_),
    .C(_6143__bF$buf3),
    .Y(_6907_)
);

NAND2X1 _17852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6904_),
    .B(_6907_),
    .Y(_6908_)
);

INVX1 _17853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [16]),
    .Y(_6909_)
);

AOI21X1 _17854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [16]),
    .B(\datapath.idinstr_17_bF$buf19 ),
    .C(_6141__bF$buf3),
    .Y(_6910_)
);

OAI21X1 _17855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6909_),
    .B(\datapath.idinstr_17_bF$buf18 ),
    .C(_6910_),
    .Y(_6911_)
);

AOI21X1 _17856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [16]),
    .B(\datapath.idinstr_17_bF$buf17 ),
    .C(\datapath.idinstr_15_bF$buf7 ),
    .Y(_6912_)
);

OAI21X1 _17857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6018_),
    .B(\datapath.idinstr_17_bF$buf16 ),
    .C(_6912_),
    .Y(_6913_)
);

NAND3X1 _17858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf2),
    .B(_6913_),
    .C(_6911_),
    .Y(_6914_)
);

AOI21X1 _17859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6908_),
    .B(_6914_),
    .C(\datapath.idinstr_18_bF$buf2 ),
    .Y(_6915_)
);

MUX2X1 _17860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [16]),
    .B(\datapath.registers.1226[29] [16]),
    .S(\datapath.idinstr_16_bF$buf22 ),
    .Y(_6916_)
);

MUX2X1 _17861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [16]),
    .B(\datapath.registers.1226[28] [16]),
    .S(\datapath.idinstr_16_bF$buf21 ),
    .Y(_6917_)
);

MUX2X1 _17862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6917_),
    .B(_6916_),
    .S(_6141__bF$buf2),
    .Y(_6918_)
);

NAND2X1 _17863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf15 ),
    .B(_6918_),
    .Y(_6919_)
);

MUX2X1 _17864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [16]),
    .B(\datapath.registers.1226[25] [16]),
    .S(\datapath.idinstr_16_bF$buf20 ),
    .Y(_6920_)
);

MUX2X1 _17865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [16]),
    .B(\datapath.registers.1226[24] [16]),
    .S(\datapath.idinstr_16_bF$buf19 ),
    .Y(_6921_)
);

MUX2X1 _17866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6921_),
    .B(_6920_),
    .S(_6141__bF$buf1),
    .Y(_6922_)
);

NAND2X1 _17867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf5),
    .B(_6922_),
    .Y(_6923_)
);

AOI21X1 _17868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6919_),
    .B(_6923_),
    .C(_6145__bF$buf5),
    .Y(_6924_)
);

OAI21X1 _17869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6924_),
    .B(_6915_),
    .C(\datapath.idinstr_19_bF$buf3 ),
    .Y(_6925_)
);

AOI21X1 _17870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6925_),
    .B(_6901_),
    .C(_6147__bF$buf3),
    .Y(\datapath.registers.rega_data [16])
);

MUX2X1 _17871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [17]),
    .B(\datapath.registers.1226[24] [17]),
    .S(\datapath.idinstr_15_bF$buf6 ),
    .Y(_6926_)
);

MUX2X1 _17872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [17]),
    .B(\datapath.registers.1226[26] [17]),
    .S(\datapath.idinstr_15_bF$buf5 ),
    .Y(_6927_)
);

MUX2X1 _17873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6927_),
    .B(_6926_),
    .S(\datapath.idinstr_16_bF$buf18 ),
    .Y(_6928_)
);

NAND2X1 _17874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf4),
    .B(_6928_),
    .Y(_6929_)
);

MUX2X1 _17875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [17]),
    .B(\datapath.registers.1226[28] [17]),
    .S(\datapath.idinstr_15_bF$buf4 ),
    .Y(_6930_)
);

MUX2X1 _17876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [17]),
    .B(\datapath.registers.1226[30] [17]),
    .S(\datapath.idinstr_15_bF$buf3 ),
    .Y(_6931_)
);

MUX2X1 _17877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6931_),
    .B(_6930_),
    .S(\datapath.idinstr_16_bF$buf17 ),
    .Y(_6932_)
);

NAND2X1 _17878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf14 ),
    .B(_6932_),
    .Y(_6933_)
);

AOI21X1 _17879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6929_),
    .B(_6933_),
    .C(_6145__bF$buf4),
    .Y(_6934_)
);

MUX2X1 _17880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [17]),
    .B(\datapath.registers.1226[16] [17]),
    .S(\datapath.idinstr_16_bF$buf16 ),
    .Y(_6935_)
);

NAND2X1 _17881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf0),
    .B(_6935_),
    .Y(_6936_)
);

MUX2X1 _17882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [17]),
    .B(\datapath.registers.1226[17] [17]),
    .S(\datapath.idinstr_16_bF$buf15 ),
    .Y(_6937_)
);

AOI21X1 _17883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf2 ),
    .B(_6937_),
    .C(\datapath.idinstr_17_bF$buf13 ),
    .Y(_6938_)
);

NAND2X1 _17884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6936_),
    .B(_6938_),
    .Y(_6939_)
);

MUX2X1 _17885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [17]),
    .B(\datapath.registers.1226[20] [17]),
    .S(\datapath.idinstr_16_bF$buf14 ),
    .Y(_6940_)
);

NAND2X1 _17886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf10),
    .B(_6940_),
    .Y(_6941_)
);

MUX2X1 _17887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [17]),
    .B(\datapath.registers.1226[21] [17]),
    .S(\datapath.idinstr_16_bF$buf13 ),
    .Y(_6942_)
);

AOI21X1 _17888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf1 ),
    .B(_6942_),
    .C(_6144__bF$buf3),
    .Y(_6943_)
);

NAND2X1 _17889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6941_),
    .B(_6943_),
    .Y(_6944_)
);

AOI21X1 _17890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6939_),
    .B(_6944_),
    .C(\datapath.idinstr_18_bF$buf1 ),
    .Y(_6945_)
);

OAI21X1 _17891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6934_),
    .B(_6945_),
    .C(\datapath.idinstr_19_bF$buf2 ),
    .Y(_6946_)
);

INVX1 _17892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [17]),
    .Y(_6947_)
);

AOI21X1 _17893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [17]),
    .B(\datapath.idinstr_17_bF$buf12 ),
    .C(_6141__bF$buf9),
    .Y(_6948_)
);

OAI21X1 _17894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf11 ),
    .B(_6947_),
    .C(_6948_),
    .Y(_6949_)
);

INVX1 _17895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [17]),
    .Y(_6950_)
);

AOI21X1 _17896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf10 ),
    .B(\datapath.registers.1226[12] [17]),
    .C(\datapath.idinstr_15_bF$buf0 ),
    .Y(_6951_)
);

OAI21X1 _17897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf9 ),
    .B(_6950_),
    .C(_6951_),
    .Y(_6952_)
);

NAND3X1 _17898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf1),
    .B(_6952_),
    .C(_6949_),
    .Y(_6953_)
);

INVX1 _17899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [17]),
    .Y(_6954_)
);

AOI21X1 _17900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [17]),
    .B(\datapath.idinstr_17_bF$buf8 ),
    .C(_6141__bF$buf8),
    .Y(_6955_)
);

OAI21X1 _17901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf7 ),
    .B(_6954_),
    .C(_6955_),
    .Y(_6956_)
);

INVX1 _17902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[10] [17]),
    .Y(_6957_)
);

AOI21X1 _17903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [17]),
    .B(\datapath.idinstr_17_bF$buf6 ),
    .C(\datapath.idinstr_15_bF$buf53 ),
    .Y(_6958_)
);

OAI21X1 _17904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf5 ),
    .B(_6957_),
    .C(_6958_),
    .Y(_6959_)
);

NAND3X1 _17905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_bF$buf12 ),
    .B(_6959_),
    .C(_6956_),
    .Y(_6960_)
);

AOI21X1 _17906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6953_),
    .B(_6960_),
    .C(_6145__bF$buf3),
    .Y(_6961_)
);

MUX2X1 _17907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [17]),
    .B(\datapath.registers.1226[0] [17]),
    .S(\datapath.idinstr_15_bF$buf52 ),
    .Y(_6962_)
);

MUX2X1 _17908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [17]),
    .B(\datapath.registers.1226[2] [17]),
    .S(\datapath.idinstr_15_bF$buf51 ),
    .Y(_6963_)
);

MUX2X1 _17909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6963_),
    .B(_6962_),
    .S(\datapath.idinstr_16_bF$buf11 ),
    .Y(_6964_)
);

NAND2X1 _17910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf2),
    .B(_6964_),
    .Y(_6965_)
);

MUX2X1 _17911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [17]),
    .B(\datapath.registers.1226[4] [17]),
    .S(\datapath.idinstr_15_bF$buf50 ),
    .Y(_6966_)
);

MUX2X1 _17912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [17]),
    .B(\datapath.registers.1226[6] [17]),
    .S(\datapath.idinstr_15_bF$buf49 ),
    .Y(_6967_)
);

MUX2X1 _17913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6967_),
    .B(_6966_),
    .S(\datapath.idinstr_16_bF$buf10 ),
    .Y(_6968_)
);

NAND2X1 _17914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf4 ),
    .B(_6968_),
    .Y(_6969_)
);

AOI21X1 _17915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6965_),
    .B(_6969_),
    .C(\datapath.idinstr_18_bF$buf0 ),
    .Y(_6970_)
);

OAI21X1 _17916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6970_),
    .B(_6961_),
    .C(_6140__bF$buf1),
    .Y(_6971_)
);

AOI21X1 _17917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6946_),
    .B(_6971_),
    .C(_6147__bF$buf2),
    .Y(\datapath.registers.rega_data [17])
);

MUX2X1 _17918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [18]),
    .B(\datapath.registers.1226[24] [18]),
    .S(\datapath.idinstr_15_bF$buf48 ),
    .Y(_6972_)
);

MUX2X1 _17919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [18]),
    .B(\datapath.registers.1226[26] [18]),
    .S(\datapath.idinstr_15_bF$buf47 ),
    .Y(_6973_)
);

MUX2X1 _17920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6973_),
    .B(_6972_),
    .S(\datapath.idinstr_16_bF$buf9 ),
    .Y(_6974_)
);

NAND2X1 _17921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf1),
    .B(_6974_),
    .Y(_6975_)
);

MUX2X1 _17922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [18]),
    .B(\datapath.registers.1226[28] [18]),
    .S(\datapath.idinstr_15_bF$buf46 ),
    .Y(_6976_)
);

MUX2X1 _17923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [18]),
    .B(\datapath.registers.1226[30] [18]),
    .S(\datapath.idinstr_15_bF$buf45 ),
    .Y(_6977_)
);

MUX2X1 _17924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6977_),
    .B(_6976_),
    .S(\datapath.idinstr_16_bF$buf8 ),
    .Y(_6978_)
);

NAND2X1 _17925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf3 ),
    .B(_6978_),
    .Y(_6979_)
);

AOI21X1 _17926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6975_),
    .B(_6979_),
    .C(_6145__bF$buf2),
    .Y(_6980_)
);

MUX2X1 _17927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [18]),
    .B(\datapath.registers.1226[16] [18]),
    .S(\datapath.idinstr_16_bF$buf7 ),
    .Y(_6981_)
);

NAND2X1 _17928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf7),
    .B(_6981_),
    .Y(_6982_)
);

MUX2X1 _17929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [18]),
    .B(\datapath.registers.1226[17] [18]),
    .S(\datapath.idinstr_16_bF$buf6 ),
    .Y(_6983_)
);

AOI21X1 _17930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf44 ),
    .B(_6983_),
    .C(\datapath.idinstr_17_bF$buf2 ),
    .Y(_6984_)
);

NAND2X1 _17931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6982_),
    .B(_6984_),
    .Y(_6985_)
);

MUX2X1 _17932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [18]),
    .B(\datapath.registers.1226[20] [18]),
    .S(\datapath.idinstr_16_bF$buf5 ),
    .Y(_6986_)
);

NAND2X1 _17933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf6),
    .B(_6986_),
    .Y(_6987_)
);

MUX2X1 _17934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [18]),
    .B(\datapath.registers.1226[21] [18]),
    .S(\datapath.idinstr_16_bF$buf4 ),
    .Y(_6988_)
);

AOI21X1 _17935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf43 ),
    .B(_6988_),
    .C(_6144__bF$buf0),
    .Y(_6989_)
);

NAND2X1 _17936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6987_),
    .B(_6989_),
    .Y(_6990_)
);

AOI21X1 _17937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6985_),
    .B(_6990_),
    .C(\datapath.idinstr_18_bF$buf7 ),
    .Y(_6991_)
);

OAI21X1 _17938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6980_),
    .B(_6991_),
    .C(\datapath.idinstr_19_bF$buf1 ),
    .Y(_6992_)
);

MUX2X1 _17939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [18]),
    .B(\datapath.registers.1226[8] [18]),
    .S(\datapath.idinstr_15_bF$buf42 ),
    .Y(_6993_)
);

MUX2X1 _17940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [18]),
    .B(\datapath.registers.1226[10] [18]),
    .S(\datapath.idinstr_15_bF$buf41 ),
    .Y(_6994_)
);

MUX2X1 _17941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6994_),
    .B(_6993_),
    .S(\datapath.idinstr_16_bF$buf3 ),
    .Y(_6995_)
);

NAND2X1 _17942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf10),
    .B(_6995_),
    .Y(_6996_)
);

AND2X2 _17943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [18]),
    .B(\datapath.idinstr_15_bF$buf40 ),
    .Y(_6997_)
);

INVX1 _17944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [18]),
    .Y(_6998_)
);

OAI21X1 _17945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6998_),
    .B(\datapath.idinstr_15_bF$buf39 ),
    .C(\datapath.idinstr_16_bF$buf2 ),
    .Y(_6999_)
);

NAND2X1 _17946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [18]),
    .B(_6141__bF$buf5),
    .Y(_7000_)
);

AOI21X1 _17947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [18]),
    .B(\datapath.idinstr_15_bF$buf38 ),
    .C(\datapath.idinstr_16_bF$buf1 ),
    .Y(_7001_)
);

AOI21X1 _17948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7001_),
    .B(_7000_),
    .C(_6144__bF$buf9),
    .Y(_7002_)
);

OAI21X1 _17949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6997_),
    .B(_6999_),
    .C(_7002_),
    .Y(_7003_)
);

AOI21X1 _17950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7003_),
    .B(_6996_),
    .C(_6145__bF$buf1),
    .Y(_7004_)
);

MUX2X1 _17951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [18]),
    .B(\datapath.registers.1226[4] [18]),
    .S(\datapath.idinstr_15_bF$buf37 ),
    .Y(_7005_)
);

MUX2X1 _17952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [18]),
    .B(\datapath.registers.1226[6] [18]),
    .S(\datapath.idinstr_15_bF$buf36 ),
    .Y(_7006_)
);

MUX2X1 _17953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7006_),
    .B(_7005_),
    .S(\datapath.idinstr_16_bF$buf0 ),
    .Y(_7007_)
);

NAND2X1 _17954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf1 ),
    .B(_7007_),
    .Y(_7008_)
);

MUX2X1 _17955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [18]),
    .B(\datapath.registers.1226[0] [18]),
    .S(\datapath.idinstr_15_bF$buf35 ),
    .Y(_7009_)
);

MUX2X1 _17956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [18]),
    .B(\datapath.registers.1226[2] [18]),
    .S(\datapath.idinstr_15_bF$buf34 ),
    .Y(_7010_)
);

MUX2X1 _17957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7010_),
    .B(_7009_),
    .S(\datapath.idinstr_16_bF$buf45 ),
    .Y(_7011_)
);

NAND2X1 _17958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf8),
    .B(_7011_),
    .Y(_7012_)
);

AOI21X1 _17959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7008_),
    .B(_7012_),
    .C(\datapath.idinstr_18_bF$buf6 ),
    .Y(_7013_)
);

OAI21X1 _17960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7013_),
    .B(_7004_),
    .C(_6140__bF$buf0),
    .Y(_7014_)
);

AOI21X1 _17961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6992_),
    .B(_7014_),
    .C(_6147__bF$buf1),
    .Y(\datapath.registers.rega_data [18])
);

MUX2X1 _17962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [19]),
    .B(\datapath.registers.1226[24] [19]),
    .S(\datapath.idinstr_15_bF$buf33 ),
    .Y(_7015_)
);

MUX2X1 _17963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [19]),
    .B(\datapath.registers.1226[26] [19]),
    .S(\datapath.idinstr_15_bF$buf32 ),
    .Y(_7016_)
);

MUX2X1 _17964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7016_),
    .B(_7015_),
    .S(\datapath.idinstr_16_bF$buf44 ),
    .Y(_7017_)
);

NAND2X1 _17965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf7),
    .B(_7017_),
    .Y(_7018_)
);

MUX2X1 _17966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [19]),
    .B(\datapath.registers.1226[28] [19]),
    .S(\datapath.idinstr_15_bF$buf31 ),
    .Y(_7019_)
);

MUX2X1 _17967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [19]),
    .B(\datapath.registers.1226[30] [19]),
    .S(\datapath.idinstr_15_bF$buf30 ),
    .Y(_7020_)
);

MUX2X1 _17968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7020_),
    .B(_7019_),
    .S(\datapath.idinstr_16_bF$buf43 ),
    .Y(_7021_)
);

NAND2X1 _17969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf0 ),
    .B(_7021_),
    .Y(_7022_)
);

AOI21X1 _17970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7018_),
    .B(_7022_),
    .C(_6145__bF$buf0),
    .Y(_7023_)
);

MUX2X1 _17971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [19]),
    .B(\datapath.registers.1226[16] [19]),
    .S(\datapath.idinstr_16_bF$buf42 ),
    .Y(_7024_)
);

NAND2X1 _17972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf4),
    .B(_7024_),
    .Y(_7025_)
);

MUX2X1 _17973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [19]),
    .B(\datapath.registers.1226[17] [19]),
    .S(\datapath.idinstr_16_bF$buf41 ),
    .Y(_7026_)
);

AOI21X1 _17974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf29 ),
    .B(_7026_),
    .C(\datapath.idinstr_17_bF$buf41 ),
    .Y(_7027_)
);

NAND2X1 _17975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7025_),
    .B(_7027_),
    .Y(_7028_)
);

MUX2X1 _17976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [19]),
    .B(\datapath.registers.1226[20] [19]),
    .S(\datapath.idinstr_16_bF$buf40 ),
    .Y(_7029_)
);

NAND2X1 _17977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf3),
    .B(_7029_),
    .Y(_7030_)
);

MUX2X1 _17978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [19]),
    .B(\datapath.registers.1226[21] [19]),
    .S(\datapath.idinstr_16_bF$buf39 ),
    .Y(_7031_)
);

AOI21X1 _17979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf28 ),
    .B(_7031_),
    .C(_6144__bF$buf6),
    .Y(_7032_)
);

NAND2X1 _17980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7030_),
    .B(_7032_),
    .Y(_7033_)
);

AOI21X1 _17981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7028_),
    .B(_7033_),
    .C(\datapath.idinstr_18_bF$buf5 ),
    .Y(_7034_)
);

OAI21X1 _17982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7023_),
    .B(_7034_),
    .C(\datapath.idinstr_19_bF$buf0 ),
    .Y(_7035_)
);

MUX2X1 _17983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [19]),
    .B(\datapath.registers.1226[8] [19]),
    .S(\datapath.idinstr_15_bF$buf27 ),
    .Y(_7036_)
);

MUX2X1 _17984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [19]),
    .B(\datapath.registers.1226[10] [19]),
    .S(\datapath.idinstr_15_bF$buf26 ),
    .Y(_7037_)
);

MUX2X1 _17985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7037_),
    .B(_7036_),
    .S(\datapath.idinstr_16_bF$buf38 ),
    .Y(_7038_)
);

NAND2X1 _17986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf5),
    .B(_7038_),
    .Y(_7039_)
);

MUX2X1 _17987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [19]),
    .B(\datapath.registers.1226[12] [19]),
    .S(\datapath.idinstr_15_bF$buf25 ),
    .Y(_7040_)
);

MUX2X1 _17988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [19]),
    .B(\datapath.registers.1226[14] [19]),
    .S(\datapath.idinstr_15_bF$buf24 ),
    .Y(_7041_)
);

MUX2X1 _17989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7041_),
    .B(_7040_),
    .S(\datapath.idinstr_16_bF$buf37 ),
    .Y(_7042_)
);

NAND2X1 _17990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf40 ),
    .B(_7042_),
    .Y(_7043_)
);

AOI21X1 _17991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7039_),
    .B(_7043_),
    .C(_6145__bF$buf7),
    .Y(_7044_)
);

INVX1 _17992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [19]),
    .Y(_7045_)
);

AOI21X1 _17993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf39 ),
    .B(\datapath.registers.1226[5] [19]),
    .C(_6141__bF$buf2),
    .Y(_7046_)
);

OAI21X1 _17994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf38 ),
    .B(_7045_),
    .C(_7046_),
    .Y(_7047_)
);

INVX1 _17995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [19]),
    .Y(_7048_)
);

AOI21X1 _17996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf37 ),
    .B(\datapath.registers.1226[4] [19]),
    .C(\datapath.idinstr_15_bF$buf23 ),
    .Y(_7049_)
);

OAI21X1 _17997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7048_),
    .B(\datapath.idinstr_17_bF$buf36 ),
    .C(_7049_),
    .Y(_7050_)
);

NAND3X1 _17998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf0),
    .B(_7050_),
    .C(_7047_),
    .Y(_7051_)
);

INVX2 _17999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [19]),
    .Y(_7052_)
);

AOI21X1 _18000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf35 ),
    .B(\datapath.registers.1226[7] [19]),
    .C(_6141__bF$buf1),
    .Y(_7053_)
);

OAI21X1 _18001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf34 ),
    .B(_7052_),
    .C(_7053_),
    .Y(_7054_)
);

INVX1 _18002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[2] [19]),
    .Y(_7055_)
);

AOI21X1 _18003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf33 ),
    .B(\datapath.registers.1226[6] [19]),
    .C(\datapath.idinstr_15_bF$buf22 ),
    .Y(_7056_)
);

OAI21X1 _18004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf32 ),
    .B(_7055_),
    .C(_7056_),
    .Y(_7057_)
);

NAND3X1 _18005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_bF$buf36 ),
    .B(_7057_),
    .C(_7054_),
    .Y(_7058_)
);

AOI21X1 _18006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7051_),
    .B(_7058_),
    .C(\datapath.idinstr_18_bF$buf4 ),
    .Y(_7059_)
);

OAI21X1 _18007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7044_),
    .B(_7059_),
    .C(_6140__bF$buf4),
    .Y(_7060_)
);

AOI21X1 _18008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7035_),
    .B(_7060_),
    .C(_6147__bF$buf0),
    .Y(\datapath.registers.rega_data [19])
);

MUX2X1 _18009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [20]),
    .B(\datapath.registers.1226[8] [20]),
    .S(\datapath.idinstr_15_bF$buf21 ),
    .Y(_7061_)
);

MUX2X1 _18010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [20]),
    .B(\datapath.registers.1226[10] [20]),
    .S(\datapath.idinstr_15_bF$buf20 ),
    .Y(_7062_)
);

MUX2X1 _18011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7062_),
    .B(_7061_),
    .S(\datapath.idinstr_16_bF$buf35 ),
    .Y(_7063_)
);

NAND2X1 _18012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf4),
    .B(_7063_),
    .Y(_7064_)
);

INVX1 _18013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [20]),
    .Y(_7065_)
);

NOR2X1 _18014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7065_),
    .B(_6141__bF$buf0),
    .Y(_7066_)
);

INVX1 _18015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [20]),
    .Y(_7067_)
);

OAI21X1 _18016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7067_),
    .B(\datapath.idinstr_15_bF$buf19 ),
    .C(\datapath.idinstr_16_bF$buf34 ),
    .Y(_7068_)
);

NAND2X1 _18017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [20]),
    .B(_6141__bF$buf10),
    .Y(_7069_)
);

AOI21X1 _18018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [20]),
    .B(\datapath.idinstr_15_bF$buf18 ),
    .C(\datapath.idinstr_16_bF$buf33 ),
    .Y(_7070_)
);

AOI21X1 _18019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7070_),
    .B(_7069_),
    .C(_6144__bF$buf3),
    .Y(_7071_)
);

OAI21X1 _18020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7066_),
    .B(_7068_),
    .C(_7071_),
    .Y(_7072_)
);

AOI21X1 _18021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7072_),
    .B(_7064_),
    .C(_6145__bF$buf6),
    .Y(_7073_)
);

MUX2X1 _18022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [20]),
    .B(\datapath.registers.1226[4] [20]),
    .S(\datapath.idinstr_15_bF$buf17 ),
    .Y(_7074_)
);

MUX2X1 _18023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [20]),
    .B(\datapath.registers.1226[6] [20]),
    .S(\datapath.idinstr_15_bF$buf16 ),
    .Y(_7075_)
);

MUX2X1 _18024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7075_),
    .B(_7074_),
    .S(\datapath.idinstr_16_bF$buf32 ),
    .Y(_7076_)
);

NAND2X1 _18025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf31 ),
    .B(_7076_),
    .Y(_7077_)
);

MUX2X1 _18026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [20]),
    .B(\datapath.registers.1226[0] [20]),
    .S(\datapath.idinstr_15_bF$buf15 ),
    .Y(_7078_)
);

MUX2X1 _18027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [20]),
    .B(\datapath.registers.1226[2] [20]),
    .S(\datapath.idinstr_15_bF$buf14 ),
    .Y(_7079_)
);

MUX2X1 _18028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7079_),
    .B(_7078_),
    .S(\datapath.idinstr_16_bF$buf31 ),
    .Y(_7080_)
);

NAND2X1 _18029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf2),
    .B(_7080_),
    .Y(_7081_)
);

AOI21X1 _18030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7077_),
    .B(_7081_),
    .C(\datapath.idinstr_18_bF$buf3 ),
    .Y(_7082_)
);

OAI21X1 _18031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7082_),
    .B(_7073_),
    .C(_6140__bF$buf3),
    .Y(_7083_)
);

INVX1 _18032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [20]),
    .Y(_7084_)
);

AOI21X1 _18033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [20]),
    .B(\datapath.idinstr_17_bF$buf30 ),
    .C(_6141__bF$buf9),
    .Y(_7085_)
);

OAI21X1 _18034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7084_),
    .B(\datapath.idinstr_17_bF$buf29 ),
    .C(_7085_),
    .Y(_7086_)
);

NAND2X1 _18035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [20]),
    .B(_6144__bF$buf1),
    .Y(_7087_)
);

AOI21X1 _18036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [20]),
    .B(\datapath.idinstr_17_bF$buf28 ),
    .C(\datapath.idinstr_15_bF$buf13 ),
    .Y(_7088_)
);

AOI21X1 _18037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7088_),
    .B(_7087_),
    .C(_6143__bF$buf4),
    .Y(_7089_)
);

NAND2X1 _18038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7086_),
    .B(_7089_),
    .Y(_7090_)
);

INVX1 _18039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [20]),
    .Y(_7091_)
);

AOI21X1 _18040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [20]),
    .B(\datapath.idinstr_17_bF$buf27 ),
    .C(_6141__bF$buf8),
    .Y(_7092_)
);

OAI21X1 _18041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7091_),
    .B(\datapath.idinstr_17_bF$buf26 ),
    .C(_7092_),
    .Y(_7093_)
);

AOI21X1 _18042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[28] [20]),
    .B(\datapath.idinstr_17_bF$buf25 ),
    .C(\datapath.idinstr_15_bF$buf12 ),
    .Y(_7094_)
);

OAI21X1 _18043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5740_),
    .B(\datapath.idinstr_17_bF$buf24 ),
    .C(_7094_),
    .Y(_7095_)
);

NAND3X1 _18044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf3),
    .B(_7095_),
    .C(_7093_),
    .Y(_7096_)
);

AOI21X1 _18045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7090_),
    .B(_7096_),
    .C(_6145__bF$buf5),
    .Y(_7097_)
);

MUX2X1 _18046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [20]),
    .B(\datapath.registers.1226[16] [20]),
    .S(\datapath.idinstr_15_bF$buf11 ),
    .Y(_7098_)
);

MUX2X1 _18047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [20]),
    .B(\datapath.registers.1226[18] [20]),
    .S(\datapath.idinstr_15_bF$buf10 ),
    .Y(_7099_)
);

MUX2X1 _18048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7099_),
    .B(_7098_),
    .S(\datapath.idinstr_16_bF$buf30 ),
    .Y(_7100_)
);

NAND2X1 _18049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf0),
    .B(_7100_),
    .Y(_7101_)
);

MUX2X1 _18050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [20]),
    .B(\datapath.registers.1226[20] [20]),
    .S(\datapath.idinstr_15_bF$buf9 ),
    .Y(_7102_)
);

MUX2X1 _18051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [20]),
    .B(\datapath.registers.1226[22] [20]),
    .S(\datapath.idinstr_15_bF$buf8 ),
    .Y(_7103_)
);

MUX2X1 _18052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7103_),
    .B(_7102_),
    .S(\datapath.idinstr_16_bF$buf29 ),
    .Y(_7104_)
);

NAND2X1 _18053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf23 ),
    .B(_7104_),
    .Y(_7105_)
);

AOI21X1 _18054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7101_),
    .B(_7105_),
    .C(\datapath.idinstr_18_bF$buf2 ),
    .Y(_7106_)
);

OAI21X1 _18055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7106_),
    .B(_7097_),
    .C(\datapath.idinstr_19_bF$buf5 ),
    .Y(_7107_)
);

AOI21X1 _18056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7107_),
    .B(_7083_),
    .C(_6147__bF$buf4),
    .Y(\datapath.registers.rega_data [20])
);

MUX2X1 _18057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [21]),
    .B(\datapath.registers.1226[8] [21]),
    .S(\datapath.idinstr_15_bF$buf7 ),
    .Y(_7108_)
);

MUX2X1 _18058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [21]),
    .B(\datapath.registers.1226[10] [21]),
    .S(\datapath.idinstr_15_bF$buf6 ),
    .Y(_7109_)
);

MUX2X1 _18059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7109_),
    .B(_7108_),
    .S(\datapath.idinstr_16_bF$buf28 ),
    .Y(_7110_)
);

NAND2X1 _18060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf10),
    .B(_7110_),
    .Y(_7111_)
);

INVX1 _18061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [21]),
    .Y(_7112_)
);

NOR2X1 _18062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7112_),
    .B(_6141__bF$buf7),
    .Y(_7113_)
);

INVX1 _18063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [21]),
    .Y(_7114_)
);

OAI21X1 _18064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7114_),
    .B(\datapath.idinstr_15_bF$buf5 ),
    .C(\datapath.idinstr_16_bF$buf27 ),
    .Y(_7115_)
);

NAND2X1 _18065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [21]),
    .B(_6141__bF$buf6),
    .Y(_7116_)
);

AOI21X1 _18066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [21]),
    .B(\datapath.idinstr_15_bF$buf4 ),
    .C(\datapath.idinstr_16_bF$buf26 ),
    .Y(_7117_)
);

AOI21X1 _18067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7117_),
    .B(_7116_),
    .C(_6144__bF$buf9),
    .Y(_7118_)
);

OAI21X1 _18068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7113_),
    .B(_7115_),
    .C(_7118_),
    .Y(_7119_)
);

AOI21X1 _18069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7119_),
    .B(_7111_),
    .C(_6145__bF$buf4),
    .Y(_7120_)
);

MUX2X1 _18070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [21]),
    .B(\datapath.registers.1226[4] [21]),
    .S(\datapath.idinstr_15_bF$buf3 ),
    .Y(_7121_)
);

MUX2X1 _18071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [21]),
    .B(\datapath.registers.1226[6] [21]),
    .S(\datapath.idinstr_15_bF$buf2 ),
    .Y(_7122_)
);

MUX2X1 _18072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7122_),
    .B(_7121_),
    .S(\datapath.idinstr_16_bF$buf25 ),
    .Y(_7123_)
);

NAND2X1 _18073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf22 ),
    .B(_7123_),
    .Y(_7124_)
);

MUX2X1 _18074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [21]),
    .B(\datapath.registers.1226[0] [21]),
    .S(\datapath.idinstr_15_bF$buf1 ),
    .Y(_7125_)
);

MUX2X1 _18075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [21]),
    .B(\datapath.registers.1226[2] [21]),
    .S(\datapath.idinstr_15_bF$buf0 ),
    .Y(_7126_)
);

MUX2X1 _18076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7126_),
    .B(_7125_),
    .S(\datapath.idinstr_16_bF$buf24 ),
    .Y(_7127_)
);

NAND2X1 _18077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf8),
    .B(_7127_),
    .Y(_7128_)
);

AOI21X1 _18078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7124_),
    .B(_7128_),
    .C(\datapath.idinstr_18_bF$buf1 ),
    .Y(_7129_)
);

OAI21X1 _18079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7129_),
    .B(_7120_),
    .C(_6140__bF$buf2),
    .Y(_7130_)
);

INVX1 _18080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [21]),
    .Y(_7131_)
);

AOI21X1 _18081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [21]),
    .B(\datapath.idinstr_17_bF$buf21 ),
    .C(_6141__bF$buf5),
    .Y(_7132_)
);

OAI21X1 _18082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7131_),
    .B(\datapath.idinstr_17_bF$buf20 ),
    .C(_7132_),
    .Y(_7133_)
);

NAND2X1 _18083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [21]),
    .B(_6144__bF$buf7),
    .Y(_7134_)
);

AOI21X1 _18084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [21]),
    .B(\datapath.idinstr_17_bF$buf19 ),
    .C(\datapath.idinstr_15_bF$buf53 ),
    .Y(_7135_)
);

AOI21X1 _18085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7135_),
    .B(_7134_),
    .C(_6143__bF$buf2),
    .Y(_7136_)
);

NAND2X1 _18086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7133_),
    .B(_7136_),
    .Y(_7137_)
);

INVX1 _18087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [21]),
    .Y(_7138_)
);

AOI21X1 _18088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [21]),
    .B(\datapath.idinstr_17_bF$buf18 ),
    .C(_6141__bF$buf4),
    .Y(_7139_)
);

OAI21X1 _18089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7138_),
    .B(\datapath.idinstr_17_bF$buf17 ),
    .C(_7139_),
    .Y(_7140_)
);

AOI21X1 _18090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [21]),
    .B(\datapath.idinstr_17_bF$buf16 ),
    .C(\datapath.idinstr_15_bF$buf52 ),
    .Y(_7141_)
);

OAI21X1 _18091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6024_),
    .B(\datapath.idinstr_17_bF$buf15 ),
    .C(_7141_),
    .Y(_7142_)
);

NAND3X1 _18092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf1),
    .B(_7142_),
    .C(_7140_),
    .Y(_7143_)
);

AOI21X1 _18093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7137_),
    .B(_7143_),
    .C(\datapath.idinstr_18_bF$buf0 ),
    .Y(_7144_)
);

MUX2X1 _18094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [21]),
    .B(\datapath.registers.1226[29] [21]),
    .S(\datapath.idinstr_16_bF$buf23 ),
    .Y(_7145_)
);

MUX2X1 _18095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [21]),
    .B(\datapath.registers.1226[28] [21]),
    .S(\datapath.idinstr_16_bF$buf22 ),
    .Y(_7146_)
);

MUX2X1 _18096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7146_),
    .B(_7145_),
    .S(_6141__bF$buf3),
    .Y(_7147_)
);

NAND2X1 _18097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf14 ),
    .B(_7147_),
    .Y(_7148_)
);

MUX2X1 _18098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [21]),
    .B(\datapath.registers.1226[25] [21]),
    .S(\datapath.idinstr_16_bF$buf21 ),
    .Y(_7149_)
);

MUX2X1 _18099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [21]),
    .B(\datapath.registers.1226[24] [21]),
    .S(\datapath.idinstr_16_bF$buf20 ),
    .Y(_7150_)
);

MUX2X1 _18100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7150_),
    .B(_7149_),
    .S(_6141__bF$buf2),
    .Y(_7151_)
);

NAND2X1 _18101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf6),
    .B(_7151_),
    .Y(_7152_)
);

AOI21X1 _18102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7148_),
    .B(_7152_),
    .C(_6145__bF$buf3),
    .Y(_7153_)
);

OAI21X1 _18103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7153_),
    .B(_7144_),
    .C(\datapath.idinstr_19_bF$buf4 ),
    .Y(_7154_)
);

AOI21X1 _18104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7154_),
    .B(_7130_),
    .C(_6147__bF$buf3),
    .Y(\datapath.registers.rega_data [21])
);

MUX2X1 _18105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [22]),
    .B(\datapath.registers.1226[24] [22]),
    .S(\datapath.idinstr_15_bF$buf51 ),
    .Y(_7155_)
);

MUX2X1 _18106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [22]),
    .B(\datapath.registers.1226[26] [22]),
    .S(\datapath.idinstr_15_bF$buf50 ),
    .Y(_7156_)
);

MUX2X1 _18107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7156_),
    .B(_7155_),
    .S(\datapath.idinstr_16_bF$buf19 ),
    .Y(_7157_)
);

NAND2X1 _18108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf5),
    .B(_7157_),
    .Y(_7158_)
);

MUX2X1 _18109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [22]),
    .B(\datapath.registers.1226[28] [22]),
    .S(\datapath.idinstr_15_bF$buf49 ),
    .Y(_7159_)
);

MUX2X1 _18110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [22]),
    .B(\datapath.registers.1226[30] [22]),
    .S(\datapath.idinstr_15_bF$buf48 ),
    .Y(_7160_)
);

MUX2X1 _18111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7160_),
    .B(_7159_),
    .S(\datapath.idinstr_16_bF$buf18 ),
    .Y(_7161_)
);

NAND2X1 _18112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf13 ),
    .B(_7161_),
    .Y(_7162_)
);

AOI21X1 _18113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7158_),
    .B(_7162_),
    .C(_6145__bF$buf2),
    .Y(_7163_)
);

MUX2X1 _18114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [22]),
    .B(\datapath.registers.1226[16] [22]),
    .S(\datapath.idinstr_16_bF$buf17 ),
    .Y(_7164_)
);

NAND2X1 _18115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf1),
    .B(_7164_),
    .Y(_7165_)
);

MUX2X1 _18116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [22]),
    .B(\datapath.registers.1226[17] [22]),
    .S(\datapath.idinstr_16_bF$buf16 ),
    .Y(_7166_)
);

AOI21X1 _18117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf47 ),
    .B(_7166_),
    .C(\datapath.idinstr_17_bF$buf12 ),
    .Y(_7167_)
);

NAND2X1 _18118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7165_),
    .B(_7167_),
    .Y(_7168_)
);

MUX2X1 _18119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [22]),
    .B(\datapath.registers.1226[20] [22]),
    .S(\datapath.idinstr_16_bF$buf15 ),
    .Y(_7169_)
);

NAND2X1 _18120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf0),
    .B(_7169_),
    .Y(_7170_)
);

MUX2X1 _18121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [22]),
    .B(\datapath.registers.1226[21] [22]),
    .S(\datapath.idinstr_16_bF$buf14 ),
    .Y(_7171_)
);

AOI21X1 _18122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf46 ),
    .B(_7171_),
    .C(_6144__bF$buf4),
    .Y(_7172_)
);

NAND2X1 _18123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7170_),
    .B(_7172_),
    .Y(_7173_)
);

AOI21X1 _18124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7168_),
    .B(_7173_),
    .C(\datapath.idinstr_18_bF$buf7 ),
    .Y(_7174_)
);

OAI21X1 _18125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7163_),
    .B(_7174_),
    .C(\datapath.idinstr_19_bF$buf3 ),
    .Y(_7175_)
);

MUX2X1 _18126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [22]),
    .B(\datapath.registers.1226[8] [22]),
    .S(\datapath.idinstr_15_bF$buf45 ),
    .Y(_7176_)
);

MUX2X1 _18127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [22]),
    .B(\datapath.registers.1226[10] [22]),
    .S(\datapath.idinstr_15_bF$buf44 ),
    .Y(_7177_)
);

MUX2X1 _18128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7177_),
    .B(_7176_),
    .S(\datapath.idinstr_16_bF$buf13 ),
    .Y(_7178_)
);

NAND2X1 _18129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf3),
    .B(_7178_),
    .Y(_7179_)
);

INVX1 _18130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [22]),
    .Y(_7180_)
);

NOR2X1 _18131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7180_),
    .B(_6141__bF$buf10),
    .Y(_7181_)
);

INVX1 _18132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [22]),
    .Y(_7182_)
);

OAI21X1 _18133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7182_),
    .B(\datapath.idinstr_15_bF$buf43 ),
    .C(\datapath.idinstr_16_bF$buf12 ),
    .Y(_7183_)
);

NAND2X1 _18134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [22]),
    .B(_6141__bF$buf9),
    .Y(_7184_)
);

AOI21X1 _18135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [22]),
    .B(\datapath.idinstr_15_bF$buf42 ),
    .C(\datapath.idinstr_16_bF$buf11 ),
    .Y(_7185_)
);

AOI21X1 _18136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7185_),
    .B(_7184_),
    .C(_6144__bF$buf2),
    .Y(_7186_)
);

OAI21X1 _18137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7181_),
    .B(_7183_),
    .C(_7186_),
    .Y(_7187_)
);

AOI21X1 _18138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7187_),
    .B(_7179_),
    .C(_6145__bF$buf1),
    .Y(_7188_)
);

MUX2X1 _18139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [22]),
    .B(\datapath.registers.1226[4] [22]),
    .S(\datapath.idinstr_15_bF$buf41 ),
    .Y(_7189_)
);

MUX2X1 _18140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [22]),
    .B(\datapath.registers.1226[6] [22]),
    .S(\datapath.idinstr_15_bF$buf40 ),
    .Y(_7190_)
);

MUX2X1 _18141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7190_),
    .B(_7189_),
    .S(\datapath.idinstr_16_bF$buf10 ),
    .Y(_7191_)
);

NAND2X1 _18142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf11 ),
    .B(_7191_),
    .Y(_7192_)
);

MUX2X1 _18143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [22]),
    .B(\datapath.registers.1226[0] [22]),
    .S(\datapath.idinstr_15_bF$buf39 ),
    .Y(_7193_)
);

MUX2X1 _18144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [22]),
    .B(\datapath.registers.1226[2] [22]),
    .S(\datapath.idinstr_15_bF$buf38 ),
    .Y(_7194_)
);

MUX2X1 _18145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7194_),
    .B(_7193_),
    .S(\datapath.idinstr_16_bF$buf9 ),
    .Y(_7195_)
);

NAND2X1 _18146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf1),
    .B(_7195_),
    .Y(_7196_)
);

AOI21X1 _18147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7192_),
    .B(_7196_),
    .C(\datapath.idinstr_18_bF$buf6 ),
    .Y(_7197_)
);

OAI21X1 _18148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7197_),
    .B(_7188_),
    .C(_6140__bF$buf1),
    .Y(_7198_)
);

AOI21X1 _18149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7175_),
    .B(_7198_),
    .C(_6147__bF$buf2),
    .Y(\datapath.registers.rega_data [22])
);

MUX2X1 _18150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [23]),
    .B(\datapath.registers.1226[24] [23]),
    .S(\datapath.idinstr_15_bF$buf37 ),
    .Y(_7199_)
);

MUX2X1 _18151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [23]),
    .B(\datapath.registers.1226[26] [23]),
    .S(\datapath.idinstr_15_bF$buf36 ),
    .Y(_7200_)
);

MUX2X1 _18152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7200_),
    .B(_7199_),
    .S(\datapath.idinstr_16_bF$buf8 ),
    .Y(_7201_)
);

NAND2X1 _18153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf0),
    .B(_7201_),
    .Y(_7202_)
);

MUX2X1 _18154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [23]),
    .B(\datapath.registers.1226[28] [23]),
    .S(\datapath.idinstr_15_bF$buf35 ),
    .Y(_7203_)
);

MUX2X1 _18155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [23]),
    .B(\datapath.registers.1226[30] [23]),
    .S(\datapath.idinstr_15_bF$buf34 ),
    .Y(_7204_)
);

MUX2X1 _18156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7204_),
    .B(_7203_),
    .S(\datapath.idinstr_16_bF$buf7 ),
    .Y(_7205_)
);

NAND2X1 _18157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf10 ),
    .B(_7205_),
    .Y(_7206_)
);

AOI21X1 _18158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7202_),
    .B(_7206_),
    .C(_6145__bF$buf0),
    .Y(_7207_)
);

MUX2X1 _18159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [23]),
    .B(\datapath.registers.1226[16] [23]),
    .S(\datapath.idinstr_16_bF$buf6 ),
    .Y(_7208_)
);

NAND2X1 _18160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf8),
    .B(_7208_),
    .Y(_7209_)
);

MUX2X1 _18161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [23]),
    .B(\datapath.registers.1226[17] [23]),
    .S(\datapath.idinstr_16_bF$buf5 ),
    .Y(_7210_)
);

AOI21X1 _18162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf33 ),
    .B(_7210_),
    .C(\datapath.idinstr_17_bF$buf9 ),
    .Y(_7211_)
);

NAND2X1 _18163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7209_),
    .B(_7211_),
    .Y(_7212_)
);

MUX2X1 _18164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [23]),
    .B(\datapath.registers.1226[20] [23]),
    .S(\datapath.idinstr_16_bF$buf4 ),
    .Y(_7213_)
);

NAND2X1 _18165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf7),
    .B(_7213_),
    .Y(_7214_)
);

MUX2X1 _18166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [23]),
    .B(\datapath.registers.1226[21] [23]),
    .S(\datapath.idinstr_16_bF$buf3 ),
    .Y(_7215_)
);

AOI21X1 _18167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf32 ),
    .B(_7215_),
    .C(_6144__bF$buf10),
    .Y(_7216_)
);

NAND2X1 _18168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7214_),
    .B(_7216_),
    .Y(_7217_)
);

AOI21X1 _18169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7212_),
    .B(_7217_),
    .C(\datapath.idinstr_18_bF$buf5 ),
    .Y(_7218_)
);

OAI21X1 _18170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7207_),
    .B(_7218_),
    .C(\datapath.idinstr_19_bF$buf2 ),
    .Y(_7219_)
);

MUX2X1 _18171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [23]),
    .B(\datapath.registers.1226[8] [23]),
    .S(\datapath.idinstr_15_bF$buf31 ),
    .Y(_7220_)
);

MUX2X1 _18172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [23]),
    .B(\datapath.registers.1226[10] [23]),
    .S(\datapath.idinstr_15_bF$buf30 ),
    .Y(_7221_)
);

MUX2X1 _18173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7221_),
    .B(_7220_),
    .S(\datapath.idinstr_16_bF$buf2 ),
    .Y(_7222_)
);

NAND2X1 _18174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf9),
    .B(_7222_),
    .Y(_7223_)
);

INVX1 _18175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [23]),
    .Y(_7224_)
);

NOR2X1 _18176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7224_),
    .B(_6141__bF$buf6),
    .Y(_7225_)
);

INVX1 _18177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [23]),
    .Y(_7226_)
);

OAI21X1 _18178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7226_),
    .B(\datapath.idinstr_15_bF$buf29 ),
    .C(\datapath.idinstr_16_bF$buf1 ),
    .Y(_7227_)
);

NAND2X1 _18179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [23]),
    .B(_6141__bF$buf5),
    .Y(_7228_)
);

AOI21X1 _18180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [23]),
    .B(\datapath.idinstr_15_bF$buf28 ),
    .C(\datapath.idinstr_16_bF$buf0 ),
    .Y(_7229_)
);

AOI21X1 _18181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7229_),
    .B(_7228_),
    .C(_6144__bF$buf8),
    .Y(_7230_)
);

OAI21X1 _18182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7225_),
    .B(_7227_),
    .C(_7230_),
    .Y(_7231_)
);

AOI21X1 _18183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7231_),
    .B(_7223_),
    .C(_6145__bF$buf7),
    .Y(_7232_)
);

MUX2X1 _18184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [23]),
    .B(\datapath.registers.1226[4] [23]),
    .S(\datapath.idinstr_15_bF$buf27 ),
    .Y(_7233_)
);

MUX2X1 _18185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [23]),
    .B(\datapath.registers.1226[6] [23]),
    .S(\datapath.idinstr_15_bF$buf26 ),
    .Y(_7234_)
);

MUX2X1 _18186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7234_),
    .B(_7233_),
    .S(\datapath.idinstr_16_bF$buf45 ),
    .Y(_7235_)
);

NAND2X1 _18187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf8 ),
    .B(_7235_),
    .Y(_7236_)
);

MUX2X1 _18188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [23]),
    .B(\datapath.registers.1226[0] [23]),
    .S(\datapath.idinstr_15_bF$buf25 ),
    .Y(_7237_)
);

MUX2X1 _18189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [23]),
    .B(\datapath.registers.1226[2] [23]),
    .S(\datapath.idinstr_15_bF$buf24 ),
    .Y(_7238_)
);

MUX2X1 _18190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7238_),
    .B(_7237_),
    .S(\datapath.idinstr_16_bF$buf44 ),
    .Y(_7239_)
);

NAND2X1 _18191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf7),
    .B(_7239_),
    .Y(_7240_)
);

AOI21X1 _18192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7236_),
    .B(_7240_),
    .C(\datapath.idinstr_18_bF$buf4 ),
    .Y(_7241_)
);

OAI21X1 _18193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7241_),
    .B(_7232_),
    .C(_6140__bF$buf0),
    .Y(_7242_)
);

AOI21X1 _18194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7219_),
    .B(_7242_),
    .C(_6147__bF$buf1),
    .Y(\datapath.registers.rega_data [23])
);

MUX2X1 _18195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [24]),
    .B(\datapath.registers.1226[24] [24]),
    .S(\datapath.idinstr_15_bF$buf23 ),
    .Y(_7243_)
);

MUX2X1 _18196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [24]),
    .B(\datapath.registers.1226[26] [24]),
    .S(\datapath.idinstr_15_bF$buf22 ),
    .Y(_7244_)
);

MUX2X1 _18197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7244_),
    .B(_7243_),
    .S(\datapath.idinstr_16_bF$buf43 ),
    .Y(_7245_)
);

NAND2X1 _18198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf6),
    .B(_7245_),
    .Y(_7246_)
);

MUX2X1 _18199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [24]),
    .B(\datapath.registers.1226[28] [24]),
    .S(\datapath.idinstr_15_bF$buf21 ),
    .Y(_7247_)
);

MUX2X1 _18200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [24]),
    .B(\datapath.registers.1226[30] [24]),
    .S(\datapath.idinstr_15_bF$buf20 ),
    .Y(_7248_)
);

MUX2X1 _18201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7248_),
    .B(_7247_),
    .S(\datapath.idinstr_16_bF$buf42 ),
    .Y(_7249_)
);

NAND2X1 _18202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf7 ),
    .B(_7249_),
    .Y(_7250_)
);

AOI21X1 _18203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7246_),
    .B(_7250_),
    .C(_6145__bF$buf6),
    .Y(_7251_)
);

MUX2X1 _18204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [24]),
    .B(\datapath.registers.1226[16] [24]),
    .S(\datapath.idinstr_16_bF$buf41 ),
    .Y(_7252_)
);

NAND2X1 _18205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf4),
    .B(_7252_),
    .Y(_7253_)
);

MUX2X1 _18206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [24]),
    .B(\datapath.registers.1226[17] [24]),
    .S(\datapath.idinstr_16_bF$buf40 ),
    .Y(_7254_)
);

AOI21X1 _18207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf19 ),
    .B(_7254_),
    .C(\datapath.idinstr_17_bF$buf6 ),
    .Y(_7255_)
);

NAND2X1 _18208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7253_),
    .B(_7255_),
    .Y(_7256_)
);

MUX2X1 _18209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [24]),
    .B(\datapath.registers.1226[20] [24]),
    .S(\datapath.idinstr_16_bF$buf39 ),
    .Y(_7257_)
);

NAND2X1 _18210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf3),
    .B(_7257_),
    .Y(_7258_)
);

MUX2X1 _18211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [24]),
    .B(\datapath.registers.1226[21] [24]),
    .S(\datapath.idinstr_16_bF$buf38 ),
    .Y(_7259_)
);

AOI21X1 _18212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf18 ),
    .B(_7259_),
    .C(_6144__bF$buf5),
    .Y(_7260_)
);

NAND2X1 _18213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7258_),
    .B(_7260_),
    .Y(_7261_)
);

AOI21X1 _18214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7256_),
    .B(_7261_),
    .C(\datapath.idinstr_18_bF$buf3 ),
    .Y(_7262_)
);

OAI21X1 _18215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7251_),
    .B(_7262_),
    .C(\datapath.idinstr_19_bF$buf1 ),
    .Y(_7263_)
);

MUX2X1 _18216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [24]),
    .B(\datapath.registers.1226[8] [24]),
    .S(\datapath.idinstr_15_bF$buf17 ),
    .Y(_7264_)
);

MUX2X1 _18217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [24]),
    .B(\datapath.registers.1226[10] [24]),
    .S(\datapath.idinstr_15_bF$buf16 ),
    .Y(_7265_)
);

MUX2X1 _18218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7265_),
    .B(_7264_),
    .S(\datapath.idinstr_16_bF$buf37 ),
    .Y(_7266_)
);

NAND2X1 _18219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf4),
    .B(_7266_),
    .Y(_7267_)
);

AND2X2 _18220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [24]),
    .B(\datapath.idinstr_15_bF$buf15 ),
    .Y(_7268_)
);

INVX1 _18221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [24]),
    .Y(_7269_)
);

OAI21X1 _18222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7269_),
    .B(\datapath.idinstr_15_bF$buf14 ),
    .C(\datapath.idinstr_16_bF$buf36 ),
    .Y(_7270_)
);

NAND2X1 _18223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [24]),
    .B(_6141__bF$buf2),
    .Y(_7271_)
);

AOI21X1 _18224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [24]),
    .B(\datapath.idinstr_15_bF$buf13 ),
    .C(\datapath.idinstr_16_bF$buf35 ),
    .Y(_7272_)
);

AOI21X1 _18225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7272_),
    .B(_7271_),
    .C(_6144__bF$buf3),
    .Y(_7273_)
);

OAI21X1 _18226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7268_),
    .B(_7270_),
    .C(_7273_),
    .Y(_7274_)
);

AOI21X1 _18227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7274_),
    .B(_7267_),
    .C(_6145__bF$buf5),
    .Y(_7275_)
);

MUX2X1 _18228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [24]),
    .B(\datapath.registers.1226[4] [24]),
    .S(\datapath.idinstr_15_bF$buf12 ),
    .Y(_7276_)
);

MUX2X1 _18229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [24]),
    .B(\datapath.registers.1226[6] [24]),
    .S(\datapath.idinstr_15_bF$buf11 ),
    .Y(_7277_)
);

MUX2X1 _18230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7277_),
    .B(_7276_),
    .S(\datapath.idinstr_16_bF$buf34 ),
    .Y(_7278_)
);

NAND2X1 _18231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf5 ),
    .B(_7278_),
    .Y(_7279_)
);

MUX2X1 _18232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [24]),
    .B(\datapath.registers.1226[0] [24]),
    .S(\datapath.idinstr_15_bF$buf10 ),
    .Y(_7280_)
);

MUX2X1 _18233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [24]),
    .B(\datapath.registers.1226[2] [24]),
    .S(\datapath.idinstr_15_bF$buf9 ),
    .Y(_7281_)
);

MUX2X1 _18234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7281_),
    .B(_7280_),
    .S(\datapath.idinstr_16_bF$buf33 ),
    .Y(_7282_)
);

NAND2X1 _18235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf2),
    .B(_7282_),
    .Y(_7283_)
);

AOI21X1 _18236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7279_),
    .B(_7283_),
    .C(\datapath.idinstr_18_bF$buf2 ),
    .Y(_7284_)
);

OAI21X1 _18237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7284_),
    .B(_7275_),
    .C(_6140__bF$buf4),
    .Y(_7285_)
);

AOI21X1 _18238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7263_),
    .B(_7285_),
    .C(_6147__bF$buf0),
    .Y(\datapath.registers.rega_data [24])
);

INVX1 _18239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [25]),
    .Y(_7286_)
);

AOI21X1 _18240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf4 ),
    .B(\datapath.registers.1226[5] [25]),
    .C(_6141__bF$buf1),
    .Y(_7287_)
);

OAI21X1 _18241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf3 ),
    .B(_7286_),
    .C(_7287_),
    .Y(_7288_)
);

INVX1 _18242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [25]),
    .Y(_7289_)
);

AOI21X1 _18243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf2 ),
    .B(\datapath.registers.1226[4] [25]),
    .C(\datapath.idinstr_15_bF$buf8 ),
    .Y(_7290_)
);

OAI21X1 _18244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7289_),
    .B(\datapath.idinstr_17_bF$buf1 ),
    .C(_7290_),
    .Y(_7291_)
);

NAND3X1 _18245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf0),
    .B(_7291_),
    .C(_7288_),
    .Y(_7292_)
);

INVX1 _18246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [25]),
    .Y(_7293_)
);

AOI21X1 _18247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf0 ),
    .B(\datapath.registers.1226[7] [25]),
    .C(_6141__bF$buf0),
    .Y(_7294_)
);

OAI21X1 _18248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf41 ),
    .B(_7293_),
    .C(_7294_),
    .Y(_7295_)
);

INVX1 _18249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[2] [25]),
    .Y(_7296_)
);

AOI21X1 _18250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf40 ),
    .B(\datapath.registers.1226[6] [25]),
    .C(\datapath.idinstr_15_bF$buf7 ),
    .Y(_7297_)
);

OAI21X1 _18251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf39 ),
    .B(_7296_),
    .C(_7297_),
    .Y(_7298_)
);

NAND3X1 _18252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_bF$buf32 ),
    .B(_7298_),
    .C(_7295_),
    .Y(_7299_)
);

AOI21X1 _18253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7292_),
    .B(_7299_),
    .C(\datapath.idinstr_18_bF$buf1 ),
    .Y(_7300_)
);

MUX2X1 _18254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [25]),
    .B(\datapath.registers.1226[8] [25]),
    .S(\datapath.idinstr_15_bF$buf6 ),
    .Y(_7301_)
);

MUX2X1 _18255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [25]),
    .B(\datapath.registers.1226[10] [25]),
    .S(\datapath.idinstr_15_bF$buf5 ),
    .Y(_7302_)
);

MUX2X1 _18256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7302_),
    .B(_7301_),
    .S(\datapath.idinstr_16_bF$buf31 ),
    .Y(_7303_)
);

NAND2X1 _18257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf1),
    .B(_7303_),
    .Y(_7304_)
);

MUX2X1 _18258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [25]),
    .B(\datapath.registers.1226[12] [25]),
    .S(\datapath.idinstr_15_bF$buf4 ),
    .Y(_7305_)
);

MUX2X1 _18259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [25]),
    .B(\datapath.registers.1226[14] [25]),
    .S(\datapath.idinstr_15_bF$buf3 ),
    .Y(_7306_)
);

MUX2X1 _18260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7306_),
    .B(_7305_),
    .S(\datapath.idinstr_16_bF$buf30 ),
    .Y(_7307_)
);

NAND2X1 _18261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf38 ),
    .B(_7307_),
    .Y(_7308_)
);

AOI21X1 _18262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7304_),
    .B(_7308_),
    .C(_6145__bF$buf4),
    .Y(_7309_)
);

OAI21X1 _18263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7309_),
    .B(_7300_),
    .C(_6140__bF$buf3),
    .Y(_7310_)
);

MUX2X1 _18264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [25]),
    .B(\datapath.registers.1226[16] [25]),
    .S(\datapath.idinstr_15_bF$buf2 ),
    .Y(_7311_)
);

MUX2X1 _18265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [25]),
    .B(\datapath.registers.1226[18] [25]),
    .S(\datapath.idinstr_15_bF$buf1 ),
    .Y(_7312_)
);

MUX2X1 _18266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7312_),
    .B(_7311_),
    .S(\datapath.idinstr_16_bF$buf29 ),
    .Y(_7313_)
);

NAND2X1 _18267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf0),
    .B(_7313_),
    .Y(_7314_)
);

MUX2X1 _18268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [25]),
    .B(\datapath.registers.1226[20] [25]),
    .S(\datapath.idinstr_15_bF$buf0 ),
    .Y(_7315_)
);

MUX2X1 _18269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [25]),
    .B(\datapath.registers.1226[22] [25]),
    .S(\datapath.idinstr_15_bF$buf53 ),
    .Y(_7316_)
);

MUX2X1 _18270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7316_),
    .B(_7315_),
    .S(\datapath.idinstr_16_bF$buf28 ),
    .Y(_7317_)
);

NAND2X1 _18271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf37 ),
    .B(_7317_),
    .Y(_7318_)
);

AOI21X1 _18272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7314_),
    .B(_7318_),
    .C(\datapath.idinstr_18_bF$buf0 ),
    .Y(_7319_)
);

INVX1 _18273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [25]),
    .Y(_7320_)
);

AOI21X1 _18274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [25]),
    .B(\datapath.idinstr_17_bF$buf36 ),
    .C(_6141__bF$buf10),
    .Y(_7321_)
);

OAI21X1 _18275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7320_),
    .B(\datapath.idinstr_17_bF$buf35 ),
    .C(_7321_),
    .Y(_7322_)
);

NAND2X1 _18276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [25]),
    .B(_6144__bF$buf10),
    .Y(_7323_)
);

AOI21X1 _18277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [25]),
    .B(\datapath.idinstr_17_bF$buf34 ),
    .C(\datapath.idinstr_15_bF$buf52 ),
    .Y(_7324_)
);

AOI21X1 _18278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7324_),
    .B(_7323_),
    .C(_6143__bF$buf4),
    .Y(_7325_)
);

NAND2X1 _18279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7322_),
    .B(_7325_),
    .Y(_7326_)
);

INVX1 _18280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [25]),
    .Y(_7327_)
);

AOI21X1 _18281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [25]),
    .B(\datapath.idinstr_17_bF$buf33 ),
    .C(_6141__bF$buf9),
    .Y(_7328_)
);

OAI21X1 _18282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7327_),
    .B(\datapath.idinstr_17_bF$buf32 ),
    .C(_7328_),
    .Y(_7329_)
);

AOI21X1 _18283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[28] [25]),
    .B(\datapath.idinstr_17_bF$buf31 ),
    .C(\datapath.idinstr_15_bF$buf51 ),
    .Y(_7330_)
);

OAI21X1 _18284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5747_),
    .B(\datapath.idinstr_17_bF$buf30 ),
    .C(_7330_),
    .Y(_7331_)
);

NAND3X1 _18285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf3),
    .B(_7331_),
    .C(_7329_),
    .Y(_7332_)
);

AOI21X1 _18286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7326_),
    .B(_7332_),
    .C(_6145__bF$buf3),
    .Y(_7333_)
);

OAI21X1 _18287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7319_),
    .B(_7333_),
    .C(\datapath.idinstr_19_bF$buf0 ),
    .Y(_7334_)
);

AOI21X1 _18288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7334_),
    .B(_7310_),
    .C(_6147__bF$buf4),
    .Y(\datapath.registers.rega_data [25])
);

MUX2X1 _18289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [26]),
    .B(\datapath.registers.1226[24] [26]),
    .S(\datapath.idinstr_15_bF$buf50 ),
    .Y(_7335_)
);

MUX2X1 _18290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [26]),
    .B(\datapath.registers.1226[26] [26]),
    .S(\datapath.idinstr_15_bF$buf49 ),
    .Y(_7336_)
);

MUX2X1 _18291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7336_),
    .B(_7335_),
    .S(\datapath.idinstr_16_bF$buf27 ),
    .Y(_7337_)
);

NAND2X1 _18292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf9),
    .B(_7337_),
    .Y(_7338_)
);

MUX2X1 _18293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [26]),
    .B(\datapath.registers.1226[28] [26]),
    .S(\datapath.idinstr_15_bF$buf48 ),
    .Y(_7339_)
);

MUX2X1 _18294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [26]),
    .B(\datapath.registers.1226[30] [26]),
    .S(\datapath.idinstr_15_bF$buf47 ),
    .Y(_7340_)
);

MUX2X1 _18295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7340_),
    .B(_7339_),
    .S(\datapath.idinstr_16_bF$buf26 ),
    .Y(_7341_)
);

NAND2X1 _18296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf29 ),
    .B(_7341_),
    .Y(_7342_)
);

AOI21X1 _18297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7338_),
    .B(_7342_),
    .C(_6145__bF$buf2),
    .Y(_7343_)
);

MUX2X1 _18298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [26]),
    .B(\datapath.registers.1226[16] [26]),
    .S(\datapath.idinstr_16_bF$buf25 ),
    .Y(_7344_)
);

NAND2X1 _18299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf8),
    .B(_7344_),
    .Y(_7345_)
);

MUX2X1 _18300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [26]),
    .B(\datapath.registers.1226[17] [26]),
    .S(\datapath.idinstr_16_bF$buf24 ),
    .Y(_7346_)
);

AOI21X1 _18301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf46 ),
    .B(_7346_),
    .C(\datapath.idinstr_17_bF$buf28 ),
    .Y(_7347_)
);

NAND2X1 _18302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7345_),
    .B(_7347_),
    .Y(_7348_)
);

MUX2X1 _18303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [26]),
    .B(\datapath.registers.1226[20] [26]),
    .S(\datapath.idinstr_16_bF$buf23 ),
    .Y(_7349_)
);

NAND2X1 _18304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf7),
    .B(_7349_),
    .Y(_7350_)
);

MUX2X1 _18305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [26]),
    .B(\datapath.registers.1226[21] [26]),
    .S(\datapath.idinstr_16_bF$buf22 ),
    .Y(_7351_)
);

AOI21X1 _18306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf45 ),
    .B(_7351_),
    .C(_6144__bF$buf8),
    .Y(_7352_)
);

NAND2X1 _18307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7350_),
    .B(_7352_),
    .Y(_7353_)
);

AOI21X1 _18308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7348_),
    .B(_7353_),
    .C(\datapath.idinstr_18_bF$buf7 ),
    .Y(_7354_)
);

OAI21X1 _18309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7343_),
    .B(_7354_),
    .C(\datapath.idinstr_19_bF$buf5 ),
    .Y(_7355_)
);

MUX2X1 _18310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [26]),
    .B(\datapath.registers.1226[8] [26]),
    .S(\datapath.idinstr_15_bF$buf44 ),
    .Y(_7356_)
);

MUX2X1 _18311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [26]),
    .B(\datapath.registers.1226[10] [26]),
    .S(\datapath.idinstr_15_bF$buf43 ),
    .Y(_7357_)
);

MUX2X1 _18312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7357_),
    .B(_7356_),
    .S(\datapath.idinstr_16_bF$buf21 ),
    .Y(_7358_)
);

NAND2X1 _18313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf7),
    .B(_7358_),
    .Y(_7359_)
);

INVX1 _18314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [26]),
    .Y(_7360_)
);

NOR2X1 _18315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7360_),
    .B(_6141__bF$buf6),
    .Y(_7361_)
);

INVX1 _18316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [26]),
    .Y(_7362_)
);

OAI21X1 _18317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7362_),
    .B(\datapath.idinstr_15_bF$buf42 ),
    .C(\datapath.idinstr_16_bF$buf20 ),
    .Y(_7363_)
);

NAND2X1 _18318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [26]),
    .B(_6141__bF$buf5),
    .Y(_7364_)
);

AOI21X1 _18319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [26]),
    .B(\datapath.idinstr_15_bF$buf41 ),
    .C(\datapath.idinstr_16_bF$buf19 ),
    .Y(_7365_)
);

AOI21X1 _18320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7365_),
    .B(_7364_),
    .C(_6144__bF$buf6),
    .Y(_7366_)
);

OAI21X1 _18321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7361_),
    .B(_7363_),
    .C(_7366_),
    .Y(_7367_)
);

AOI21X1 _18322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7367_),
    .B(_7359_),
    .C(_6145__bF$buf1),
    .Y(_7368_)
);

MUX2X1 _18323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [26]),
    .B(\datapath.registers.1226[4] [26]),
    .S(\datapath.idinstr_15_bF$buf40 ),
    .Y(_7369_)
);

MUX2X1 _18324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [26]),
    .B(\datapath.registers.1226[6] [26]),
    .S(\datapath.idinstr_15_bF$buf39 ),
    .Y(_7370_)
);

MUX2X1 _18325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7370_),
    .B(_7369_),
    .S(\datapath.idinstr_16_bF$buf18 ),
    .Y(_7371_)
);

NAND2X1 _18326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf27 ),
    .B(_7371_),
    .Y(_7372_)
);

MUX2X1 _18327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [26]),
    .B(\datapath.registers.1226[0] [26]),
    .S(\datapath.idinstr_15_bF$buf38 ),
    .Y(_7373_)
);

MUX2X1 _18328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [26]),
    .B(\datapath.registers.1226[2] [26]),
    .S(\datapath.idinstr_15_bF$buf37 ),
    .Y(_7374_)
);

MUX2X1 _18329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7374_),
    .B(_7373_),
    .S(\datapath.idinstr_16_bF$buf17 ),
    .Y(_7375_)
);

NAND2X1 _18330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf5),
    .B(_7375_),
    .Y(_7376_)
);

AOI21X1 _18331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7372_),
    .B(_7376_),
    .C(\datapath.idinstr_18_bF$buf6 ),
    .Y(_7377_)
);

OAI21X1 _18332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7377_),
    .B(_7368_),
    .C(_6140__bF$buf2),
    .Y(_7378_)
);

AOI21X1 _18333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7355_),
    .B(_7378_),
    .C(_6147__bF$buf3),
    .Y(\datapath.registers.rega_data [26])
);

MUX2X1 _18334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [27]),
    .B(\datapath.registers.1226[8] [27]),
    .S(\datapath.idinstr_15_bF$buf36 ),
    .Y(_7379_)
);

MUX2X1 _18335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [27]),
    .B(\datapath.registers.1226[10] [27]),
    .S(\datapath.idinstr_15_bF$buf35 ),
    .Y(_7380_)
);

MUX2X1 _18336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7380_),
    .B(_7379_),
    .S(\datapath.idinstr_16_bF$buf16 ),
    .Y(_7381_)
);

NAND2X1 _18337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf4),
    .B(_7381_),
    .Y(_7382_)
);

MUX2X1 _18338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [27]),
    .B(\datapath.registers.1226[12] [27]),
    .S(\datapath.idinstr_15_bF$buf34 ),
    .Y(_7383_)
);

MUX2X1 _18339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [27]),
    .B(\datapath.registers.1226[14] [27]),
    .S(\datapath.idinstr_15_bF$buf33 ),
    .Y(_7384_)
);

MUX2X1 _18340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7384_),
    .B(_7383_),
    .S(\datapath.idinstr_16_bF$buf15 ),
    .Y(_7385_)
);

NAND2X1 _18341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf26 ),
    .B(_7385_),
    .Y(_7386_)
);

AOI21X1 _18342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7382_),
    .B(_7386_),
    .C(_6145__bF$buf0),
    .Y(_7387_)
);

INVX1 _18343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [27]),
    .Y(_7388_)
);

AOI21X1 _18344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf25 ),
    .B(\datapath.registers.1226[5] [27]),
    .C(_6141__bF$buf4),
    .Y(_7389_)
);

OAI21X1 _18345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf24 ),
    .B(_7388_),
    .C(_7389_),
    .Y(_7390_)
);

NAND2X1 _18346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [27]),
    .B(_6144__bF$buf3),
    .Y(_7391_)
);

AOI21X1 _18347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf23 ),
    .B(\datapath.registers.1226[4] [27]),
    .C(\datapath.idinstr_15_bF$buf32 ),
    .Y(_7392_)
);

AOI21X1 _18348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7392_),
    .B(_7391_),
    .C(\datapath.idinstr_16_bF$buf14 ),
    .Y(_7393_)
);

NAND2X1 _18349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7390_),
    .B(_7393_),
    .Y(_7394_)
);

INVX1 _18350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [27]),
    .Y(_7395_)
);

AOI21X1 _18351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf22 ),
    .B(\datapath.registers.1226[7] [27]),
    .C(_6141__bF$buf3),
    .Y(_7396_)
);

OAI21X1 _18352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf21 ),
    .B(_7395_),
    .C(_7396_),
    .Y(_7397_)
);

INVX1 _18353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[2] [27]),
    .Y(_7398_)
);

AOI21X1 _18354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf20 ),
    .B(\datapath.registers.1226[6] [27]),
    .C(\datapath.idinstr_15_bF$buf31 ),
    .Y(_7399_)
);

OAI21X1 _18355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf19 ),
    .B(_7398_),
    .C(_7399_),
    .Y(_7400_)
);

NAND3X1 _18356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_bF$buf13 ),
    .B(_7400_),
    .C(_7397_),
    .Y(_7401_)
);

AOI21X1 _18357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7394_),
    .B(_7401_),
    .C(\datapath.idinstr_18_bF$buf5 ),
    .Y(_7402_)
);

OAI21X1 _18358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7387_),
    .B(_7402_),
    .C(_6140__bF$buf1),
    .Y(_7403_)
);

MUX2X1 _18359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [27]),
    .B(\datapath.registers.1226[29] [27]),
    .S(\datapath.idinstr_16_bF$buf12 ),
    .Y(_7404_)
);

MUX2X1 _18360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [27]),
    .B(\datapath.registers.1226[28] [27]),
    .S(\datapath.idinstr_16_bF$buf11 ),
    .Y(_7405_)
);

MUX2X1 _18361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7405_),
    .B(_7404_),
    .S(_6141__bF$buf2),
    .Y(_7406_)
);

NAND2X1 _18362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf18 ),
    .B(_7406_),
    .Y(_7407_)
);

MUX2X1 _18363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [27]),
    .B(\datapath.registers.1226[25] [27]),
    .S(\datapath.idinstr_16_bF$buf10 ),
    .Y(_7408_)
);

MUX2X1 _18364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [27]),
    .B(\datapath.registers.1226[24] [27]),
    .S(\datapath.idinstr_16_bF$buf9 ),
    .Y(_7409_)
);

MUX2X1 _18365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7409_),
    .B(_7408_),
    .S(_6141__bF$buf1),
    .Y(_7410_)
);

NAND2X1 _18366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf2),
    .B(_7410_),
    .Y(_7411_)
);

AOI21X1 _18367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7407_),
    .B(_7411_),
    .C(_6145__bF$buf7),
    .Y(_7412_)
);

INVX1 _18368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [27]),
    .Y(_7413_)
);

AOI21X1 _18369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [27]),
    .B(\datapath.idinstr_17_bF$buf17 ),
    .C(_6141__bF$buf0),
    .Y(_7414_)
);

OAI21X1 _18370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7413_),
    .B(\datapath.idinstr_17_bF$buf16 ),
    .C(_7414_),
    .Y(_7415_)
);

INVX1 _18371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [27]),
    .Y(_7416_)
);

AOI21X1 _18372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [27]),
    .B(\datapath.idinstr_17_bF$buf15 ),
    .C(\datapath.idinstr_15_bF$buf30 ),
    .Y(_7417_)
);

OAI21X1 _18373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7416_),
    .B(\datapath.idinstr_17_bF$buf14 ),
    .C(_7417_),
    .Y(_7418_)
);

NAND3X1 _18374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_bF$buf8 ),
    .B(_7418_),
    .C(_7415_),
    .Y(_7419_)
);

INVX1 _18375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [27]),
    .Y(_7420_)
);

AOI21X1 _18376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [27]),
    .B(\datapath.idinstr_17_bF$buf13 ),
    .C(_6141__bF$buf10),
    .Y(_7421_)
);

OAI21X1 _18377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7420_),
    .B(\datapath.idinstr_17_bF$buf12 ),
    .C(_7421_),
    .Y(_7422_)
);

AOI21X1 _18378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [27]),
    .B(\datapath.idinstr_17_bF$buf11 ),
    .C(\datapath.idinstr_15_bF$buf29 ),
    .Y(_7423_)
);

OAI21X1 _18379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6032_),
    .B(\datapath.idinstr_17_bF$buf10 ),
    .C(_7423_),
    .Y(_7424_)
);

NAND3X1 _18380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf2),
    .B(_7424_),
    .C(_7422_),
    .Y(_7425_)
);

AOI21X1 _18381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7419_),
    .B(_7425_),
    .C(\datapath.idinstr_18_bF$buf4 ),
    .Y(_7426_)
);

OAI21X1 _18382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7412_),
    .B(_7426_),
    .C(\datapath.idinstr_19_bF$buf4 ),
    .Y(_7427_)
);

AOI21X1 _18383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7403_),
    .B(_7427_),
    .C(_6147__bF$buf2),
    .Y(\datapath.registers.rega_data [27])
);

MUX2X1 _18384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [28]),
    .B(\datapath.registers.1226[24] [28]),
    .S(\datapath.idinstr_15_bF$buf28 ),
    .Y(_7428_)
);

MUX2X1 _18385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [28]),
    .B(\datapath.registers.1226[26] [28]),
    .S(\datapath.idinstr_15_bF$buf27 ),
    .Y(_7429_)
);

MUX2X1 _18386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7429_),
    .B(_7428_),
    .S(\datapath.idinstr_16_bF$buf7 ),
    .Y(_7430_)
);

NAND2X1 _18387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf1),
    .B(_7430_),
    .Y(_7431_)
);

MUX2X1 _18388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [28]),
    .B(\datapath.registers.1226[28] [28]),
    .S(\datapath.idinstr_15_bF$buf26 ),
    .Y(_7432_)
);

MUX2X1 _18389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [28]),
    .B(\datapath.registers.1226[30] [28]),
    .S(\datapath.idinstr_15_bF$buf25 ),
    .Y(_7433_)
);

MUX2X1 _18390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7433_),
    .B(_7432_),
    .S(\datapath.idinstr_16_bF$buf6 ),
    .Y(_7434_)
);

NAND2X1 _18391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf9 ),
    .B(_7434_),
    .Y(_7435_)
);

AOI21X1 _18392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7431_),
    .B(_7435_),
    .C(_6145__bF$buf6),
    .Y(_7436_)
);

MUX2X1 _18393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [28]),
    .B(\datapath.registers.1226[16] [28]),
    .S(\datapath.idinstr_16_bF$buf5 ),
    .Y(_7437_)
);

NAND2X1 _18394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf9),
    .B(_7437_),
    .Y(_7438_)
);

MUX2X1 _18395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [28]),
    .B(\datapath.registers.1226[17] [28]),
    .S(\datapath.idinstr_16_bF$buf4 ),
    .Y(_7439_)
);

AOI21X1 _18396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf24 ),
    .B(_7439_),
    .C(\datapath.idinstr_17_bF$buf8 ),
    .Y(_7440_)
);

NAND2X1 _18397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7438_),
    .B(_7440_),
    .Y(_7441_)
);

MUX2X1 _18398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [28]),
    .B(\datapath.registers.1226[20] [28]),
    .S(\datapath.idinstr_16_bF$buf3 ),
    .Y(_7442_)
);

NAND2X1 _18399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf8),
    .B(_7442_),
    .Y(_7443_)
);

MUX2X1 _18400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [28]),
    .B(\datapath.registers.1226[21] [28]),
    .S(\datapath.idinstr_16_bF$buf2 ),
    .Y(_7444_)
);

AOI21X1 _18401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf23 ),
    .B(_7444_),
    .C(_6144__bF$buf0),
    .Y(_7445_)
);

NAND2X1 _18402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7443_),
    .B(_7445_),
    .Y(_7446_)
);

AOI21X1 _18403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7441_),
    .B(_7446_),
    .C(\datapath.idinstr_18_bF$buf3 ),
    .Y(_7447_)
);

OAI21X1 _18404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7436_),
    .B(_7447_),
    .C(\datapath.idinstr_19_bF$buf3 ),
    .Y(_7448_)
);

MUX2X1 _18405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [28]),
    .B(\datapath.registers.1226[8] [28]),
    .S(\datapath.idinstr_15_bF$buf22 ),
    .Y(_7449_)
);

MUX2X1 _18406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [28]),
    .B(\datapath.registers.1226[10] [28]),
    .S(\datapath.idinstr_15_bF$buf21 ),
    .Y(_7450_)
);

MUX2X1 _18407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7450_),
    .B(_7449_),
    .S(\datapath.idinstr_16_bF$buf1 ),
    .Y(_7451_)
);

NAND2X1 _18408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf10),
    .B(_7451_),
    .Y(_7452_)
);

MUX2X1 _18409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [28]),
    .B(\datapath.registers.1226[12] [28]),
    .S(\datapath.idinstr_15_bF$buf20 ),
    .Y(_7453_)
);

MUX2X1 _18410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [28]),
    .B(\datapath.registers.1226[14] [28]),
    .S(\datapath.idinstr_15_bF$buf19 ),
    .Y(_7454_)
);

MUX2X1 _18411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7454_),
    .B(_7453_),
    .S(\datapath.idinstr_16_bF$buf0 ),
    .Y(_7455_)
);

NAND2X1 _18412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf7 ),
    .B(_7455_),
    .Y(_7456_)
);

AOI21X1 _18413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7452_),
    .B(_7456_),
    .C(_6145__bF$buf5),
    .Y(_7457_)
);

INVX1 _18414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [28]),
    .Y(_7458_)
);

AOI21X1 _18415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf6 ),
    .B(\datapath.registers.1226[5] [28]),
    .C(_6141__bF$buf7),
    .Y(_7459_)
);

OAI21X1 _18416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf5 ),
    .B(_7458_),
    .C(_7459_),
    .Y(_7460_)
);

INVX1 _18417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [28]),
    .Y(_7461_)
);

AOI21X1 _18418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf4 ),
    .B(\datapath.registers.1226[4] [28]),
    .C(\datapath.idinstr_15_bF$buf18 ),
    .Y(_7462_)
);

OAI21X1 _18419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7461_),
    .B(\datapath.idinstr_17_bF$buf3 ),
    .C(_7462_),
    .Y(_7463_)
);

NAND3X1 _18420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf1),
    .B(_7463_),
    .C(_7460_),
    .Y(_7464_)
);

INVX1 _18421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [28]),
    .Y(_7465_)
);

AOI21X1 _18422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf2 ),
    .B(\datapath.registers.1226[7] [28]),
    .C(_6141__bF$buf6),
    .Y(_7466_)
);

OAI21X1 _18423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf1 ),
    .B(_7465_),
    .C(_7466_),
    .Y(_7467_)
);

INVX1 _18424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[2] [28]),
    .Y(_7468_)
);

AOI21X1 _18425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf0 ),
    .B(\datapath.registers.1226[6] [28]),
    .C(\datapath.idinstr_15_bF$buf17 ),
    .Y(_7469_)
);

OAI21X1 _18426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf41 ),
    .B(_7468_),
    .C(_7469_),
    .Y(_7470_)
);

NAND3X1 _18427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_bF$buf45 ),
    .B(_7470_),
    .C(_7467_),
    .Y(_7471_)
);

AOI21X1 _18428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7464_),
    .B(_7471_),
    .C(\datapath.idinstr_18_bF$buf2 ),
    .Y(_7472_)
);

OAI21X1 _18429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7457_),
    .B(_7472_),
    .C(_6140__bF$buf0),
    .Y(_7473_)
);

AOI21X1 _18430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7448_),
    .B(_7473_),
    .C(_6147__bF$buf1),
    .Y(\datapath.registers.rega_data [28])
);

MUX2X1 _18431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [29]),
    .B(\datapath.registers.1226[24] [29]),
    .S(\datapath.idinstr_15_bF$buf16 ),
    .Y(_7474_)
);

MUX2X1 _18432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [29]),
    .B(\datapath.registers.1226[26] [29]),
    .S(\datapath.idinstr_15_bF$buf15 ),
    .Y(_7475_)
);

MUX2X1 _18433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7475_),
    .B(_7474_),
    .S(\datapath.idinstr_16_bF$buf44 ),
    .Y(_7476_)
);

NAND2X1 _18434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf9),
    .B(_7476_),
    .Y(_7477_)
);

MUX2X1 _18435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [29]),
    .B(\datapath.registers.1226[28] [29]),
    .S(\datapath.idinstr_15_bF$buf14 ),
    .Y(_7478_)
);

MUX2X1 _18436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [29]),
    .B(\datapath.registers.1226[30] [29]),
    .S(\datapath.idinstr_15_bF$buf13 ),
    .Y(_7479_)
);

MUX2X1 _18437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7479_),
    .B(_7478_),
    .S(\datapath.idinstr_16_bF$buf43 ),
    .Y(_7480_)
);

NAND2X1 _18438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf40 ),
    .B(_7480_),
    .Y(_7481_)
);

AOI21X1 _18439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7477_),
    .B(_7481_),
    .C(_6145__bF$buf4),
    .Y(_7482_)
);

MUX2X1 _18440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [29]),
    .B(\datapath.registers.1226[16] [29]),
    .S(\datapath.idinstr_16_bF$buf42 ),
    .Y(_7483_)
);

NAND2X1 _18441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf5),
    .B(_7483_),
    .Y(_7484_)
);

MUX2X1 _18442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [29]),
    .B(\datapath.registers.1226[17] [29]),
    .S(\datapath.idinstr_16_bF$buf41 ),
    .Y(_7485_)
);

AOI21X1 _18443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf12 ),
    .B(_7485_),
    .C(\datapath.idinstr_17_bF$buf39 ),
    .Y(_7486_)
);

NAND2X1 _18444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7484_),
    .B(_7486_),
    .Y(_7487_)
);

MUX2X1 _18445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [29]),
    .B(\datapath.registers.1226[20] [29]),
    .S(\datapath.idinstr_16_bF$buf40 ),
    .Y(_7488_)
);

NAND2X1 _18446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf4),
    .B(_7488_),
    .Y(_7489_)
);

MUX2X1 _18447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [29]),
    .B(\datapath.registers.1226[21] [29]),
    .S(\datapath.idinstr_16_bF$buf39 ),
    .Y(_7490_)
);

AOI21X1 _18448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf11 ),
    .B(_7490_),
    .C(_6144__bF$buf8),
    .Y(_7491_)
);

NAND2X1 _18449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7489_),
    .B(_7491_),
    .Y(_7492_)
);

AOI21X1 _18450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7487_),
    .B(_7492_),
    .C(\datapath.idinstr_18_bF$buf1 ),
    .Y(_7493_)
);

OAI21X1 _18451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7482_),
    .B(_7493_),
    .C(\datapath.idinstr_19_bF$buf2 ),
    .Y(_7494_)
);

MUX2X1 _18452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [29]),
    .B(\datapath.registers.1226[8] [29]),
    .S(\datapath.idinstr_15_bF$buf10 ),
    .Y(_7495_)
);

MUX2X1 _18453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [29]),
    .B(\datapath.registers.1226[10] [29]),
    .S(\datapath.idinstr_15_bF$buf9 ),
    .Y(_7496_)
);

MUX2X1 _18454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7496_),
    .B(_7495_),
    .S(\datapath.idinstr_16_bF$buf38 ),
    .Y(_7497_)
);

NAND2X1 _18455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf7),
    .B(_7497_),
    .Y(_7498_)
);

AND2X2 _18456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [29]),
    .B(\datapath.idinstr_15_bF$buf8 ),
    .Y(_7499_)
);

INVX1 _18457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [29]),
    .Y(_7500_)
);

OAI21X1 _18458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7500_),
    .B(\datapath.idinstr_15_bF$buf7 ),
    .C(\datapath.idinstr_16_bF$buf37 ),
    .Y(_7501_)
);

NAND2X1 _18459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [29]),
    .B(_6141__bF$buf3),
    .Y(_7502_)
);

AOI21X1 _18460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [29]),
    .B(\datapath.idinstr_15_bF$buf6 ),
    .C(\datapath.idinstr_16_bF$buf36 ),
    .Y(_7503_)
);

AOI21X1 _18461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7503_),
    .B(_7502_),
    .C(_6144__bF$buf6),
    .Y(_7504_)
);

OAI21X1 _18462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7499_),
    .B(_7501_),
    .C(_7504_),
    .Y(_7505_)
);

AOI21X1 _18463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7505_),
    .B(_7498_),
    .C(_6145__bF$buf3),
    .Y(_7506_)
);

MUX2X1 _18464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [29]),
    .B(\datapath.registers.1226[4] [29]),
    .S(\datapath.idinstr_15_bF$buf5 ),
    .Y(_7507_)
);

MUX2X1 _18465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [29]),
    .B(\datapath.registers.1226[6] [29]),
    .S(\datapath.idinstr_15_bF$buf4 ),
    .Y(_7508_)
);

MUX2X1 _18466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7508_),
    .B(_7507_),
    .S(\datapath.idinstr_16_bF$buf35 ),
    .Y(_7509_)
);

NAND2X1 _18467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf38 ),
    .B(_7509_),
    .Y(_7510_)
);

MUX2X1 _18468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [29]),
    .B(\datapath.registers.1226[0] [29]),
    .S(\datapath.idinstr_15_bF$buf3 ),
    .Y(_7511_)
);

MUX2X1 _18469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [29]),
    .B(\datapath.registers.1226[2] [29]),
    .S(\datapath.idinstr_15_bF$buf2 ),
    .Y(_7512_)
);

MUX2X1 _18470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7512_),
    .B(_7511_),
    .S(\datapath.idinstr_16_bF$buf34 ),
    .Y(_7513_)
);

NAND2X1 _18471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf5),
    .B(_7513_),
    .Y(_7514_)
);

AOI21X1 _18472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7510_),
    .B(_7514_),
    .C(\datapath.idinstr_18_bF$buf0 ),
    .Y(_7515_)
);

OAI21X1 _18473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7515_),
    .B(_7506_),
    .C(_6140__bF$buf4),
    .Y(_7516_)
);

AOI21X1 _18474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7494_),
    .B(_7516_),
    .C(_6147__bF$buf0),
    .Y(\datapath.registers.rega_data [29])
);

MUX2X1 _18475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [30]),
    .B(\datapath.registers.1226[24] [30]),
    .S(\datapath.idinstr_15_bF$buf1 ),
    .Y(_7517_)
);

MUX2X1 _18476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [30]),
    .B(\datapath.registers.1226[26] [30]),
    .S(\datapath.idinstr_15_bF$buf0 ),
    .Y(_7518_)
);

MUX2X1 _18477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7518_),
    .B(_7517_),
    .S(\datapath.idinstr_16_bF$buf33 ),
    .Y(_7519_)
);

NAND2X1 _18478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf4),
    .B(_7519_),
    .Y(_7520_)
);

MUX2X1 _18479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [30]),
    .B(\datapath.registers.1226[28] [30]),
    .S(\datapath.idinstr_15_bF$buf53 ),
    .Y(_7521_)
);

MUX2X1 _18480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [30]),
    .B(\datapath.registers.1226[30] [30]),
    .S(\datapath.idinstr_15_bF$buf52 ),
    .Y(_7522_)
);

MUX2X1 _18481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7522_),
    .B(_7521_),
    .S(\datapath.idinstr_16_bF$buf32 ),
    .Y(_7523_)
);

NAND2X1 _18482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf37 ),
    .B(_7523_),
    .Y(_7524_)
);

AOI21X1 _18483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7520_),
    .B(_7524_),
    .C(_6145__bF$buf2),
    .Y(_7525_)
);

MUX2X1 _18484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [30]),
    .B(\datapath.registers.1226[16] [30]),
    .S(\datapath.idinstr_16_bF$buf31 ),
    .Y(_7526_)
);

NAND2X1 _18485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf2),
    .B(_7526_),
    .Y(_7527_)
);

MUX2X1 _18486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [30]),
    .B(\datapath.registers.1226[17] [30]),
    .S(\datapath.idinstr_16_bF$buf30 ),
    .Y(_7528_)
);

AOI21X1 _18487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf51 ),
    .B(_7528_),
    .C(\datapath.idinstr_17_bF$buf36 ),
    .Y(_7529_)
);

NAND2X1 _18488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7527_),
    .B(_7529_),
    .Y(_7530_)
);

MUX2X1 _18489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [30]),
    .B(\datapath.registers.1226[20] [30]),
    .S(\datapath.idinstr_16_bF$buf29 ),
    .Y(_7531_)
);

NAND2X1 _18490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf1),
    .B(_7531_),
    .Y(_7532_)
);

MUX2X1 _18491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [30]),
    .B(\datapath.registers.1226[21] [30]),
    .S(\datapath.idinstr_16_bF$buf28 ),
    .Y(_7533_)
);

AOI21X1 _18492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf50 ),
    .B(_7533_),
    .C(_6144__bF$buf3),
    .Y(_7534_)
);

NAND2X1 _18493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7532_),
    .B(_7534_),
    .Y(_7535_)
);

AOI21X1 _18494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7530_),
    .B(_7535_),
    .C(\datapath.idinstr_18_bF$buf7 ),
    .Y(_7536_)
);

OAI21X1 _18495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7525_),
    .B(_7536_),
    .C(\datapath.idinstr_19_bF$buf1 ),
    .Y(_7537_)
);

MUX2X1 _18496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [30]),
    .B(\datapath.registers.1226[8] [30]),
    .S(\datapath.idinstr_15_bF$buf49 ),
    .Y(_7538_)
);

MUX2X1 _18497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [30]),
    .B(\datapath.registers.1226[10] [30]),
    .S(\datapath.idinstr_15_bF$buf48 ),
    .Y(_7539_)
);

MUX2X1 _18498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7539_),
    .B(_7538_),
    .S(\datapath.idinstr_16_bF$buf27 ),
    .Y(_7540_)
);

NAND2X1 _18499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf2),
    .B(_7540_),
    .Y(_7541_)
);

MUX2X1 _18500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [30]),
    .B(\datapath.registers.1226[12] [30]),
    .S(\datapath.idinstr_15_bF$buf47 ),
    .Y(_7542_)
);

MUX2X1 _18501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [30]),
    .B(\datapath.registers.1226[14] [30]),
    .S(\datapath.idinstr_15_bF$buf46 ),
    .Y(_7543_)
);

MUX2X1 _18502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7543_),
    .B(_7542_),
    .S(\datapath.idinstr_16_bF$buf26 ),
    .Y(_7544_)
);

NAND2X1 _18503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf35 ),
    .B(_7544_),
    .Y(_7545_)
);

AOI21X1 _18504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7541_),
    .B(_7545_),
    .C(_6145__bF$buf1),
    .Y(_7546_)
);

INVX1 _18505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [30]),
    .Y(_7547_)
);

AOI21X1 _18506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf34 ),
    .B(\datapath.registers.1226[5] [30]),
    .C(_6141__bF$buf0),
    .Y(_7548_)
);

OAI21X1 _18507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf33 ),
    .B(_7547_),
    .C(_7548_),
    .Y(_7549_)
);

INVX1 _18508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [30]),
    .Y(_7550_)
);

AOI21X1 _18509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf32 ),
    .B(\datapath.registers.1226[4] [30]),
    .C(\datapath.idinstr_15_bF$buf45 ),
    .Y(_7551_)
);

OAI21X1 _18510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7550_),
    .B(\datapath.idinstr_17_bF$buf31 ),
    .C(_7551_),
    .Y(_7552_)
);

NAND3X1 _18511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143__bF$buf0),
    .B(_7552_),
    .C(_7549_),
    .Y(_7553_)
);

INVX1 _18512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [30]),
    .Y(_7554_)
);

AOI21X1 _18513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf30 ),
    .B(\datapath.registers.1226[7] [30]),
    .C(_6141__bF$buf10),
    .Y(_7555_)
);

OAI21X1 _18514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf29 ),
    .B(_7554_),
    .C(_7555_),
    .Y(_7556_)
);

INVX1 _18515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[2] [30]),
    .Y(_7557_)
);

AOI21X1 _18516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf28 ),
    .B(\datapath.registers.1226[6] [30]),
    .C(\datapath.idinstr_15_bF$buf44 ),
    .Y(_7558_)
);

OAI21X1 _18517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf27 ),
    .B(_7557_),
    .C(_7558_),
    .Y(_7559_)
);

NAND3X1 _18518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_bF$buf25 ),
    .B(_7559_),
    .C(_7556_),
    .Y(_7560_)
);

AOI21X1 _18519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7553_),
    .B(_7560_),
    .C(\datapath.idinstr_18_bF$buf6 ),
    .Y(_7561_)
);

OAI21X1 _18520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7546_),
    .B(_7561_),
    .C(_6140__bF$buf3),
    .Y(_7562_)
);

AOI21X1 _18521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7537_),
    .B(_7562_),
    .C(_6147__bF$buf4),
    .Y(\datapath.registers.rega_data [30])
);

MUX2X1 _18522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [31]),
    .B(\datapath.registers.1226[24] [31]),
    .S(\datapath.idinstr_15_bF$buf43 ),
    .Y(_7563_)
);

MUX2X1 _18523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [31]),
    .B(\datapath.registers.1226[26] [31]),
    .S(\datapath.idinstr_15_bF$buf42 ),
    .Y(_7564_)
);

MUX2X1 _18524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7564_),
    .B(_7563_),
    .S(\datapath.idinstr_16_bF$buf24 ),
    .Y(_7565_)
);

NAND2X1 _18525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf1),
    .B(_7565_),
    .Y(_7566_)
);

MUX2X1 _18526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [31]),
    .B(\datapath.registers.1226[28] [31]),
    .S(\datapath.idinstr_15_bF$buf41 ),
    .Y(_7567_)
);

MUX2X1 _18527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [31]),
    .B(\datapath.registers.1226[30] [31]),
    .S(\datapath.idinstr_15_bF$buf40 ),
    .Y(_7568_)
);

MUX2X1 _18528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7568_),
    .B(_7567_),
    .S(\datapath.idinstr_16_bF$buf23 ),
    .Y(_7569_)
);

NAND2X1 _18529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf26 ),
    .B(_7569_),
    .Y(_7570_)
);

AOI21X1 _18530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7566_),
    .B(_7570_),
    .C(_6145__bF$buf0),
    .Y(_7571_)
);

MUX2X1 _18531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [31]),
    .B(\datapath.registers.1226[16] [31]),
    .S(\datapath.idinstr_16_bF$buf22 ),
    .Y(_7572_)
);

NAND2X1 _18532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf9),
    .B(_7572_),
    .Y(_7573_)
);

MUX2X1 _18533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [31]),
    .B(\datapath.registers.1226[17] [31]),
    .S(\datapath.idinstr_16_bF$buf21 ),
    .Y(_7574_)
);

AOI21X1 _18534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf39 ),
    .B(_7574_),
    .C(\datapath.idinstr_17_bF$buf25 ),
    .Y(_7575_)
);

NAND2X1 _18535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7573_),
    .B(_7575_),
    .Y(_7576_)
);

MUX2X1 _18536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [31]),
    .B(\datapath.registers.1226[20] [31]),
    .S(\datapath.idinstr_16_bF$buf20 ),
    .Y(_7577_)
);

NAND2X1 _18537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141__bF$buf8),
    .B(_7577_),
    .Y(_7578_)
);

MUX2X1 _18538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [31]),
    .B(\datapath.registers.1226[21] [31]),
    .S(\datapath.idinstr_16_bF$buf19 ),
    .Y(_7579_)
);

AOI21X1 _18539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf38 ),
    .B(_7579_),
    .C(_6144__bF$buf0),
    .Y(_7580_)
);

NAND2X1 _18540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7578_),
    .B(_7580_),
    .Y(_7581_)
);

AOI21X1 _18541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7576_),
    .B(_7581_),
    .C(\datapath.idinstr_18_bF$buf5 ),
    .Y(_7582_)
);

OAI21X1 _18542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7571_),
    .B(_7582_),
    .C(\datapath.idinstr_19_bF$buf0 ),
    .Y(_7583_)
);

MUX2X1 _18543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [31]),
    .B(\datapath.registers.1226[8] [31]),
    .S(\datapath.idinstr_15_bF$buf37 ),
    .Y(_7584_)
);

MUX2X1 _18544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [31]),
    .B(\datapath.registers.1226[10] [31]),
    .S(\datapath.idinstr_15_bF$buf36 ),
    .Y(_7585_)
);

MUX2X1 _18545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7585_),
    .B(_7584_),
    .S(\datapath.idinstr_16_bF$buf18 ),
    .Y(_7586_)
);

NAND2X1 _18546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf10),
    .B(_7586_),
    .Y(_7587_)
);

INVX1 _18547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [31]),
    .Y(_7588_)
);

NOR2X1 _18548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7588_),
    .B(_6141__bF$buf7),
    .Y(_7589_)
);

INVX1 _18549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [31]),
    .Y(_7590_)
);

OAI21X1 _18550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7590_),
    .B(\datapath.idinstr_15_bF$buf35 ),
    .C(\datapath.idinstr_16_bF$buf17 ),
    .Y(_7591_)
);

NAND2X1 _18551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [31]),
    .B(_6141__bF$buf6),
    .Y(_7592_)
);

AOI21X1 _18552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [31]),
    .B(\datapath.idinstr_15_bF$buf34 ),
    .C(\datapath.idinstr_16_bF$buf16 ),
    .Y(_7593_)
);

AOI21X1 _18553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7593_),
    .B(_7592_),
    .C(_6144__bF$buf9),
    .Y(_7594_)
);

OAI21X1 _18554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7589_),
    .B(_7591_),
    .C(_7594_),
    .Y(_7595_)
);

AOI21X1 _18555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7595_),
    .B(_7587_),
    .C(_6145__bF$buf7),
    .Y(_7596_)
);

MUX2X1 _18556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [31]),
    .B(\datapath.registers.1226[4] [31]),
    .S(\datapath.idinstr_15_bF$buf33 ),
    .Y(_7597_)
);

MUX2X1 _18557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [31]),
    .B(\datapath.registers.1226[6] [31]),
    .S(\datapath.idinstr_15_bF$buf32 ),
    .Y(_7598_)
);

MUX2X1 _18558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7598_),
    .B(_7597_),
    .S(\datapath.idinstr_16_bF$buf15 ),
    .Y(_7599_)
);

NAND2X1 _18559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf24 ),
    .B(_7599_),
    .Y(_7600_)
);

MUX2X1 _18560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [31]),
    .B(\datapath.registers.1226[0] [31]),
    .S(\datapath.idinstr_15_bF$buf31 ),
    .Y(_7601_)
);

MUX2X1 _18561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [31]),
    .B(\datapath.registers.1226[2] [31]),
    .S(\datapath.idinstr_15_bF$buf30 ),
    .Y(_7602_)
);

MUX2X1 _18562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7602_),
    .B(_7601_),
    .S(\datapath.idinstr_16_bF$buf14 ),
    .Y(_7603_)
);

NAND2X1 _18563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144__bF$buf8),
    .B(_7603_),
    .Y(_7604_)
);

AOI21X1 _18564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7600_),
    .B(_7604_),
    .C(\datapath.idinstr_18_bF$buf4 ),
    .Y(_7605_)
);

OAI21X1 _18565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7605_),
    .B(_7596_),
    .C(_6140__bF$buf2),
    .Y(_7606_)
);

AOI21X1 _18566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7583_),
    .B(_7606_),
    .C(_6147__bF$buf3),
    .Y(\datapath.registers.rega_data [31])
);

INVX8 _18567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_24_bF$buf1 ),
    .Y(_7607_)
);

INVX8 _18568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf49 ),
    .Y(_7608_)
);

NAND2X1 _18569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7607__bF$buf4),
    .B(_7608__bF$buf10),
    .Y(_7609_)
);

INVX8 _18570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf38 ),
    .Y(_7610_)
);

INVX8 _18571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf37 ),
    .Y(_7611_)
);

INVX8 _18572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_23_bF$buf2 ),
    .Y(_7612_)
);

NAND3X1 _18573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf4),
    .B(_7611__bF$buf10),
    .C(_7612__bF$buf7),
    .Y(_7613_)
);

NOR2X1 _18574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7609_),
    .B(_7613_),
    .Y(_7614_)
);

MUX2X1 _18575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [0]),
    .B(\datapath.registers.1226[24] [0]),
    .S(\datapath.idinstr_20_bF$buf48 ),
    .Y(_7615_)
);

MUX2X1 _18576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [0]),
    .B(\datapath.registers.1226[26] [0]),
    .S(\datapath.idinstr_20_bF$buf47 ),
    .Y(_7616_)
);

MUX2X1 _18577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7616_),
    .B(_7615_),
    .S(\datapath.idinstr_21_bF$buf37 ),
    .Y(_7617_)
);

NAND2X1 _18578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf9),
    .B(_7617_),
    .Y(_7618_)
);

MUX2X1 _18579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [0]),
    .B(\datapath.registers.1226[28] [0]),
    .S(\datapath.idinstr_20_bF$buf46 ),
    .Y(_7619_)
);

MUX2X1 _18580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [0]),
    .B(\datapath.registers.1226[30] [0]),
    .S(\datapath.idinstr_20_bF$buf45 ),
    .Y(_7620_)
);

MUX2X1 _18581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7620_),
    .B(_7619_),
    .S(\datapath.idinstr_21_bF$buf36 ),
    .Y(_7621_)
);

NAND2X1 _18582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf36 ),
    .B(_7621_),
    .Y(_7622_)
);

AOI21X1 _18583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7618_),
    .B(_7622_),
    .C(_7612__bF$buf6),
    .Y(_7623_)
);

MUX2X1 _18584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [0]),
    .B(\datapath.registers.1226[16] [0]),
    .S(\datapath.idinstr_21_bF$buf35 ),
    .Y(_7624_)
);

NAND2X1 _18585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf9),
    .B(_7624_),
    .Y(_7625_)
);

MUX2X1 _18586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [0]),
    .B(\datapath.registers.1226[17] [0]),
    .S(\datapath.idinstr_21_bF$buf34 ),
    .Y(_7626_)
);

AOI21X1 _18587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf44 ),
    .B(_7626_),
    .C(\datapath.idinstr_22_bF$buf35 ),
    .Y(_7627_)
);

NAND2X1 _18588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7625_),
    .B(_7627_),
    .Y(_7628_)
);

MUX2X1 _18589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [0]),
    .B(\datapath.registers.1226[20] [0]),
    .S(\datapath.idinstr_21_bF$buf33 ),
    .Y(_7629_)
);

NAND2X1 _18590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf8),
    .B(_7629_),
    .Y(_7630_)
);

MUX2X1 _18591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [0]),
    .B(\datapath.registers.1226[21] [0]),
    .S(\datapath.idinstr_21_bF$buf32 ),
    .Y(_7631_)
);

AOI21X1 _18592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf43 ),
    .B(_7631_),
    .C(_7611__bF$buf8),
    .Y(_7632_)
);

NAND2X1 _18593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7630_),
    .B(_7632_),
    .Y(_7633_)
);

AOI21X1 _18594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7628_),
    .B(_7633_),
    .C(\datapath.idinstr_23_bF$buf1 ),
    .Y(_7634_)
);

OAI21X1 _18595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7623_),
    .B(_7634_),
    .C(\datapath.idinstr_24_bF$buf0 ),
    .Y(_7635_)
);

MUX2X1 _18596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [0]),
    .B(\datapath.registers.1226[8] [0]),
    .S(\datapath.idinstr_20_bF$buf42 ),
    .Y(_7636_)
);

MUX2X1 _18597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [0]),
    .B(\datapath.registers.1226[10] [0]),
    .S(\datapath.idinstr_20_bF$buf41 ),
    .Y(_7637_)
);

MUX2X1 _18598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7637_),
    .B(_7636_),
    .S(\datapath.idinstr_21_bF$buf31 ),
    .Y(_7638_)
);

NAND2X1 _18599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf7),
    .B(_7638_),
    .Y(_7639_)
);

MUX2X1 _18600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [0]),
    .B(\datapath.registers.1226[12] [0]),
    .S(\datapath.idinstr_20_bF$buf40 ),
    .Y(_7640_)
);

MUX2X1 _18601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [0]),
    .B(\datapath.registers.1226[14] [0]),
    .S(\datapath.idinstr_20_bF$buf39 ),
    .Y(_7641_)
);

MUX2X1 _18602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7641_),
    .B(_7640_),
    .S(\datapath.idinstr_21_bF$buf30 ),
    .Y(_7642_)
);

NAND2X1 _18603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf34 ),
    .B(_7642_),
    .Y(_7643_)
);

AOI21X1 _18604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7639_),
    .B(_7643_),
    .C(_7612__bF$buf5),
    .Y(_7644_)
);

AOI21X1 _18605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [0]),
    .B(\datapath.idinstr_22_bF$buf33 ),
    .C(_7608__bF$buf7),
    .Y(_7645_)
);

OAI21X1 _18606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6148_),
    .B(\datapath.idinstr_22_bF$buf32 ),
    .C(_7645_),
    .Y(_7646_)
);

AOI21X1 _18607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [0]),
    .B(\datapath.idinstr_22_bF$buf31 ),
    .C(\datapath.idinstr_20_bF$buf38 ),
    .Y(_7647_)
);

OAI21X1 _18608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6151_),
    .B(\datapath.idinstr_22_bF$buf30 ),
    .C(_7647_),
    .Y(_7648_)
);

NAND3X1 _18609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf3),
    .B(_7648_),
    .C(_7646_),
    .Y(_7649_)
);

AOI21X1 _18610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [0]),
    .B(\datapath.idinstr_22_bF$buf29 ),
    .C(_7608__bF$buf6),
    .Y(_7650_)
);

OAI21X1 _18611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6155_),
    .B(\datapath.idinstr_22_bF$buf28 ),
    .C(_7650_),
    .Y(_7651_)
);

AOI21X1 _18612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[6] [0]),
    .B(\datapath.idinstr_22_bF$buf27 ),
    .C(\datapath.idinstr_20_bF$buf37 ),
    .Y(_7652_)
);

OAI21X1 _18613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6158_),
    .B(\datapath.idinstr_22_bF$buf26 ),
    .C(_7652_),
    .Y(_7653_)
);

NAND3X1 _18614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf29 ),
    .B(_7653_),
    .C(_7651_),
    .Y(_7654_)
);

AOI21X1 _18615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7649_),
    .B(_7654_),
    .C(\datapath.idinstr_23_bF$buf0 ),
    .Y(_7655_)
);

OAI21X1 _18616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7644_),
    .B(_7655_),
    .C(_7607__bF$buf3),
    .Y(_7656_)
);

AOI21X1 _18617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7635_),
    .B(_7656_),
    .C(_7614__bF$buf4),
    .Y(\datapath.registers.regb_data [0])
);

MUX2X1 _18618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [1]),
    .B(\datapath.registers.1226[24] [1]),
    .S(\datapath.idinstr_20_bF$buf36 ),
    .Y(_7657_)
);

MUX2X1 _18619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [1]),
    .B(\datapath.registers.1226[26] [1]),
    .S(\datapath.idinstr_20_bF$buf35 ),
    .Y(_7658_)
);

MUX2X1 _18620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7658_),
    .B(_7657_),
    .S(\datapath.idinstr_21_bF$buf28 ),
    .Y(_7659_)
);

NAND2X1 _18621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf6),
    .B(_7659_),
    .Y(_7660_)
);

MUX2X1 _18622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [1]),
    .B(\datapath.registers.1226[28] [1]),
    .S(\datapath.idinstr_20_bF$buf34 ),
    .Y(_7661_)
);

MUX2X1 _18623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [1]),
    .B(\datapath.registers.1226[30] [1]),
    .S(\datapath.idinstr_20_bF$buf33 ),
    .Y(_7662_)
);

MUX2X1 _18624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7662_),
    .B(_7661_),
    .S(\datapath.idinstr_21_bF$buf27 ),
    .Y(_7663_)
);

NAND2X1 _18625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf25 ),
    .B(_7663_),
    .Y(_7664_)
);

AOI21X1 _18626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7660_),
    .B(_7664_),
    .C(_7612__bF$buf4),
    .Y(_7665_)
);

MUX2X1 _18627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [1]),
    .B(\datapath.registers.1226[16] [1]),
    .S(\datapath.idinstr_21_bF$buf26 ),
    .Y(_7666_)
);

NAND2X1 _18628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf5),
    .B(_7666_),
    .Y(_7667_)
);

MUX2X1 _18629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [1]),
    .B(\datapath.registers.1226[17] [1]),
    .S(\datapath.idinstr_21_bF$buf25 ),
    .Y(_7668_)
);

AOI21X1 _18630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf32 ),
    .B(_7668_),
    .C(\datapath.idinstr_22_bF$buf24 ),
    .Y(_7669_)
);

NAND2X1 _18631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7667_),
    .B(_7669_),
    .Y(_7670_)
);

MUX2X1 _18632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [1]),
    .B(\datapath.registers.1226[20] [1]),
    .S(\datapath.idinstr_21_bF$buf24 ),
    .Y(_7671_)
);

NAND2X1 _18633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf4),
    .B(_7671_),
    .Y(_7672_)
);

MUX2X1 _18634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [1]),
    .B(\datapath.registers.1226[21] [1]),
    .S(\datapath.idinstr_21_bF$buf23 ),
    .Y(_7673_)
);

AOI21X1 _18635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf31 ),
    .B(_7673_),
    .C(_7611__bF$buf5),
    .Y(_7674_)
);

NAND2X1 _18636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7672_),
    .B(_7674_),
    .Y(_7675_)
);

AOI21X1 _18637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7670_),
    .B(_7675_),
    .C(\datapath.idinstr_23_bF$buf7 ),
    .Y(_7676_)
);

OAI21X1 _18638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7665_),
    .B(_7676_),
    .C(\datapath.idinstr_24_bF$buf5 ),
    .Y(_7677_)
);

MUX2X1 _18639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [1]),
    .B(\datapath.registers.1226[8] [1]),
    .S(\datapath.idinstr_20_bF$buf30 ),
    .Y(_7678_)
);

MUX2X1 _18640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [1]),
    .B(\datapath.registers.1226[10] [1]),
    .S(\datapath.idinstr_20_bF$buf29 ),
    .Y(_7679_)
);

MUX2X1 _18641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7679_),
    .B(_7678_),
    .S(\datapath.idinstr_21_bF$buf22 ),
    .Y(_7680_)
);

NAND2X1 _18642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf4),
    .B(_7680_),
    .Y(_7681_)
);

MUX2X1 _18643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [1]),
    .B(\datapath.registers.1226[12] [1]),
    .S(\datapath.idinstr_20_bF$buf28 ),
    .Y(_7682_)
);

MUX2X1 _18644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [1]),
    .B(\datapath.registers.1226[14] [1]),
    .S(\datapath.idinstr_20_bF$buf27 ),
    .Y(_7683_)
);

MUX2X1 _18645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7683_),
    .B(_7682_),
    .S(\datapath.idinstr_21_bF$buf21 ),
    .Y(_7684_)
);

NAND2X1 _18646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf23 ),
    .B(_7684_),
    .Y(_7685_)
);

AOI21X1 _18647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7681_),
    .B(_7685_),
    .C(_7612__bF$buf3),
    .Y(_7686_)
);

AOI21X1 _18648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [1]),
    .B(\datapath.idinstr_22_bF$buf22 ),
    .C(_7608__bF$buf3),
    .Y(_7687_)
);

OAI21X1 _18649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6206_),
    .B(\datapath.idinstr_22_bF$buf21 ),
    .C(_7687_),
    .Y(_7688_)
);

INVX1 _18650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [1]),
    .Y(_7689_)
);

AOI21X1 _18651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [1]),
    .B(\datapath.idinstr_22_bF$buf20 ),
    .C(\datapath.idinstr_20_bF$buf26 ),
    .Y(_7690_)
);

OAI21X1 _18652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7689_),
    .B(\datapath.idinstr_22_bF$buf19 ),
    .C(_7690_),
    .Y(_7691_)
);

NAND3X1 _18653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf2),
    .B(_7691_),
    .C(_7688_),
    .Y(_7692_)
);

AOI21X1 _18654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [1]),
    .B(\datapath.idinstr_22_bF$buf18 ),
    .C(_7608__bF$buf2),
    .Y(_7693_)
);

OAI21X1 _18655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6213_),
    .B(\datapath.idinstr_22_bF$buf17 ),
    .C(_7693_),
    .Y(_7694_)
);

AOI21X1 _18656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[6] [1]),
    .B(\datapath.idinstr_22_bF$buf16 ),
    .C(\datapath.idinstr_20_bF$buf25 ),
    .Y(_7695_)
);

OAI21X1 _18657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6216_),
    .B(\datapath.idinstr_22_bF$buf15 ),
    .C(_7695_),
    .Y(_7696_)
);

NAND3X1 _18658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf20 ),
    .B(_7696_),
    .C(_7694_),
    .Y(_7697_)
);

AOI21X1 _18659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7692_),
    .B(_7697_),
    .C(\datapath.idinstr_23_bF$buf6 ),
    .Y(_7698_)
);

OAI21X1 _18660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7686_),
    .B(_7698_),
    .C(_7607__bF$buf2),
    .Y(_7699_)
);

AOI21X1 _18661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7677_),
    .B(_7699_),
    .C(_7614__bF$buf3),
    .Y(\datapath.registers.regb_data [1])
);

MUX2X1 _18662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [2]),
    .B(\datapath.registers.1226[24] [2]),
    .S(\datapath.idinstr_20_bF$buf24 ),
    .Y(_7700_)
);

MUX2X1 _18663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [2]),
    .B(\datapath.registers.1226[26] [2]),
    .S(\datapath.idinstr_20_bF$buf23 ),
    .Y(_7701_)
);

MUX2X1 _18664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7701_),
    .B(_7700_),
    .S(\datapath.idinstr_21_bF$buf19 ),
    .Y(_7702_)
);

NAND2X1 _18665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf3),
    .B(_7702_),
    .Y(_7703_)
);

MUX2X1 _18666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [2]),
    .B(\datapath.registers.1226[28] [2]),
    .S(\datapath.idinstr_20_bF$buf22 ),
    .Y(_7704_)
);

MUX2X1 _18667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [2]),
    .B(\datapath.registers.1226[30] [2]),
    .S(\datapath.idinstr_20_bF$buf21 ),
    .Y(_7705_)
);

MUX2X1 _18668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7705_),
    .B(_7704_),
    .S(\datapath.idinstr_21_bF$buf18 ),
    .Y(_7706_)
);

NAND2X1 _18669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf14 ),
    .B(_7706_),
    .Y(_7707_)
);

AOI21X1 _18670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7703_),
    .B(_7707_),
    .C(_7612__bF$buf2),
    .Y(_7708_)
);

MUX2X1 _18671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [2]),
    .B(\datapath.registers.1226[16] [2]),
    .S(\datapath.idinstr_21_bF$buf17 ),
    .Y(_7709_)
);

NAND2X1 _18672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf1),
    .B(_7709_),
    .Y(_7710_)
);

MUX2X1 _18673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [2]),
    .B(\datapath.registers.1226[17] [2]),
    .S(\datapath.idinstr_21_bF$buf16 ),
    .Y(_7711_)
);

AOI21X1 _18674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf20 ),
    .B(_7711_),
    .C(\datapath.idinstr_22_bF$buf13 ),
    .Y(_7712_)
);

NAND2X1 _18675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7710_),
    .B(_7712_),
    .Y(_7713_)
);

MUX2X1 _18676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [2]),
    .B(\datapath.registers.1226[20] [2]),
    .S(\datapath.idinstr_21_bF$buf15 ),
    .Y(_7714_)
);

NAND2X1 _18677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf0),
    .B(_7714_),
    .Y(_7715_)
);

MUX2X1 _18678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [2]),
    .B(\datapath.registers.1226[21] [2]),
    .S(\datapath.idinstr_21_bF$buf14 ),
    .Y(_7716_)
);

AOI21X1 _18679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf19 ),
    .B(_7716_),
    .C(_7611__bF$buf2),
    .Y(_7717_)
);

NAND2X1 _18680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7715_),
    .B(_7717_),
    .Y(_7718_)
);

AOI21X1 _18681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7713_),
    .B(_7718_),
    .C(\datapath.idinstr_23_bF$buf5 ),
    .Y(_7719_)
);

OAI21X1 _18682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7708_),
    .B(_7719_),
    .C(\datapath.idinstr_24_bF$buf4 ),
    .Y(_7720_)
);

MUX2X1 _18683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [2]),
    .B(\datapath.registers.1226[8] [2]),
    .S(\datapath.idinstr_20_bF$buf18 ),
    .Y(_7721_)
);

MUX2X1 _18684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [2]),
    .B(\datapath.registers.1226[10] [2]),
    .S(\datapath.idinstr_20_bF$buf17 ),
    .Y(_7722_)
);

MUX2X1 _18685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7722_),
    .B(_7721_),
    .S(\datapath.idinstr_21_bF$buf13 ),
    .Y(_7723_)
);

NAND2X1 _18686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf1),
    .B(_7723_),
    .Y(_7724_)
);

AND2X2 _18687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [2]),
    .B(\datapath.idinstr_20_bF$buf16 ),
    .Y(_7725_)
);

INVX1 _18688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [2]),
    .Y(_7726_)
);

OAI21X1 _18689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7726_),
    .B(\datapath.idinstr_20_bF$buf15 ),
    .C(\datapath.idinstr_21_bF$buf12 ),
    .Y(_7727_)
);

NAND2X1 _18690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [2]),
    .B(_7608__bF$buf10),
    .Y(_7728_)
);

AOI21X1 _18691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [2]),
    .B(\datapath.idinstr_20_bF$buf14 ),
    .C(\datapath.idinstr_21_bF$buf11 ),
    .Y(_7729_)
);

AOI21X1 _18692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7729_),
    .B(_7728_),
    .C(_7611__bF$buf0),
    .Y(_7730_)
);

OAI21X1 _18693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7725_),
    .B(_7727_),
    .C(_7730_),
    .Y(_7731_)
);

AOI21X1 _18694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7731_),
    .B(_7724_),
    .C(_7612__bF$buf1),
    .Y(_7732_)
);

MUX2X1 _18695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [2]),
    .B(\datapath.registers.1226[4] [2]),
    .S(\datapath.idinstr_20_bF$buf13 ),
    .Y(_7733_)
);

MUX2X1 _18696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [2]),
    .B(\datapath.registers.1226[6] [2]),
    .S(\datapath.idinstr_20_bF$buf12 ),
    .Y(_7734_)
);

MUX2X1 _18697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7734_),
    .B(_7733_),
    .S(\datapath.idinstr_21_bF$buf10 ),
    .Y(_7735_)
);

NAND2X1 _18698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf12 ),
    .B(_7735_),
    .Y(_7736_)
);

MUX2X1 _18699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [2]),
    .B(\datapath.registers.1226[0] [2]),
    .S(\datapath.idinstr_20_bF$buf11 ),
    .Y(_7737_)
);

MUX2X1 _18700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [2]),
    .B(\datapath.registers.1226[2] [2]),
    .S(\datapath.idinstr_20_bF$buf10 ),
    .Y(_7738_)
);

MUX2X1 _18701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7738_),
    .B(_7737_),
    .S(\datapath.idinstr_21_bF$buf9 ),
    .Y(_7739_)
);

NAND2X1 _18702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf10),
    .B(_7739_),
    .Y(_7740_)
);

AOI21X1 _18703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7736_),
    .B(_7740_),
    .C(\datapath.idinstr_23_bF$buf4 ),
    .Y(_7741_)
);

OAI21X1 _18704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7741_),
    .B(_7732_),
    .C(_7607__bF$buf1),
    .Y(_7742_)
);

AOI21X1 _18705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7720_),
    .B(_7742_),
    .C(_7614__bF$buf2),
    .Y(\datapath.registers.regb_data [2])
);

MUX2X1 _18706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [3]),
    .B(\datapath.registers.1226[0] [3]),
    .S(\datapath.idinstr_20_bF$buf9 ),
    .Y(_7743_)
);

MUX2X1 _18707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [3]),
    .B(\datapath.registers.1226[2] [3]),
    .S(\datapath.idinstr_20_bF$buf8 ),
    .Y(_7744_)
);

MUX2X1 _18708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7744_),
    .B(_7743_),
    .S(\datapath.idinstr_21_bF$buf8 ),
    .Y(_7745_)
);

NAND2X1 _18709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf9),
    .B(_7745_),
    .Y(_7746_)
);

MUX2X1 _18710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [3]),
    .B(\datapath.registers.1226[4] [3]),
    .S(\datapath.idinstr_20_bF$buf7 ),
    .Y(_7747_)
);

MUX2X1 _18711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [3]),
    .B(\datapath.registers.1226[6] [3]),
    .S(\datapath.idinstr_20_bF$buf6 ),
    .Y(_7748_)
);

MUX2X1 _18712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7748_),
    .B(_7747_),
    .S(\datapath.idinstr_21_bF$buf7 ),
    .Y(_7749_)
);

NAND2X1 _18713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf11 ),
    .B(_7749_),
    .Y(_7750_)
);

AOI21X1 _18714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7746_),
    .B(_7750_),
    .C(\datapath.idinstr_23_bF$buf3 ),
    .Y(_7751_)
);

INVX1 _18715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [3]),
    .Y(_7752_)
);

AOI21X1 _18716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [3]),
    .B(\datapath.idinstr_22_bF$buf10 ),
    .C(_7608__bF$buf9),
    .Y(_7753_)
);

OAI21X1 _18717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7752_),
    .B(\datapath.idinstr_22_bF$buf9 ),
    .C(_7753_),
    .Y(_7754_)
);

NAND2X1 _18718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [3]),
    .B(_7611__bF$buf8),
    .Y(_7755_)
);

AOI21X1 _18719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [3]),
    .B(\datapath.idinstr_22_bF$buf8 ),
    .C(\datapath.idinstr_20_bF$buf5 ),
    .Y(_7756_)
);

AOI21X1 _18720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7756_),
    .B(_7755_),
    .C(\datapath.idinstr_21_bF$buf6 ),
    .Y(_7757_)
);

NAND2X1 _18721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7754_),
    .B(_7757_),
    .Y(_7758_)
);

INVX1 _18722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [3]),
    .Y(_7759_)
);

AOI21X1 _18723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [3]),
    .B(\datapath.idinstr_22_bF$buf7 ),
    .C(_7608__bF$buf8),
    .Y(_7760_)
);

OAI21X1 _18724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7759_),
    .B(\datapath.idinstr_22_bF$buf6 ),
    .C(_7760_),
    .Y(_7761_)
);

INVX1 _18725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[10] [3]),
    .Y(_7762_)
);

AOI21X1 _18726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [3]),
    .B(\datapath.idinstr_22_bF$buf5 ),
    .C(\datapath.idinstr_20_bF$buf4 ),
    .Y(_7763_)
);

OAI21X1 _18727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7762_),
    .B(\datapath.idinstr_22_bF$buf4 ),
    .C(_7763_),
    .Y(_7764_)
);

NAND3X1 _18728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf5 ),
    .B(_7764_),
    .C(_7761_),
    .Y(_7765_)
);

AOI21X1 _18729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7758_),
    .B(_7765_),
    .C(_7612__bF$buf0),
    .Y(_7766_)
);

OAI21X1 _18730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7751_),
    .B(_7766_),
    .C(_7607__bF$buf0),
    .Y(_7767_)
);

MUX2X1 _18731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [3]),
    .B(\datapath.registers.1226[16] [3]),
    .S(\datapath.idinstr_20_bF$buf3 ),
    .Y(_7768_)
);

MUX2X1 _18732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [3]),
    .B(\datapath.registers.1226[18] [3]),
    .S(\datapath.idinstr_20_bF$buf2 ),
    .Y(_7769_)
);

MUX2X1 _18733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7769_),
    .B(_7768_),
    .S(\datapath.idinstr_21_bF$buf4 ),
    .Y(_7770_)
);

NAND2X1 _18734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf7),
    .B(_7770_),
    .Y(_7771_)
);

MUX2X1 _18735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [3]),
    .B(\datapath.registers.1226[20] [3]),
    .S(\datapath.idinstr_20_bF$buf1 ),
    .Y(_7772_)
);

MUX2X1 _18736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [3]),
    .B(\datapath.registers.1226[22] [3]),
    .S(\datapath.idinstr_20_bF$buf0 ),
    .Y(_7773_)
);

MUX2X1 _18737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7773_),
    .B(_7772_),
    .S(\datapath.idinstr_21_bF$buf3 ),
    .Y(_7774_)
);

NAND2X1 _18738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf3 ),
    .B(_7774_),
    .Y(_7775_)
);

AOI21X1 _18739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7771_),
    .B(_7775_),
    .C(\datapath.idinstr_23_bF$buf2 ),
    .Y(_7776_)
);

INVX1 _18740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [3]),
    .Y(_7777_)
);

AOI21X1 _18741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [3]),
    .B(\datapath.idinstr_22_bF$buf2 ),
    .C(_7608__bF$buf7),
    .Y(_7778_)
);

OAI21X1 _18742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7777_),
    .B(\datapath.idinstr_22_bF$buf1 ),
    .C(_7778_),
    .Y(_7779_)
);

INVX1 _18743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [3]),
    .Y(_7780_)
);

AOI21X1 _18744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [3]),
    .B(\datapath.idinstr_22_bF$buf0 ),
    .C(\datapath.idinstr_20_bF$buf55 ),
    .Y(_7781_)
);

OAI21X1 _18745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7780_),
    .B(\datapath.idinstr_22_bF$buf43 ),
    .C(_7781_),
    .Y(_7782_)
);

NAND3X1 _18746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf2 ),
    .B(_7782_),
    .C(_7779_),
    .Y(_7783_)
);

INVX1 _18747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [3]),
    .Y(_7784_)
);

AOI21X1 _18748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [3]),
    .B(\datapath.idinstr_22_bF$buf42 ),
    .C(_7608__bF$buf6),
    .Y(_7785_)
);

OAI21X1 _18749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7784_),
    .B(\datapath.idinstr_22_bF$buf41 ),
    .C(_7785_),
    .Y(_7786_)
);

AOI21X1 _18750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[28] [3]),
    .B(\datapath.idinstr_22_bF$buf40 ),
    .C(\datapath.idinstr_20_bF$buf54 ),
    .Y(_7787_)
);

OAI21X1 _18751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5719_),
    .B(\datapath.idinstr_22_bF$buf39 ),
    .C(_7787_),
    .Y(_7788_)
);

NAND3X1 _18752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf1),
    .B(_7788_),
    .C(_7786_),
    .Y(_7789_)
);

AOI21X1 _18753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7783_),
    .B(_7789_),
    .C(_7612__bF$buf7),
    .Y(_7790_)
);

OAI21X1 _18754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7776_),
    .B(_7790_),
    .C(\datapath.idinstr_24_bF$buf3 ),
    .Y(_7791_)
);

AOI21X1 _18755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7767_),
    .B(_7791_),
    .C(_7614__bF$buf1),
    .Y(\datapath.registers.regb_data [3])
);

MUX2X1 _18756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [4]),
    .B(\datapath.registers.1226[24] [4]),
    .S(\datapath.idinstr_20_bF$buf53 ),
    .Y(_7792_)
);

MUX2X1 _18757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [4]),
    .B(\datapath.registers.1226[26] [4]),
    .S(\datapath.idinstr_20_bF$buf52 ),
    .Y(_7793_)
);

MUX2X1 _18758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7793_),
    .B(_7792_),
    .S(\datapath.idinstr_21_bF$buf1 ),
    .Y(_7794_)
);

NAND2X1 _18759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf6),
    .B(_7794_),
    .Y(_7795_)
);

MUX2X1 _18760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [4]),
    .B(\datapath.registers.1226[28] [4]),
    .S(\datapath.idinstr_20_bF$buf51 ),
    .Y(_7796_)
);

MUX2X1 _18761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [4]),
    .B(\datapath.registers.1226[30] [4]),
    .S(\datapath.idinstr_20_bF$buf50 ),
    .Y(_7797_)
);

MUX2X1 _18762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7797_),
    .B(_7796_),
    .S(\datapath.idinstr_21_bF$buf0 ),
    .Y(_7798_)
);

NAND2X1 _18763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf38 ),
    .B(_7798_),
    .Y(_7799_)
);

AOI21X1 _18764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7795_),
    .B(_7799_),
    .C(_7612__bF$buf6),
    .Y(_7800_)
);

MUX2X1 _18765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [4]),
    .B(\datapath.registers.1226[16] [4]),
    .S(\datapath.idinstr_21_bF$buf44 ),
    .Y(_7801_)
);

NAND2X1 _18766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf5),
    .B(_7801_),
    .Y(_7802_)
);

MUX2X1 _18767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [4]),
    .B(\datapath.registers.1226[17] [4]),
    .S(\datapath.idinstr_21_bF$buf43 ),
    .Y(_7803_)
);

AOI21X1 _18768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf49 ),
    .B(_7803_),
    .C(\datapath.idinstr_22_bF$buf37 ),
    .Y(_7804_)
);

NAND2X1 _18769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7802_),
    .B(_7804_),
    .Y(_7805_)
);

MUX2X1 _18770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [4]),
    .B(\datapath.registers.1226[20] [4]),
    .S(\datapath.idinstr_21_bF$buf42 ),
    .Y(_7806_)
);

NAND2X1 _18771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf4),
    .B(_7806_),
    .Y(_7807_)
);

MUX2X1 _18772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [4]),
    .B(\datapath.registers.1226[21] [4]),
    .S(\datapath.idinstr_21_bF$buf41 ),
    .Y(_7808_)
);

AOI21X1 _18773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf48 ),
    .B(_7808_),
    .C(_7611__bF$buf5),
    .Y(_7809_)
);

NAND2X1 _18774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7807_),
    .B(_7809_),
    .Y(_7810_)
);

AOI21X1 _18775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7805_),
    .B(_7810_),
    .C(\datapath.idinstr_23_bF$buf1 ),
    .Y(_7811_)
);

OAI21X1 _18776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7800_),
    .B(_7811_),
    .C(\datapath.idinstr_24_bF$buf2 ),
    .Y(_7812_)
);

MUX2X1 _18777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [4]),
    .B(\datapath.registers.1226[8] [4]),
    .S(\datapath.idinstr_20_bF$buf47 ),
    .Y(_7813_)
);

MUX2X1 _18778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [4]),
    .B(\datapath.registers.1226[10] [4]),
    .S(\datapath.idinstr_20_bF$buf46 ),
    .Y(_7814_)
);

MUX2X1 _18779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7814_),
    .B(_7813_),
    .S(\datapath.idinstr_21_bF$buf40 ),
    .Y(_7815_)
);

NAND2X1 _18780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf4),
    .B(_7815_),
    .Y(_7816_)
);

NOR2X1 _18781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6363_),
    .B(_7608__bF$buf3),
    .Y(_7817_)
);

OAI21X1 _18782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6365_),
    .B(\datapath.idinstr_20_bF$buf45 ),
    .C(\datapath.idinstr_21_bF$buf39 ),
    .Y(_7818_)
);

NAND2X1 _18783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [4]),
    .B(_7608__bF$buf2),
    .Y(_7819_)
);

AOI21X1 _18784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [4]),
    .B(\datapath.idinstr_20_bF$buf44 ),
    .C(\datapath.idinstr_21_bF$buf38 ),
    .Y(_7820_)
);

AOI21X1 _18785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7820_),
    .B(_7819_),
    .C(_7611__bF$buf3),
    .Y(_7821_)
);

OAI21X1 _18786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7817_),
    .B(_7818_),
    .C(_7821_),
    .Y(_7822_)
);

AOI21X1 _18787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7822_),
    .B(_7816_),
    .C(_7612__bF$buf5),
    .Y(_7823_)
);

MUX2X1 _18788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [4]),
    .B(\datapath.registers.1226[4] [4]),
    .S(\datapath.idinstr_20_bF$buf43 ),
    .Y(_7824_)
);

MUX2X1 _18789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [4]),
    .B(\datapath.registers.1226[6] [4]),
    .S(\datapath.idinstr_20_bF$buf42 ),
    .Y(_7825_)
);

MUX2X1 _18790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7825_),
    .B(_7824_),
    .S(\datapath.idinstr_21_bF$buf37 ),
    .Y(_7826_)
);

NAND2X1 _18791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf36 ),
    .B(_7826_),
    .Y(_7827_)
);

MUX2X1 _18792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [4]),
    .B(\datapath.registers.1226[0] [4]),
    .S(\datapath.idinstr_20_bF$buf41 ),
    .Y(_7828_)
);

MUX2X1 _18793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [4]),
    .B(\datapath.registers.1226[2] [4]),
    .S(\datapath.idinstr_20_bF$buf40 ),
    .Y(_7829_)
);

MUX2X1 _18794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7829_),
    .B(_7828_),
    .S(\datapath.idinstr_21_bF$buf36 ),
    .Y(_7830_)
);

NAND2X1 _18795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf2),
    .B(_7830_),
    .Y(_7831_)
);

AOI21X1 _18796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7827_),
    .B(_7831_),
    .C(\datapath.idinstr_23_bF$buf0 ),
    .Y(_7832_)
);

OAI21X1 _18797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7832_),
    .B(_7823_),
    .C(_7607__bF$buf4),
    .Y(_7833_)
);

AOI21X1 _18798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7812_),
    .B(_7833_),
    .C(_7614__bF$buf0),
    .Y(\datapath.registers.regb_data [4])
);

MUX2X1 _18799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [5]),
    .B(\datapath.registers.1226[24] [5]),
    .S(\datapath.idinstr_20_bF$buf39 ),
    .Y(_7834_)
);

MUX2X1 _18800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [5]),
    .B(\datapath.registers.1226[26] [5]),
    .S(\datapath.idinstr_20_bF$buf38 ),
    .Y(_7835_)
);

MUX2X1 _18801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7835_),
    .B(_7834_),
    .S(\datapath.idinstr_21_bF$buf35 ),
    .Y(_7836_)
);

NAND2X1 _18802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf1),
    .B(_7836_),
    .Y(_7837_)
);

MUX2X1 _18803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [5]),
    .B(\datapath.registers.1226[28] [5]),
    .S(\datapath.idinstr_20_bF$buf37 ),
    .Y(_7838_)
);

MUX2X1 _18804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [5]),
    .B(\datapath.registers.1226[30] [5]),
    .S(\datapath.idinstr_20_bF$buf36 ),
    .Y(_7839_)
);

MUX2X1 _18805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7839_),
    .B(_7838_),
    .S(\datapath.idinstr_21_bF$buf34 ),
    .Y(_7840_)
);

NAND2X1 _18806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf35 ),
    .B(_7840_),
    .Y(_7841_)
);

AOI21X1 _18807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7837_),
    .B(_7841_),
    .C(_7612__bF$buf4),
    .Y(_7842_)
);

MUX2X1 _18808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [5]),
    .B(\datapath.registers.1226[16] [5]),
    .S(\datapath.idinstr_21_bF$buf33 ),
    .Y(_7843_)
);

NAND2X1 _18809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf1),
    .B(_7843_),
    .Y(_7844_)
);

MUX2X1 _18810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [5]),
    .B(\datapath.registers.1226[17] [5]),
    .S(\datapath.idinstr_21_bF$buf32 ),
    .Y(_7845_)
);

AOI21X1 _18811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf35 ),
    .B(_7845_),
    .C(\datapath.idinstr_22_bF$buf34 ),
    .Y(_7846_)
);

NAND2X1 _18812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7844_),
    .B(_7846_),
    .Y(_7847_)
);

MUX2X1 _18813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [5]),
    .B(\datapath.registers.1226[20] [5]),
    .S(\datapath.idinstr_21_bF$buf31 ),
    .Y(_7848_)
);

NAND2X1 _18814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf0),
    .B(_7848_),
    .Y(_7849_)
);

MUX2X1 _18815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [5]),
    .B(\datapath.registers.1226[21] [5]),
    .S(\datapath.idinstr_21_bF$buf30 ),
    .Y(_7850_)
);

AOI21X1 _18816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf34 ),
    .B(_7850_),
    .C(_7611__bF$buf0),
    .Y(_7851_)
);

NAND2X1 _18817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7849_),
    .B(_7851_),
    .Y(_7852_)
);

AOI21X1 _18818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7847_),
    .B(_7852_),
    .C(\datapath.idinstr_23_bF$buf7 ),
    .Y(_7853_)
);

OAI21X1 _18819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7842_),
    .B(_7853_),
    .C(\datapath.idinstr_24_bF$buf1 ),
    .Y(_7854_)
);

MUX2X1 _18820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [5]),
    .B(\datapath.registers.1226[8] [5]),
    .S(\datapath.idinstr_20_bF$buf33 ),
    .Y(_7855_)
);

MUX2X1 _18821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [5]),
    .B(\datapath.registers.1226[10] [5]),
    .S(\datapath.idinstr_20_bF$buf32 ),
    .Y(_7856_)
);

MUX2X1 _18822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7856_),
    .B(_7855_),
    .S(\datapath.idinstr_21_bF$buf29 ),
    .Y(_7857_)
);

NAND2X1 _18823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf10),
    .B(_7857_),
    .Y(_7858_)
);

AND2X2 _18824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [5]),
    .B(\datapath.idinstr_20_bF$buf31 ),
    .Y(_7859_)
);

INVX1 _18825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [5]),
    .Y(_7860_)
);

OAI21X1 _18826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7860_),
    .B(\datapath.idinstr_20_bF$buf30 ),
    .C(\datapath.idinstr_21_bF$buf28 ),
    .Y(_7861_)
);

NAND2X1 _18827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [5]),
    .B(_7608__bF$buf10),
    .Y(_7862_)
);

AOI21X1 _18828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [5]),
    .B(\datapath.idinstr_20_bF$buf29 ),
    .C(\datapath.idinstr_21_bF$buf27 ),
    .Y(_7863_)
);

AOI21X1 _18829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7863_),
    .B(_7862_),
    .C(_7611__bF$buf9),
    .Y(_7864_)
);

OAI21X1 _18830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7859_),
    .B(_7861_),
    .C(_7864_),
    .Y(_7865_)
);

AOI21X1 _18831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7865_),
    .B(_7858_),
    .C(_7612__bF$buf3),
    .Y(_7866_)
);

MUX2X1 _18832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [5]),
    .B(\datapath.registers.1226[4] [5]),
    .S(\datapath.idinstr_20_bF$buf28 ),
    .Y(_7867_)
);

MUX2X1 _18833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [5]),
    .B(\datapath.registers.1226[6] [5]),
    .S(\datapath.idinstr_20_bF$buf27 ),
    .Y(_7868_)
);

MUX2X1 _18834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7868_),
    .B(_7867_),
    .S(\datapath.idinstr_21_bF$buf26 ),
    .Y(_7869_)
);

NAND2X1 _18835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf33 ),
    .B(_7869_),
    .Y(_7870_)
);

MUX2X1 _18836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [5]),
    .B(\datapath.registers.1226[0] [5]),
    .S(\datapath.idinstr_20_bF$buf26 ),
    .Y(_7871_)
);

MUX2X1 _18837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [5]),
    .B(\datapath.registers.1226[2] [5]),
    .S(\datapath.idinstr_20_bF$buf25 ),
    .Y(_7872_)
);

MUX2X1 _18838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7872_),
    .B(_7871_),
    .S(\datapath.idinstr_21_bF$buf25 ),
    .Y(_7873_)
);

NAND2X1 _18839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf8),
    .B(_7873_),
    .Y(_7874_)
);

AOI21X1 _18840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7870_),
    .B(_7874_),
    .C(\datapath.idinstr_23_bF$buf6 ),
    .Y(_7875_)
);

OAI21X1 _18841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7875_),
    .B(_7866_),
    .C(_7607__bF$buf3),
    .Y(_7876_)
);

AOI21X1 _18842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7854_),
    .B(_7876_),
    .C(_7614__bF$buf4),
    .Y(\datapath.registers.regb_data [5])
);

MUX2X1 _18843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [6]),
    .B(\datapath.registers.1226[8] [6]),
    .S(\datapath.idinstr_20_bF$buf24 ),
    .Y(_7877_)
);

MUX2X1 _18844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [6]),
    .B(\datapath.registers.1226[10] [6]),
    .S(\datapath.idinstr_20_bF$buf23 ),
    .Y(_7878_)
);

MUX2X1 _18845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7878_),
    .B(_7877_),
    .S(\datapath.idinstr_21_bF$buf24 ),
    .Y(_7879_)
);

NAND2X1 _18846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf7),
    .B(_7879_),
    .Y(_7880_)
);

MUX2X1 _18847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [6]),
    .B(\datapath.registers.1226[12] [6]),
    .S(\datapath.idinstr_20_bF$buf22 ),
    .Y(_7881_)
);

MUX2X1 _18848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [6]),
    .B(\datapath.registers.1226[14] [6]),
    .S(\datapath.idinstr_20_bF$buf21 ),
    .Y(_7882_)
);

MUX2X1 _18849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7882_),
    .B(_7881_),
    .S(\datapath.idinstr_21_bF$buf23 ),
    .Y(_7883_)
);

NAND2X1 _18850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf32 ),
    .B(_7883_),
    .Y(_7884_)
);

AOI21X1 _18851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7880_),
    .B(_7884_),
    .C(_7612__bF$buf2),
    .Y(_7885_)
);

INVX1 _18852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [6]),
    .Y(_7886_)
);

AOI21X1 _18853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [6]),
    .B(\datapath.idinstr_22_bF$buf31 ),
    .C(_7608__bF$buf9),
    .Y(_7887_)
);

OAI21X1 _18854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7886_),
    .B(\datapath.idinstr_22_bF$buf30 ),
    .C(_7887_),
    .Y(_7888_)
);

NAND2X1 _18855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [6]),
    .B(_7611__bF$buf6),
    .Y(_7889_)
);

AOI21X1 _18856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [6]),
    .B(\datapath.idinstr_22_bF$buf29 ),
    .C(\datapath.idinstr_20_bF$buf20 ),
    .Y(_7890_)
);

AOI21X1 _18857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7890_),
    .B(_7889_),
    .C(\datapath.idinstr_21_bF$buf22 ),
    .Y(_7891_)
);

NAND2X1 _18858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7888_),
    .B(_7891_),
    .Y(_7892_)
);

INVX1 _18859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [6]),
    .Y(_7893_)
);

AOI21X1 _18860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [6]),
    .B(\datapath.idinstr_22_bF$buf28 ),
    .C(_7608__bF$buf8),
    .Y(_7894_)
);

OAI21X1 _18861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7893_),
    .B(\datapath.idinstr_22_bF$buf27 ),
    .C(_7894_),
    .Y(_7895_)
);

INVX1 _18862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[2] [6]),
    .Y(_7896_)
);

AOI21X1 _18863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[6] [6]),
    .B(\datapath.idinstr_22_bF$buf26 ),
    .C(\datapath.idinstr_20_bF$buf19 ),
    .Y(_7897_)
);

OAI21X1 _18864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7896_),
    .B(\datapath.idinstr_22_bF$buf25 ),
    .C(_7897_),
    .Y(_7898_)
);

NAND3X1 _18865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf21 ),
    .B(_7898_),
    .C(_7895_),
    .Y(_7899_)
);

AOI21X1 _18866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7892_),
    .B(_7899_),
    .C(\datapath.idinstr_23_bF$buf5 ),
    .Y(_7900_)
);

OAI21X1 _18867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7885_),
    .B(_7900_),
    .C(_7607__bF$buf2),
    .Y(_7901_)
);

MUX2X1 _18868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [6]),
    .B(\datapath.registers.1226[29] [6]),
    .S(\datapath.idinstr_21_bF$buf20 ),
    .Y(_7902_)
);

MUX2X1 _18869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [6]),
    .B(\datapath.registers.1226[28] [6]),
    .S(\datapath.idinstr_21_bF$buf19 ),
    .Y(_7903_)
);

MUX2X1 _18870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7903_),
    .B(_7902_),
    .S(_7608__bF$buf7),
    .Y(_7904_)
);

NAND2X1 _18871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf24 ),
    .B(_7904_),
    .Y(_7905_)
);

MUX2X1 _18872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [6]),
    .B(\datapath.registers.1226[25] [6]),
    .S(\datapath.idinstr_21_bF$buf18 ),
    .Y(_7906_)
);

MUX2X1 _18873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [6]),
    .B(\datapath.registers.1226[24] [6]),
    .S(\datapath.idinstr_21_bF$buf17 ),
    .Y(_7907_)
);

MUX2X1 _18874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7907_),
    .B(_7906_),
    .S(_7608__bF$buf6),
    .Y(_7908_)
);

NAND2X1 _18875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf5),
    .B(_7908_),
    .Y(_7909_)
);

AOI21X1 _18876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7905_),
    .B(_7909_),
    .C(_7612__bF$buf1),
    .Y(_7910_)
);

AOI21X1 _18877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [6]),
    .B(\datapath.idinstr_22_bF$buf23 ),
    .C(_7608__bF$buf5),
    .Y(_7911_)
);

OAI21X1 _18878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6462_),
    .B(\datapath.idinstr_22_bF$buf22 ),
    .C(_7911_),
    .Y(_7912_)
);

AOI21X1 _18879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [6]),
    .B(\datapath.idinstr_22_bF$buf21 ),
    .C(\datapath.idinstr_20_bF$buf18 ),
    .Y(_7913_)
);

OAI21X1 _18880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6465_),
    .B(\datapath.idinstr_22_bF$buf20 ),
    .C(_7913_),
    .Y(_7914_)
);

NAND3X1 _18881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf16 ),
    .B(_7914_),
    .C(_7912_),
    .Y(_7915_)
);

AOI21X1 _18882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [6]),
    .B(\datapath.idinstr_22_bF$buf19 ),
    .C(_7608__bF$buf4),
    .Y(_7916_)
);

OAI21X1 _18883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6469_),
    .B(\datapath.idinstr_22_bF$buf18 ),
    .C(_7916_),
    .Y(_7917_)
);

AOI21X1 _18884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [6]),
    .B(\datapath.idinstr_22_bF$buf17 ),
    .C(\datapath.idinstr_20_bF$buf17 ),
    .Y(_7918_)
);

OAI21X1 _18885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6002_),
    .B(\datapath.idinstr_22_bF$buf16 ),
    .C(_7918_),
    .Y(_7919_)
);

NAND3X1 _18886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf0),
    .B(_7919_),
    .C(_7917_),
    .Y(_7920_)
);

AOI21X1 _18887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7915_),
    .B(_7920_),
    .C(\datapath.idinstr_23_bF$buf4 ),
    .Y(_7921_)
);

OAI21X1 _18888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7910_),
    .B(_7921_),
    .C(\datapath.idinstr_24_bF$buf0 ),
    .Y(_7922_)
);

AOI21X1 _18889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7901_),
    .B(_7922_),
    .C(_7614__bF$buf3),
    .Y(\datapath.registers.regb_data [6])
);

MUX2X1 _18890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [7]),
    .B(\datapath.registers.1226[8] [7]),
    .S(\datapath.idinstr_20_bF$buf16 ),
    .Y(_7923_)
);

MUX2X1 _18891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [7]),
    .B(\datapath.registers.1226[10] [7]),
    .S(\datapath.idinstr_20_bF$buf15 ),
    .Y(_7924_)
);

MUX2X1 _18892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7924_),
    .B(_7923_),
    .S(\datapath.idinstr_21_bF$buf15 ),
    .Y(_7925_)
);

NAND2X1 _18893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf4),
    .B(_7925_),
    .Y(_7926_)
);

MUX2X1 _18894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [7]),
    .B(\datapath.registers.1226[12] [7]),
    .S(\datapath.idinstr_20_bF$buf14 ),
    .Y(_7927_)
);

MUX2X1 _18895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [7]),
    .B(\datapath.registers.1226[14] [7]),
    .S(\datapath.idinstr_20_bF$buf13 ),
    .Y(_7928_)
);

MUX2X1 _18896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7928_),
    .B(_7927_),
    .S(\datapath.idinstr_21_bF$buf14 ),
    .Y(_7929_)
);

NAND2X1 _18897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf15 ),
    .B(_7929_),
    .Y(_7930_)
);

AOI21X1 _18898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7926_),
    .B(_7930_),
    .C(_7612__bF$buf0),
    .Y(_7931_)
);

INVX1 _18899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [7]),
    .Y(_7932_)
);

AOI21X1 _18900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [7]),
    .B(\datapath.idinstr_22_bF$buf14 ),
    .C(_7608__bF$buf3),
    .Y(_7933_)
);

OAI21X1 _18901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7932_),
    .B(\datapath.idinstr_22_bF$buf13 ),
    .C(_7933_),
    .Y(_7934_)
);

NAND2X1 _18902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [7]),
    .B(_7611__bF$buf3),
    .Y(_7935_)
);

AOI21X1 _18903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [7]),
    .B(\datapath.idinstr_22_bF$buf12 ),
    .C(\datapath.idinstr_20_bF$buf12 ),
    .Y(_7936_)
);

AOI21X1 _18904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7936_),
    .B(_7935_),
    .C(\datapath.idinstr_21_bF$buf13 ),
    .Y(_7937_)
);

NAND2X1 _18905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7934_),
    .B(_7937_),
    .Y(_7938_)
);

INVX1 _18906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [7]),
    .Y(_7939_)
);

AOI21X1 _18907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [7]),
    .B(\datapath.idinstr_22_bF$buf11 ),
    .C(_7608__bF$buf2),
    .Y(_7940_)
);

OAI21X1 _18908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7939_),
    .B(\datapath.idinstr_22_bF$buf10 ),
    .C(_7940_),
    .Y(_7941_)
);

INVX1 _18909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[2] [7]),
    .Y(_7942_)
);

AOI21X1 _18910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[6] [7]),
    .B(\datapath.idinstr_22_bF$buf9 ),
    .C(\datapath.idinstr_20_bF$buf11 ),
    .Y(_7943_)
);

OAI21X1 _18911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7942_),
    .B(\datapath.idinstr_22_bF$buf8 ),
    .C(_7943_),
    .Y(_7944_)
);

NAND3X1 _18912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf12 ),
    .B(_7944_),
    .C(_7941_),
    .Y(_7945_)
);

AOI21X1 _18913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7938_),
    .B(_7945_),
    .C(\datapath.idinstr_23_bF$buf3 ),
    .Y(_7946_)
);

OAI21X1 _18914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7931_),
    .B(_7946_),
    .C(_7607__bF$buf1),
    .Y(_7947_)
);

MUX2X1 _18915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [7]),
    .B(\datapath.registers.1226[29] [7]),
    .S(\datapath.idinstr_21_bF$buf11 ),
    .Y(_7948_)
);

MUX2X1 _18916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [7]),
    .B(\datapath.registers.1226[28] [7]),
    .S(\datapath.idinstr_21_bF$buf10 ),
    .Y(_7949_)
);

MUX2X1 _18917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7949_),
    .B(_7948_),
    .S(_7608__bF$buf1),
    .Y(_7950_)
);

NAND2X1 _18918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf7 ),
    .B(_7950_),
    .Y(_7951_)
);

MUX2X1 _18919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [7]),
    .B(\datapath.registers.1226[25] [7]),
    .S(\datapath.idinstr_21_bF$buf9 ),
    .Y(_7952_)
);

MUX2X1 _18920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [7]),
    .B(\datapath.registers.1226[24] [7]),
    .S(\datapath.idinstr_21_bF$buf8 ),
    .Y(_7953_)
);

MUX2X1 _18921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7953_),
    .B(_7952_),
    .S(_7608__bF$buf0),
    .Y(_7954_)
);

NAND2X1 _18922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf2),
    .B(_7954_),
    .Y(_7955_)
);

AOI21X1 _18923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7951_),
    .B(_7955_),
    .C(_7612__bF$buf7),
    .Y(_7956_)
);

INVX1 _18924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [7]),
    .Y(_7957_)
);

AOI21X1 _18925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [7]),
    .B(\datapath.idinstr_22_bF$buf6 ),
    .C(_7608__bF$buf10),
    .Y(_7958_)
);

OAI21X1 _18926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7957_),
    .B(\datapath.idinstr_22_bF$buf5 ),
    .C(_7958_),
    .Y(_7959_)
);

INVX1 _18927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [7]),
    .Y(_7960_)
);

AOI21X1 _18928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [7]),
    .B(\datapath.idinstr_22_bF$buf4 ),
    .C(\datapath.idinstr_20_bF$buf10 ),
    .Y(_7961_)
);

OAI21X1 _18929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7960_),
    .B(\datapath.idinstr_22_bF$buf3 ),
    .C(_7961_),
    .Y(_7962_)
);

NAND3X1 _18930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf7 ),
    .B(_7962_),
    .C(_7959_),
    .Y(_7963_)
);

INVX1 _18931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [7]),
    .Y(_7964_)
);

AOI21X1 _18932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [7]),
    .B(\datapath.idinstr_22_bF$buf2 ),
    .C(_7608__bF$buf9),
    .Y(_7965_)
);

OAI21X1 _18933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7964_),
    .B(\datapath.idinstr_22_bF$buf1 ),
    .C(_7965_),
    .Y(_7966_)
);

AOI21X1 _18934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [7]),
    .B(\datapath.idinstr_22_bF$buf0 ),
    .C(\datapath.idinstr_20_bF$buf9 ),
    .Y(_7967_)
);

OAI21X1 _18935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6004_),
    .B(\datapath.idinstr_22_bF$buf43 ),
    .C(_7967_),
    .Y(_7968_)
);

NAND3X1 _18936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf4),
    .B(_7968_),
    .C(_7966_),
    .Y(_7969_)
);

AOI21X1 _18937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7963_),
    .B(_7969_),
    .C(\datapath.idinstr_23_bF$buf2 ),
    .Y(_7970_)
);

OAI21X1 _18938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7956_),
    .B(_7970_),
    .C(\datapath.idinstr_24_bF$buf5 ),
    .Y(_7971_)
);

AOI21X1 _18939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7947_),
    .B(_7971_),
    .C(_7614__bF$buf2),
    .Y(\datapath.registers.regb_data [7])
);

MUX2X1 _18940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [8]),
    .B(\datapath.registers.1226[24] [8]),
    .S(\datapath.idinstr_20_bF$buf8 ),
    .Y(_7972_)
);

MUX2X1 _18941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [8]),
    .B(\datapath.registers.1226[26] [8]),
    .S(\datapath.idinstr_20_bF$buf7 ),
    .Y(_7973_)
);

MUX2X1 _18942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7973_),
    .B(_7972_),
    .S(\datapath.idinstr_21_bF$buf6 ),
    .Y(_7974_)
);

NAND2X1 _18943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf1),
    .B(_7974_),
    .Y(_7975_)
);

MUX2X1 _18944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [8]),
    .B(\datapath.registers.1226[28] [8]),
    .S(\datapath.idinstr_20_bF$buf6 ),
    .Y(_7976_)
);

MUX2X1 _18945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [8]),
    .B(\datapath.registers.1226[30] [8]),
    .S(\datapath.idinstr_20_bF$buf5 ),
    .Y(_7977_)
);

MUX2X1 _18946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7977_),
    .B(_7976_),
    .S(\datapath.idinstr_21_bF$buf5 ),
    .Y(_7978_)
);

NAND2X1 _18947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf42 ),
    .B(_7978_),
    .Y(_7979_)
);

AOI21X1 _18948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7975_),
    .B(_7979_),
    .C(_7612__bF$buf6),
    .Y(_7980_)
);

MUX2X1 _18949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [8]),
    .B(\datapath.registers.1226[16] [8]),
    .S(\datapath.idinstr_21_bF$buf4 ),
    .Y(_7981_)
);

NAND2X1 _18950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf8),
    .B(_7981_),
    .Y(_7982_)
);

MUX2X1 _18951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [8]),
    .B(\datapath.registers.1226[17] [8]),
    .S(\datapath.idinstr_21_bF$buf3 ),
    .Y(_7983_)
);

AOI21X1 _18952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf4 ),
    .B(_7983_),
    .C(\datapath.idinstr_22_bF$buf41 ),
    .Y(_7984_)
);

NAND2X1 _18953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7982_),
    .B(_7984_),
    .Y(_7985_)
);

MUX2X1 _18954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [8]),
    .B(\datapath.registers.1226[20] [8]),
    .S(\datapath.idinstr_21_bF$buf2 ),
    .Y(_7986_)
);

NAND2X1 _18955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf7),
    .B(_7986_),
    .Y(_7987_)
);

MUX2X1 _18956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [8]),
    .B(\datapath.registers.1226[21] [8]),
    .S(\datapath.idinstr_21_bF$buf1 ),
    .Y(_7988_)
);

AOI21X1 _18957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf3 ),
    .B(_7988_),
    .C(_7611__bF$buf0),
    .Y(_7989_)
);

NAND2X1 _18958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7987_),
    .B(_7989_),
    .Y(_7990_)
);

AOI21X1 _18959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7985_),
    .B(_7990_),
    .C(\datapath.idinstr_23_bF$buf1 ),
    .Y(_7991_)
);

OAI21X1 _18960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7980_),
    .B(_7991_),
    .C(\datapath.idinstr_24_bF$buf4 ),
    .Y(_7992_)
);

MUX2X1 _18961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [8]),
    .B(\datapath.registers.1226[8] [8]),
    .S(\datapath.idinstr_20_bF$buf2 ),
    .Y(_7993_)
);

MUX2X1 _18962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [8]),
    .B(\datapath.registers.1226[10] [8]),
    .S(\datapath.idinstr_20_bF$buf1 ),
    .Y(_7994_)
);

MUX2X1 _18963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7994_),
    .B(_7993_),
    .S(\datapath.idinstr_21_bF$buf0 ),
    .Y(_7995_)
);

NAND2X1 _18964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf10),
    .B(_7995_),
    .Y(_7996_)
);

MUX2X1 _18965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [8]),
    .B(\datapath.registers.1226[12] [8]),
    .S(\datapath.idinstr_20_bF$buf0 ),
    .Y(_7997_)
);

MUX2X1 _18966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [8]),
    .B(\datapath.registers.1226[14] [8]),
    .S(\datapath.idinstr_20_bF$buf55 ),
    .Y(_7998_)
);

MUX2X1 _18967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7998_),
    .B(_7997_),
    .S(\datapath.idinstr_21_bF$buf44 ),
    .Y(_7999_)
);

NAND2X1 _18968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf40 ),
    .B(_7999_),
    .Y(_8000_)
);

AOI21X1 _18969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7996_),
    .B(_8000_),
    .C(_7612__bF$buf5),
    .Y(_8001_)
);

INVX1 _18970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [8]),
    .Y(_8002_)
);

AOI21X1 _18971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [8]),
    .B(\datapath.idinstr_22_bF$buf39 ),
    .C(_7608__bF$buf6),
    .Y(_8003_)
);

OAI21X1 _18972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8002_),
    .B(\datapath.idinstr_22_bF$buf38 ),
    .C(_8003_),
    .Y(_8004_)
);

INVX1 _18973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [8]),
    .Y(_8005_)
);

AOI21X1 _18974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [8]),
    .B(\datapath.idinstr_22_bF$buf37 ),
    .C(\datapath.idinstr_20_bF$buf54 ),
    .Y(_8006_)
);

OAI21X1 _18975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8005_),
    .B(\datapath.idinstr_22_bF$buf36 ),
    .C(_8006_),
    .Y(_8007_)
);

NAND3X1 _18976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf3),
    .B(_8007_),
    .C(_8004_),
    .Y(_8008_)
);

INVX1 _18977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [8]),
    .Y(_8009_)
);

AOI21X1 _18978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [8]),
    .B(\datapath.idinstr_22_bF$buf35 ),
    .C(_7608__bF$buf5),
    .Y(_8010_)
);

OAI21X1 _18979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8009_),
    .B(\datapath.idinstr_22_bF$buf34 ),
    .C(_8010_),
    .Y(_8011_)
);

INVX1 _18980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[2] [8]),
    .Y(_8012_)
);

AOI21X1 _18981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[6] [8]),
    .B(\datapath.idinstr_22_bF$buf33 ),
    .C(\datapath.idinstr_20_bF$buf53 ),
    .Y(_8013_)
);

OAI21X1 _18982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8012_),
    .B(\datapath.idinstr_22_bF$buf32 ),
    .C(_8013_),
    .Y(_8014_)
);

NAND3X1 _18983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf43 ),
    .B(_8014_),
    .C(_8011_),
    .Y(_8015_)
);

AOI21X1 _18984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8008_),
    .B(_8015_),
    .C(\datapath.idinstr_23_bF$buf0 ),
    .Y(_8016_)
);

OAI21X1 _18985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8001_),
    .B(_8016_),
    .C(_7607__bF$buf0),
    .Y(_8017_)
);

AOI21X1 _18986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7992_),
    .B(_8017_),
    .C(_7614__bF$buf1),
    .Y(\datapath.registers.regb_data [8])
);

MUX2X1 _18987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [9]),
    .B(\datapath.registers.1226[24] [9]),
    .S(\datapath.idinstr_20_bF$buf52 ),
    .Y(_8018_)
);

MUX2X1 _18988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [9]),
    .B(\datapath.registers.1226[26] [9]),
    .S(\datapath.idinstr_20_bF$buf51 ),
    .Y(_8019_)
);

MUX2X1 _18989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8019_),
    .B(_8018_),
    .S(\datapath.idinstr_21_bF$buf42 ),
    .Y(_8020_)
);

NAND2X1 _18990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf9),
    .B(_8020_),
    .Y(_8021_)
);

MUX2X1 _18991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [9]),
    .B(\datapath.registers.1226[28] [9]),
    .S(\datapath.idinstr_20_bF$buf50 ),
    .Y(_8022_)
);

MUX2X1 _18992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [9]),
    .B(\datapath.registers.1226[30] [9]),
    .S(\datapath.idinstr_20_bF$buf49 ),
    .Y(_8023_)
);

MUX2X1 _18993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8023_),
    .B(_8022_),
    .S(\datapath.idinstr_21_bF$buf41 ),
    .Y(_8024_)
);

NAND2X1 _18994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf31 ),
    .B(_8024_),
    .Y(_8025_)
);

AOI21X1 _18995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8021_),
    .B(_8025_),
    .C(_7612__bF$buf4),
    .Y(_8026_)
);

MUX2X1 _18996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [9]),
    .B(\datapath.registers.1226[16] [9]),
    .S(\datapath.idinstr_21_bF$buf40 ),
    .Y(_8027_)
);

NAND2X1 _18997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf4),
    .B(_8027_),
    .Y(_8028_)
);

MUX2X1 _18998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [9]),
    .B(\datapath.registers.1226[17] [9]),
    .S(\datapath.idinstr_21_bF$buf39 ),
    .Y(_8029_)
);

AOI21X1 _18999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf48 ),
    .B(_8029_),
    .C(\datapath.idinstr_22_bF$buf30 ),
    .Y(_8030_)
);

NAND2X1 _19000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8028_),
    .B(_8030_),
    .Y(_8031_)
);

MUX2X1 _19001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [9]),
    .B(\datapath.registers.1226[20] [9]),
    .S(\datapath.idinstr_21_bF$buf38 ),
    .Y(_8032_)
);

NAND2X1 _19002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf3),
    .B(_8032_),
    .Y(_8033_)
);

MUX2X1 _19003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [9]),
    .B(\datapath.registers.1226[21] [9]),
    .S(\datapath.idinstr_21_bF$buf37 ),
    .Y(_8034_)
);

AOI21X1 _19004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf47 ),
    .B(_8034_),
    .C(_7611__bF$buf8),
    .Y(_8035_)
);

NAND2X1 _19005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8033_),
    .B(_8035_),
    .Y(_8036_)
);

AOI21X1 _19006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8031_),
    .B(_8036_),
    .C(\datapath.idinstr_23_bF$buf7 ),
    .Y(_8037_)
);

OAI21X1 _19007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8026_),
    .B(_8037_),
    .C(\datapath.idinstr_24_bF$buf3 ),
    .Y(_8038_)
);

MUX2X1 _19008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [9]),
    .B(\datapath.registers.1226[8] [9]),
    .S(\datapath.idinstr_20_bF$buf46 ),
    .Y(_8039_)
);

MUX2X1 _19009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [9]),
    .B(\datapath.registers.1226[10] [9]),
    .S(\datapath.idinstr_20_bF$buf45 ),
    .Y(_8040_)
);

MUX2X1 _19010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8040_),
    .B(_8039_),
    .S(\datapath.idinstr_21_bF$buf36 ),
    .Y(_8041_)
);

NAND2X1 _19011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf7),
    .B(_8041_),
    .Y(_8042_)
);

NOR2X1 _19012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6591_),
    .B(_7608__bF$buf2),
    .Y(_8043_)
);

OAI21X1 _19013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6593_),
    .B(\datapath.idinstr_20_bF$buf44 ),
    .C(\datapath.idinstr_21_bF$buf35 ),
    .Y(_8044_)
);

NAND2X1 _19014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [9]),
    .B(_7608__bF$buf1),
    .Y(_8045_)
);

AOI21X1 _19015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [9]),
    .B(\datapath.idinstr_20_bF$buf43 ),
    .C(\datapath.idinstr_21_bF$buf34 ),
    .Y(_8046_)
);

AOI21X1 _19016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8046_),
    .B(_8045_),
    .C(_7611__bF$buf6),
    .Y(_8047_)
);

OAI21X1 _19017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8043_),
    .B(_8044_),
    .C(_8047_),
    .Y(_8048_)
);

AOI21X1 _19018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8048_),
    .B(_8042_),
    .C(_7612__bF$buf3),
    .Y(_8049_)
);

MUX2X1 _19019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [9]),
    .B(\datapath.registers.1226[4] [9]),
    .S(\datapath.idinstr_20_bF$buf42 ),
    .Y(_8050_)
);

MUX2X1 _19020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [9]),
    .B(\datapath.registers.1226[6] [9]),
    .S(\datapath.idinstr_20_bF$buf41 ),
    .Y(_8051_)
);

MUX2X1 _19021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8051_),
    .B(_8050_),
    .S(\datapath.idinstr_21_bF$buf33 ),
    .Y(_8052_)
);

NAND2X1 _19022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf29 ),
    .B(_8052_),
    .Y(_8053_)
);

MUX2X1 _19023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [9]),
    .B(\datapath.registers.1226[0] [9]),
    .S(\datapath.idinstr_20_bF$buf40 ),
    .Y(_8054_)
);

MUX2X1 _19024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [9]),
    .B(\datapath.registers.1226[2] [9]),
    .S(\datapath.idinstr_20_bF$buf39 ),
    .Y(_8055_)
);

MUX2X1 _19025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8055_),
    .B(_8054_),
    .S(\datapath.idinstr_21_bF$buf32 ),
    .Y(_8056_)
);

NAND2X1 _19026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf5),
    .B(_8056_),
    .Y(_8057_)
);

AOI21X1 _19027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8053_),
    .B(_8057_),
    .C(\datapath.idinstr_23_bF$buf6 ),
    .Y(_8058_)
);

OAI21X1 _19028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8058_),
    .B(_8049_),
    .C(_7607__bF$buf4),
    .Y(_8059_)
);

AOI21X1 _19029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8038_),
    .B(_8059_),
    .C(_7614__bF$buf0),
    .Y(\datapath.registers.regb_data [9])
);

MUX2X1 _19030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [10]),
    .B(\datapath.registers.1226[8] [10]),
    .S(\datapath.idinstr_20_bF$buf38 ),
    .Y(_8060_)
);

MUX2X1 _19031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [10]),
    .B(\datapath.registers.1226[10] [10]),
    .S(\datapath.idinstr_20_bF$buf37 ),
    .Y(_8061_)
);

MUX2X1 _19032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8061_),
    .B(_8060_),
    .S(\datapath.idinstr_21_bF$buf31 ),
    .Y(_8062_)
);

NAND2X1 _19033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf4),
    .B(_8062_),
    .Y(_8063_)
);

NOR2X1 _19034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6614_),
    .B(_7608__bF$buf0),
    .Y(_8064_)
);

OAI21X1 _19035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6616_),
    .B(\datapath.idinstr_20_bF$buf36 ),
    .C(\datapath.idinstr_21_bF$buf30 ),
    .Y(_8065_)
);

NAND2X1 _19036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [10]),
    .B(_7608__bF$buf10),
    .Y(_8066_)
);

AOI21X1 _19037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [10]),
    .B(\datapath.idinstr_20_bF$buf35 ),
    .C(\datapath.idinstr_21_bF$buf29 ),
    .Y(_8067_)
);

AOI21X1 _19038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8067_),
    .B(_8066_),
    .C(_7611__bF$buf3),
    .Y(_8068_)
);

OAI21X1 _19039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8064_),
    .B(_8065_),
    .C(_8068_),
    .Y(_8069_)
);

AOI21X1 _19040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8069_),
    .B(_8063_),
    .C(_7612__bF$buf2),
    .Y(_8070_)
);

MUX2X1 _19041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [10]),
    .B(\datapath.registers.1226[4] [10]),
    .S(\datapath.idinstr_20_bF$buf34 ),
    .Y(_8071_)
);

MUX2X1 _19042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [10]),
    .B(\datapath.registers.1226[6] [10]),
    .S(\datapath.idinstr_20_bF$buf33 ),
    .Y(_8072_)
);

MUX2X1 _19043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8072_),
    .B(_8071_),
    .S(\datapath.idinstr_21_bF$buf28 ),
    .Y(_8073_)
);

NAND2X1 _19044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf28 ),
    .B(_8073_),
    .Y(_8074_)
);

MUX2X1 _19045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [10]),
    .B(\datapath.registers.1226[0] [10]),
    .S(\datapath.idinstr_20_bF$buf32 ),
    .Y(_8075_)
);

MUX2X1 _19046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [10]),
    .B(\datapath.registers.1226[2] [10]),
    .S(\datapath.idinstr_20_bF$buf31 ),
    .Y(_8076_)
);

MUX2X1 _19047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8076_),
    .B(_8075_),
    .S(\datapath.idinstr_21_bF$buf27 ),
    .Y(_8077_)
);

NAND2X1 _19048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf2),
    .B(_8077_),
    .Y(_8078_)
);

AOI21X1 _19049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8074_),
    .B(_8078_),
    .C(\datapath.idinstr_23_bF$buf5 ),
    .Y(_8079_)
);

OAI21X1 _19050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8079_),
    .B(_8070_),
    .C(_7607__bF$buf3),
    .Y(_8080_)
);

INVX1 _19051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [10]),
    .Y(_8081_)
);

AOI21X1 _19052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [10]),
    .B(\datapath.idinstr_22_bF$buf27 ),
    .C(_7608__bF$buf9),
    .Y(_8082_)
);

OAI21X1 _19053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8081_),
    .B(\datapath.idinstr_22_bF$buf26 ),
    .C(_8082_),
    .Y(_8083_)
);

NAND2X1 _19054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [10]),
    .B(_7611__bF$buf1),
    .Y(_8084_)
);

AOI21X1 _19055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [10]),
    .B(\datapath.idinstr_22_bF$buf25 ),
    .C(\datapath.idinstr_20_bF$buf30 ),
    .Y(_8085_)
);

AOI21X1 _19056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8085_),
    .B(_8084_),
    .C(_7610__bF$buf2),
    .Y(_8086_)
);

NAND2X1 _19057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8083_),
    .B(_8086_),
    .Y(_8087_)
);

INVX1 _19058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [10]),
    .Y(_8088_)
);

AOI21X1 _19059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [10]),
    .B(\datapath.idinstr_22_bF$buf24 ),
    .C(_7608__bF$buf8),
    .Y(_8089_)
);

OAI21X1 _19060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8088_),
    .B(\datapath.idinstr_22_bF$buf23 ),
    .C(_8089_),
    .Y(_8090_)
);

AOI21X1 _19061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[28] [10]),
    .B(\datapath.idinstr_22_bF$buf22 ),
    .C(\datapath.idinstr_20_bF$buf29 ),
    .Y(_8091_)
);

OAI21X1 _19062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5727_),
    .B(\datapath.idinstr_22_bF$buf21 ),
    .C(_8091_),
    .Y(_8092_)
);

NAND3X1 _19063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf1),
    .B(_8092_),
    .C(_8090_),
    .Y(_8093_)
);

AOI21X1 _19064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8087_),
    .B(_8093_),
    .C(_7612__bF$buf1),
    .Y(_8094_)
);

MUX2X1 _19065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [10]),
    .B(\datapath.registers.1226[16] [10]),
    .S(\datapath.idinstr_20_bF$buf28 ),
    .Y(_8095_)
);

MUX2X1 _19066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [10]),
    .B(\datapath.registers.1226[18] [10]),
    .S(\datapath.idinstr_20_bF$buf27 ),
    .Y(_8096_)
);

MUX2X1 _19067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8096_),
    .B(_8095_),
    .S(\datapath.idinstr_21_bF$buf26 ),
    .Y(_8097_)
);

NAND2X1 _19068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf0),
    .B(_8097_),
    .Y(_8098_)
);

MUX2X1 _19069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [10]),
    .B(\datapath.registers.1226[20] [10]),
    .S(\datapath.idinstr_20_bF$buf26 ),
    .Y(_8099_)
);

MUX2X1 _19070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [10]),
    .B(\datapath.registers.1226[22] [10]),
    .S(\datapath.idinstr_20_bF$buf25 ),
    .Y(_8100_)
);

MUX2X1 _19071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8100_),
    .B(_8099_),
    .S(\datapath.idinstr_21_bF$buf25 ),
    .Y(_8101_)
);

NAND2X1 _19072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf20 ),
    .B(_8101_),
    .Y(_8102_)
);

AOI21X1 _19073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8098_),
    .B(_8102_),
    .C(\datapath.idinstr_23_bF$buf4 ),
    .Y(_8103_)
);

OAI21X1 _19074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8103_),
    .B(_8094_),
    .C(\datapath.idinstr_24_bF$buf2 ),
    .Y(_8104_)
);

AOI21X1 _19075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8104_),
    .B(_8080_),
    .C(_7614__bF$buf4),
    .Y(\datapath.registers.regb_data [10])
);

MUX2X1 _19076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [11]),
    .B(\datapath.registers.1226[24] [11]),
    .S(\datapath.idinstr_20_bF$buf24 ),
    .Y(_8105_)
);

MUX2X1 _19077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [11]),
    .B(\datapath.registers.1226[26] [11]),
    .S(\datapath.idinstr_20_bF$buf23 ),
    .Y(_8106_)
);

MUX2X1 _19078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8106_),
    .B(_8105_),
    .S(\datapath.idinstr_21_bF$buf24 ),
    .Y(_8107_)
);

NAND2X1 _19079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf10),
    .B(_8107_),
    .Y(_8108_)
);

MUX2X1 _19080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [11]),
    .B(\datapath.registers.1226[28] [11]),
    .S(\datapath.idinstr_20_bF$buf22 ),
    .Y(_8109_)
);

MUX2X1 _19081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [11]),
    .B(\datapath.registers.1226[30] [11]),
    .S(\datapath.idinstr_20_bF$buf21 ),
    .Y(_8110_)
);

MUX2X1 _19082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8110_),
    .B(_8109_),
    .S(\datapath.idinstr_21_bF$buf23 ),
    .Y(_8111_)
);

NAND2X1 _19083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf19 ),
    .B(_8111_),
    .Y(_8112_)
);

AOI21X1 _19084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8108_),
    .B(_8112_),
    .C(_7612__bF$buf0),
    .Y(_8113_)
);

MUX2X1 _19085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [11]),
    .B(\datapath.registers.1226[16] [11]),
    .S(\datapath.idinstr_21_bF$buf22 ),
    .Y(_8114_)
);

NAND2X1 _19086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf7),
    .B(_8114_),
    .Y(_8115_)
);

MUX2X1 _19087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [11]),
    .B(\datapath.registers.1226[17] [11]),
    .S(\datapath.idinstr_21_bF$buf21 ),
    .Y(_8116_)
);

AOI21X1 _19088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf20 ),
    .B(_8116_),
    .C(\datapath.idinstr_22_bF$buf18 ),
    .Y(_8117_)
);

NAND2X1 _19089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8115_),
    .B(_8117_),
    .Y(_8118_)
);

MUX2X1 _19090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [11]),
    .B(\datapath.registers.1226[20] [11]),
    .S(\datapath.idinstr_21_bF$buf20 ),
    .Y(_8119_)
);

NAND2X1 _19091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf6),
    .B(_8119_),
    .Y(_8120_)
);

MUX2X1 _19092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [11]),
    .B(\datapath.registers.1226[21] [11]),
    .S(\datapath.idinstr_21_bF$buf19 ),
    .Y(_8121_)
);

AOI21X1 _19093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf19 ),
    .B(_8121_),
    .C(_7611__bF$buf9),
    .Y(_8122_)
);

NAND2X1 _19094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8120_),
    .B(_8122_),
    .Y(_8123_)
);

AOI21X1 _19095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8118_),
    .B(_8123_),
    .C(\datapath.idinstr_23_bF$buf3 ),
    .Y(_8124_)
);

OAI21X1 _19096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8113_),
    .B(_8124_),
    .C(\datapath.idinstr_24_bF$buf1 ),
    .Y(_8125_)
);

INVX1 _19097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [11]),
    .Y(_8126_)
);

AOI21X1 _19098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [11]),
    .B(\datapath.idinstr_22_bF$buf17 ),
    .C(_7608__bF$buf5),
    .Y(_8127_)
);

OAI21X1 _19099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8126_),
    .B(\datapath.idinstr_22_bF$buf16 ),
    .C(_8127_),
    .Y(_8128_)
);

INVX1 _19100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [11]),
    .Y(_8129_)
);

AOI21X1 _19101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [11]),
    .B(\datapath.idinstr_22_bF$buf15 ),
    .C(\datapath.idinstr_20_bF$buf18 ),
    .Y(_8130_)
);

OAI21X1 _19102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8129_),
    .B(\datapath.idinstr_22_bF$buf14 ),
    .C(_8130_),
    .Y(_8131_)
);

NAND3X1 _19103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf0),
    .B(_8131_),
    .C(_8128_),
    .Y(_8132_)
);

INVX1 _19104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [11]),
    .Y(_8133_)
);

AOI21X1 _19105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [11]),
    .B(\datapath.idinstr_22_bF$buf13 ),
    .C(_7608__bF$buf4),
    .Y(_8134_)
);

OAI21X1 _19106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8133_),
    .B(\datapath.idinstr_22_bF$buf12 ),
    .C(_8134_),
    .Y(_8135_)
);

INVX1 _19107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[10] [11]),
    .Y(_8136_)
);

AOI21X1 _19108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [11]),
    .B(\datapath.idinstr_22_bF$buf11 ),
    .C(\datapath.idinstr_20_bF$buf17 ),
    .Y(_8137_)
);

OAI21X1 _19109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8136_),
    .B(\datapath.idinstr_22_bF$buf10 ),
    .C(_8137_),
    .Y(_8138_)
);

NAND3X1 _19110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf18 ),
    .B(_8138_),
    .C(_8135_),
    .Y(_8139_)
);

AOI21X1 _19111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8132_),
    .B(_8139_),
    .C(_7612__bF$buf7),
    .Y(_8140_)
);

MUX2X1 _19112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [11]),
    .B(\datapath.registers.1226[0] [11]),
    .S(\datapath.idinstr_20_bF$buf16 ),
    .Y(_8141_)
);

MUX2X1 _19113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [11]),
    .B(\datapath.registers.1226[2] [11]),
    .S(\datapath.idinstr_20_bF$buf15 ),
    .Y(_8142_)
);

MUX2X1 _19114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8142_),
    .B(_8141_),
    .S(\datapath.idinstr_21_bF$buf17 ),
    .Y(_8143_)
);

NAND2X1 _19115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf8),
    .B(_8143_),
    .Y(_8144_)
);

MUX2X1 _19116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [11]),
    .B(\datapath.registers.1226[4] [11]),
    .S(\datapath.idinstr_20_bF$buf14 ),
    .Y(_8145_)
);

MUX2X1 _19117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [11]),
    .B(\datapath.registers.1226[6] [11]),
    .S(\datapath.idinstr_20_bF$buf13 ),
    .Y(_8146_)
);

MUX2X1 _19118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8146_),
    .B(_8145_),
    .S(\datapath.idinstr_21_bF$buf16 ),
    .Y(_8147_)
);

NAND2X1 _19119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf9 ),
    .B(_8147_),
    .Y(_8148_)
);

AOI21X1 _19120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8144_),
    .B(_8148_),
    .C(\datapath.idinstr_23_bF$buf2 ),
    .Y(_8149_)
);

OAI21X1 _19121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8149_),
    .B(_8140_),
    .C(_7607__bF$buf2),
    .Y(_8150_)
);

AOI21X1 _19122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8125_),
    .B(_8150_),
    .C(_7614__bF$buf3),
    .Y(\datapath.registers.regb_data [11])
);

MUX2X1 _19123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [12]),
    .B(\datapath.registers.1226[8] [12]),
    .S(\datapath.idinstr_20_bF$buf12 ),
    .Y(_8151_)
);

MUX2X1 _19124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [12]),
    .B(\datapath.registers.1226[10] [12]),
    .S(\datapath.idinstr_20_bF$buf11 ),
    .Y(_8152_)
);

MUX2X1 _19125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8152_),
    .B(_8151_),
    .S(\datapath.idinstr_21_bF$buf15 ),
    .Y(_8153_)
);

NAND2X1 _19126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf7),
    .B(_8153_),
    .Y(_8154_)
);

AND2X2 _19127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [12]),
    .B(\datapath.idinstr_20_bF$buf10 ),
    .Y(_8155_)
);

INVX1 _19128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [12]),
    .Y(_8156_)
);

OAI21X1 _19129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8156_),
    .B(\datapath.idinstr_20_bF$buf9 ),
    .C(\datapath.idinstr_21_bF$buf14 ),
    .Y(_8157_)
);

NAND2X1 _19130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [12]),
    .B(_7608__bF$buf3),
    .Y(_8158_)
);

AOI21X1 _19131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [12]),
    .B(\datapath.idinstr_20_bF$buf8 ),
    .C(\datapath.idinstr_21_bF$buf13 ),
    .Y(_8159_)
);

AOI21X1 _19132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8159_),
    .B(_8158_),
    .C(_7611__bF$buf6),
    .Y(_8160_)
);

OAI21X1 _19133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8155_),
    .B(_8157_),
    .C(_8160_),
    .Y(_8161_)
);

AOI21X1 _19134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8161_),
    .B(_8154_),
    .C(_7612__bF$buf6),
    .Y(_8162_)
);

MUX2X1 _19135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [12]),
    .B(\datapath.registers.1226[4] [12]),
    .S(\datapath.idinstr_20_bF$buf7 ),
    .Y(_8163_)
);

MUX2X1 _19136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [12]),
    .B(\datapath.registers.1226[6] [12]),
    .S(\datapath.idinstr_20_bF$buf6 ),
    .Y(_8164_)
);

MUX2X1 _19137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8164_),
    .B(_8163_),
    .S(\datapath.idinstr_21_bF$buf12 ),
    .Y(_8165_)
);

NAND2X1 _19138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf8 ),
    .B(_8165_),
    .Y(_8166_)
);

MUX2X1 _19139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [12]),
    .B(\datapath.registers.1226[0] [12]),
    .S(\datapath.idinstr_20_bF$buf5 ),
    .Y(_8167_)
);

MUX2X1 _19140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [12]),
    .B(\datapath.registers.1226[2] [12]),
    .S(\datapath.idinstr_20_bF$buf4 ),
    .Y(_8168_)
);

MUX2X1 _19141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8168_),
    .B(_8167_),
    .S(\datapath.idinstr_21_bF$buf11 ),
    .Y(_8169_)
);

NAND2X1 _19142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf5),
    .B(_8169_),
    .Y(_8170_)
);

AOI21X1 _19143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8166_),
    .B(_8170_),
    .C(\datapath.idinstr_23_bF$buf1 ),
    .Y(_8171_)
);

OAI21X1 _19144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8171_),
    .B(_8162_),
    .C(_7607__bF$buf1),
    .Y(_8172_)
);

INVX1 _19145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [12]),
    .Y(_8173_)
);

AOI21X1 _19146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [12]),
    .B(\datapath.idinstr_22_bF$buf7 ),
    .C(_7608__bF$buf2),
    .Y(_8174_)
);

OAI21X1 _19147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8173_),
    .B(\datapath.idinstr_22_bF$buf6 ),
    .C(_8174_),
    .Y(_8175_)
);

NAND2X1 _19148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [12]),
    .B(_7611__bF$buf4),
    .Y(_8176_)
);

AOI21X1 _19149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [12]),
    .B(\datapath.idinstr_22_bF$buf5 ),
    .C(\datapath.idinstr_20_bF$buf3 ),
    .Y(_8177_)
);

AOI21X1 _19150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8177_),
    .B(_8176_),
    .C(_7610__bF$buf4),
    .Y(_8178_)
);

NAND2X1 _19151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8175_),
    .B(_8178_),
    .Y(_8179_)
);

INVX1 _19152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [12]),
    .Y(_8180_)
);

AOI21X1 _19153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [12]),
    .B(\datapath.idinstr_22_bF$buf4 ),
    .C(_7608__bF$buf1),
    .Y(_8181_)
);

OAI21X1 _19154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8180_),
    .B(\datapath.idinstr_22_bF$buf3 ),
    .C(_8181_),
    .Y(_8182_)
);

AOI21X1 _19155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [12]),
    .B(\datapath.idinstr_22_bF$buf2 ),
    .C(\datapath.idinstr_20_bF$buf2 ),
    .Y(_8183_)
);

OAI21X1 _19156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6012_),
    .B(\datapath.idinstr_22_bF$buf1 ),
    .C(_8183_),
    .Y(_8184_)
);

NAND3X1 _19157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf3),
    .B(_8184_),
    .C(_8182_),
    .Y(_8185_)
);

AOI21X1 _19158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8179_),
    .B(_8185_),
    .C(\datapath.idinstr_23_bF$buf0 ),
    .Y(_8186_)
);

MUX2X1 _19159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [12]),
    .B(\datapath.registers.1226[29] [12]),
    .S(\datapath.idinstr_21_bF$buf10 ),
    .Y(_8187_)
);

MUX2X1 _19160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [12]),
    .B(\datapath.registers.1226[28] [12]),
    .S(\datapath.idinstr_21_bF$buf9 ),
    .Y(_8188_)
);

MUX2X1 _19161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8188_),
    .B(_8187_),
    .S(_7608__bF$buf0),
    .Y(_8189_)
);

NAND2X1 _19162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf0 ),
    .B(_8189_),
    .Y(_8190_)
);

MUX2X1 _19163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [12]),
    .B(\datapath.registers.1226[25] [12]),
    .S(\datapath.idinstr_21_bF$buf8 ),
    .Y(_8191_)
);

MUX2X1 _19164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [12]),
    .B(\datapath.registers.1226[24] [12]),
    .S(\datapath.idinstr_21_bF$buf7 ),
    .Y(_8192_)
);

MUX2X1 _19165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8192_),
    .B(_8191_),
    .S(_7608__bF$buf10),
    .Y(_8193_)
);

NAND2X1 _19166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf3),
    .B(_8193_),
    .Y(_8194_)
);

AOI21X1 _19167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8190_),
    .B(_8194_),
    .C(_7612__bF$buf5),
    .Y(_8195_)
);

OAI21X1 _19168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8195_),
    .B(_8186_),
    .C(\datapath.idinstr_24_bF$buf0 ),
    .Y(_8196_)
);

AOI21X1 _19169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8196_),
    .B(_8172_),
    .C(_7614__bF$buf2),
    .Y(\datapath.registers.regb_data [12])
);

MUX2X1 _19170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [13]),
    .B(\datapath.registers.1226[0] [13]),
    .S(\datapath.idinstr_20_bF$buf1 ),
    .Y(_8197_)
);

MUX2X1 _19171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [13]),
    .B(\datapath.registers.1226[2] [13]),
    .S(\datapath.idinstr_20_bF$buf0 ),
    .Y(_8198_)
);

MUX2X1 _19172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8198_),
    .B(_8197_),
    .S(\datapath.idinstr_21_bF$buf6 ),
    .Y(_8199_)
);

NAND2X1 _19173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf2),
    .B(_8199_),
    .Y(_8200_)
);

MUX2X1 _19174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [13]),
    .B(\datapath.registers.1226[4] [13]),
    .S(\datapath.idinstr_20_bF$buf55 ),
    .Y(_8201_)
);

MUX2X1 _19175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [13]),
    .B(\datapath.registers.1226[6] [13]),
    .S(\datapath.idinstr_20_bF$buf54 ),
    .Y(_8202_)
);

MUX2X1 _19176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8202_),
    .B(_8201_),
    .S(\datapath.idinstr_21_bF$buf5 ),
    .Y(_8203_)
);

NAND2X1 _19177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf43 ),
    .B(_8203_),
    .Y(_8204_)
);

AOI21X1 _19178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8200_),
    .B(_8204_),
    .C(\datapath.idinstr_23_bF$buf7 ),
    .Y(_8205_)
);

AOI21X1 _19179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [13]),
    .B(\datapath.idinstr_22_bF$buf42 ),
    .C(_7608__bF$buf9),
    .Y(_8206_)
);

OAI21X1 _19180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6767_),
    .B(\datapath.idinstr_22_bF$buf41 ),
    .C(_8206_),
    .Y(_8207_)
);

NAND2X1 _19181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [13]),
    .B(_7611__bF$buf1),
    .Y(_8208_)
);

AOI21X1 _19182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [13]),
    .B(\datapath.idinstr_22_bF$buf40 ),
    .C(\datapath.idinstr_20_bF$buf53 ),
    .Y(_8209_)
);

AOI21X1 _19183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8209_),
    .B(_8208_),
    .C(\datapath.idinstr_21_bF$buf4 ),
    .Y(_8210_)
);

NAND2X1 _19184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8207_),
    .B(_8210_),
    .Y(_8211_)
);

AOI21X1 _19185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [13]),
    .B(\datapath.idinstr_22_bF$buf39 ),
    .C(_7608__bF$buf8),
    .Y(_8212_)
);

OAI21X1 _19186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6774_),
    .B(\datapath.idinstr_22_bF$buf38 ),
    .C(_8212_),
    .Y(_8213_)
);

AOI21X1 _19187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [13]),
    .B(\datapath.idinstr_22_bF$buf37 ),
    .C(\datapath.idinstr_20_bF$buf52 ),
    .Y(_8214_)
);

OAI21X1 _19188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6777_),
    .B(\datapath.idinstr_22_bF$buf36 ),
    .C(_8214_),
    .Y(_8215_)
);

NAND3X1 _19189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf3 ),
    .B(_8215_),
    .C(_8213_),
    .Y(_8216_)
);

AOI21X1 _19190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8211_),
    .B(_8216_),
    .C(_7612__bF$buf4),
    .Y(_8217_)
);

OAI21X1 _19191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8205_),
    .B(_8217_),
    .C(_7607__bF$buf0),
    .Y(_8218_)
);

MUX2X1 _19192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [13]),
    .B(\datapath.registers.1226[29] [13]),
    .S(\datapath.idinstr_21_bF$buf2 ),
    .Y(_8219_)
);

MUX2X1 _19193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [13]),
    .B(\datapath.registers.1226[28] [13]),
    .S(\datapath.idinstr_21_bF$buf1 ),
    .Y(_8220_)
);

MUX2X1 _19194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8220_),
    .B(_8219_),
    .S(_7608__bF$buf7),
    .Y(_8221_)
);

NAND2X1 _19195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf35 ),
    .B(_8221_),
    .Y(_8222_)
);

MUX2X1 _19196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [13]),
    .B(\datapath.registers.1226[25] [13]),
    .S(\datapath.idinstr_21_bF$buf0 ),
    .Y(_8223_)
);

MUX2X1 _19197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [13]),
    .B(\datapath.registers.1226[24] [13]),
    .S(\datapath.idinstr_21_bF$buf44 ),
    .Y(_8224_)
);

MUX2X1 _19198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8224_),
    .B(_8223_),
    .S(_7608__bF$buf6),
    .Y(_8225_)
);

NAND2X1 _19199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf0),
    .B(_8225_),
    .Y(_8226_)
);

AOI21X1 _19200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8222_),
    .B(_8226_),
    .C(_7612__bF$buf3),
    .Y(_8227_)
);

INVX1 _19201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [13]),
    .Y(_8228_)
);

AOI21X1 _19202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [13]),
    .B(\datapath.idinstr_22_bF$buf34 ),
    .C(_7608__bF$buf5),
    .Y(_8229_)
);

OAI21X1 _19203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8228_),
    .B(\datapath.idinstr_22_bF$buf33 ),
    .C(_8229_),
    .Y(_8230_)
);

INVX1 _19204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [13]),
    .Y(_8231_)
);

AOI21X1 _19205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [13]),
    .B(\datapath.idinstr_22_bF$buf32 ),
    .C(\datapath.idinstr_20_bF$buf51 ),
    .Y(_8232_)
);

OAI21X1 _19206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8231_),
    .B(\datapath.idinstr_22_bF$buf31 ),
    .C(_8232_),
    .Y(_8233_)
);

NAND3X1 _19207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf43 ),
    .B(_8233_),
    .C(_8230_),
    .Y(_8234_)
);

INVX1 _19208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [13]),
    .Y(_8235_)
);

AOI21X1 _19209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [13]),
    .B(\datapath.idinstr_22_bF$buf30 ),
    .C(_7608__bF$buf4),
    .Y(_8236_)
);

OAI21X1 _19210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8235_),
    .B(\datapath.idinstr_22_bF$buf29 ),
    .C(_8236_),
    .Y(_8237_)
);

AOI21X1 _19211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [13]),
    .B(\datapath.idinstr_22_bF$buf28 ),
    .C(\datapath.idinstr_20_bF$buf50 ),
    .Y(_8238_)
);

OAI21X1 _19212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6014_),
    .B(\datapath.idinstr_22_bF$buf27 ),
    .C(_8238_),
    .Y(_8239_)
);

NAND3X1 _19213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf2),
    .B(_8239_),
    .C(_8237_),
    .Y(_8240_)
);

AOI21X1 _19214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8234_),
    .B(_8240_),
    .C(\datapath.idinstr_23_bF$buf6 ),
    .Y(_8241_)
);

OAI21X1 _19215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8227_),
    .B(_8241_),
    .C(\datapath.idinstr_24_bF$buf5 ),
    .Y(_8242_)
);

AOI21X1 _19216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8218_),
    .B(_8242_),
    .C(_7614__bF$buf1),
    .Y(\datapath.registers.regb_data [13])
);

MUX2X1 _19217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [14]),
    .B(\datapath.registers.1226[24] [14]),
    .S(\datapath.idinstr_20_bF$buf49 ),
    .Y(_8243_)
);

MUX2X1 _19218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [14]),
    .B(\datapath.registers.1226[26] [14]),
    .S(\datapath.idinstr_20_bF$buf48 ),
    .Y(_8244_)
);

MUX2X1 _19219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8244_),
    .B(_8243_),
    .S(\datapath.idinstr_21_bF$buf42 ),
    .Y(_8245_)
);

NAND2X1 _19220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf10),
    .B(_8245_),
    .Y(_8246_)
);

MUX2X1 _19221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [14]),
    .B(\datapath.registers.1226[28] [14]),
    .S(\datapath.idinstr_20_bF$buf47 ),
    .Y(_8247_)
);

MUX2X1 _19222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [14]),
    .B(\datapath.registers.1226[30] [14]),
    .S(\datapath.idinstr_20_bF$buf46 ),
    .Y(_8248_)
);

MUX2X1 _19223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8248_),
    .B(_8247_),
    .S(\datapath.idinstr_21_bF$buf41 ),
    .Y(_8249_)
);

NAND2X1 _19224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf26 ),
    .B(_8249_),
    .Y(_8250_)
);

AOI21X1 _19225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8246_),
    .B(_8250_),
    .C(_7612__bF$buf2),
    .Y(_8251_)
);

MUX2X1 _19226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [14]),
    .B(\datapath.registers.1226[16] [14]),
    .S(\datapath.idinstr_21_bF$buf40 ),
    .Y(_8252_)
);

NAND2X1 _19227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf3),
    .B(_8252_),
    .Y(_8253_)
);

MUX2X1 _19228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [14]),
    .B(\datapath.registers.1226[17] [14]),
    .S(\datapath.idinstr_21_bF$buf39 ),
    .Y(_8254_)
);

AOI21X1 _19229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf45 ),
    .B(_8254_),
    .C(\datapath.idinstr_22_bF$buf25 ),
    .Y(_8255_)
);

NAND2X1 _19230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8253_),
    .B(_8255_),
    .Y(_8256_)
);

MUX2X1 _19231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [14]),
    .B(\datapath.registers.1226[20] [14]),
    .S(\datapath.idinstr_21_bF$buf38 ),
    .Y(_8257_)
);

NAND2X1 _19232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf2),
    .B(_8257_),
    .Y(_8258_)
);

MUX2X1 _19233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [14]),
    .B(\datapath.registers.1226[21] [14]),
    .S(\datapath.idinstr_21_bF$buf37 ),
    .Y(_8259_)
);

AOI21X1 _19234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf44 ),
    .B(_8259_),
    .C(_7611__bF$buf9),
    .Y(_8260_)
);

NAND2X1 _19235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8258_),
    .B(_8260_),
    .Y(_8261_)
);

AOI21X1 _19236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8256_),
    .B(_8261_),
    .C(\datapath.idinstr_23_bF$buf5 ),
    .Y(_8262_)
);

OAI21X1 _19237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8251_),
    .B(_8262_),
    .C(\datapath.idinstr_24_bF$buf4 ),
    .Y(_8263_)
);

MUX2X1 _19238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [14]),
    .B(\datapath.registers.1226[8] [14]),
    .S(\datapath.idinstr_20_bF$buf43 ),
    .Y(_8264_)
);

MUX2X1 _19239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [14]),
    .B(\datapath.registers.1226[10] [14]),
    .S(\datapath.idinstr_20_bF$buf42 ),
    .Y(_8265_)
);

MUX2X1 _19240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8265_),
    .B(_8264_),
    .S(\datapath.idinstr_21_bF$buf36 ),
    .Y(_8266_)
);

NAND2X1 _19241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf8),
    .B(_8266_),
    .Y(_8267_)
);

MUX2X1 _19242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [14]),
    .B(\datapath.registers.1226[12] [14]),
    .S(\datapath.idinstr_20_bF$buf41 ),
    .Y(_8268_)
);

MUX2X1 _19243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [14]),
    .B(\datapath.registers.1226[14] [14]),
    .S(\datapath.idinstr_20_bF$buf40 ),
    .Y(_8269_)
);

MUX2X1 _19244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8269_),
    .B(_8268_),
    .S(\datapath.idinstr_21_bF$buf35 ),
    .Y(_8270_)
);

NAND2X1 _19245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf24 ),
    .B(_8270_),
    .Y(_8271_)
);

AOI21X1 _19246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8267_),
    .B(_8271_),
    .C(_7612__bF$buf1),
    .Y(_8272_)
);

INVX1 _19247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [14]),
    .Y(_8273_)
);

AOI21X1 _19248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [14]),
    .B(\datapath.idinstr_22_bF$buf23 ),
    .C(_7608__bF$buf1),
    .Y(_8274_)
);

OAI21X1 _19249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8273_),
    .B(\datapath.idinstr_22_bF$buf22 ),
    .C(_8274_),
    .Y(_8275_)
);

INVX1 _19250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [14]),
    .Y(_8276_)
);

AOI21X1 _19251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [14]),
    .B(\datapath.idinstr_22_bF$buf21 ),
    .C(\datapath.idinstr_20_bF$buf39 ),
    .Y(_8277_)
);

OAI21X1 _19252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8276_),
    .B(\datapath.idinstr_22_bF$buf20 ),
    .C(_8277_),
    .Y(_8278_)
);

NAND3X1 _19253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf1),
    .B(_8278_),
    .C(_8275_),
    .Y(_8279_)
);

INVX1 _19254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [14]),
    .Y(_8280_)
);

AOI21X1 _19255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [14]),
    .B(\datapath.idinstr_22_bF$buf19 ),
    .C(_7608__bF$buf0),
    .Y(_8281_)
);

OAI21X1 _19256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8280_),
    .B(\datapath.idinstr_22_bF$buf18 ),
    .C(_8281_),
    .Y(_8282_)
);

INVX1 _19257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[2] [14]),
    .Y(_8283_)
);

AOI21X1 _19258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[6] [14]),
    .B(\datapath.idinstr_22_bF$buf17 ),
    .C(\datapath.idinstr_20_bF$buf38 ),
    .Y(_8284_)
);

OAI21X1 _19259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8283_),
    .B(\datapath.idinstr_22_bF$buf16 ),
    .C(_8284_),
    .Y(_8285_)
);

NAND3X1 _19260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf34 ),
    .B(_8285_),
    .C(_8282_),
    .Y(_8286_)
);

AOI21X1 _19261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8279_),
    .B(_8286_),
    .C(\datapath.idinstr_23_bF$buf4 ),
    .Y(_8287_)
);

OAI21X1 _19262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8272_),
    .B(_8287_),
    .C(_7607__bF$buf4),
    .Y(_8288_)
);

AOI21X1 _19263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8263_),
    .B(_8288_),
    .C(_7614__bF$buf0),
    .Y(\datapath.registers.regb_data [14])
);

MUX2X1 _19264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [15]),
    .B(\datapath.registers.1226[24] [15]),
    .S(\datapath.idinstr_20_bF$buf37 ),
    .Y(_8289_)
);

MUX2X1 _19265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [15]),
    .B(\datapath.registers.1226[26] [15]),
    .S(\datapath.idinstr_20_bF$buf36 ),
    .Y(_8290_)
);

MUX2X1 _19266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8290_),
    .B(_8289_),
    .S(\datapath.idinstr_21_bF$buf33 ),
    .Y(_8291_)
);

NAND2X1 _19267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf7),
    .B(_8291_),
    .Y(_8292_)
);

MUX2X1 _19268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [15]),
    .B(\datapath.registers.1226[28] [15]),
    .S(\datapath.idinstr_20_bF$buf35 ),
    .Y(_8293_)
);

MUX2X1 _19269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [15]),
    .B(\datapath.registers.1226[30] [15]),
    .S(\datapath.idinstr_20_bF$buf34 ),
    .Y(_8294_)
);

MUX2X1 _19270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8294_),
    .B(_8293_),
    .S(\datapath.idinstr_21_bF$buf32 ),
    .Y(_8295_)
);

NAND2X1 _19271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf15 ),
    .B(_8295_),
    .Y(_8296_)
);

AOI21X1 _19272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8292_),
    .B(_8296_),
    .C(_7612__bF$buf0),
    .Y(_8297_)
);

MUX2X1 _19273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [15]),
    .B(\datapath.registers.1226[16] [15]),
    .S(\datapath.idinstr_21_bF$buf31 ),
    .Y(_8298_)
);

NAND2X1 _19274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf10),
    .B(_8298_),
    .Y(_8299_)
);

MUX2X1 _19275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [15]),
    .B(\datapath.registers.1226[17] [15]),
    .S(\datapath.idinstr_21_bF$buf30 ),
    .Y(_8300_)
);

AOI21X1 _19276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf33 ),
    .B(_8300_),
    .C(\datapath.idinstr_22_bF$buf14 ),
    .Y(_8301_)
);

NAND2X1 _19277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8299_),
    .B(_8301_),
    .Y(_8302_)
);

MUX2X1 _19278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [15]),
    .B(\datapath.registers.1226[20] [15]),
    .S(\datapath.idinstr_21_bF$buf29 ),
    .Y(_8303_)
);

NAND2X1 _19279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf9),
    .B(_8303_),
    .Y(_8304_)
);

MUX2X1 _19280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [15]),
    .B(\datapath.registers.1226[21] [15]),
    .S(\datapath.idinstr_21_bF$buf28 ),
    .Y(_8305_)
);

AOI21X1 _19281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf32 ),
    .B(_8305_),
    .C(_7611__bF$buf6),
    .Y(_8306_)
);

NAND2X1 _19282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8304_),
    .B(_8306_),
    .Y(_8307_)
);

AOI21X1 _19283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8302_),
    .B(_8307_),
    .C(\datapath.idinstr_23_bF$buf3 ),
    .Y(_8308_)
);

OAI21X1 _19284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8297_),
    .B(_8308_),
    .C(\datapath.idinstr_24_bF$buf3 ),
    .Y(_8309_)
);

MUX2X1 _19285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [15]),
    .B(\datapath.registers.1226[8] [15]),
    .S(\datapath.idinstr_20_bF$buf31 ),
    .Y(_8310_)
);

MUX2X1 _19286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [15]),
    .B(\datapath.registers.1226[10] [15]),
    .S(\datapath.idinstr_20_bF$buf30 ),
    .Y(_8311_)
);

MUX2X1 _19287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8311_),
    .B(_8310_),
    .S(\datapath.idinstr_21_bF$buf27 ),
    .Y(_8312_)
);

NAND2X1 _19288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf5),
    .B(_8312_),
    .Y(_8313_)
);

NOR2X1 _19289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6860_),
    .B(_7608__bF$buf8),
    .Y(_8314_)
);

OAI21X1 _19290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6862_),
    .B(\datapath.idinstr_20_bF$buf29 ),
    .C(\datapath.idinstr_21_bF$buf26 ),
    .Y(_8315_)
);

NAND2X1 _19291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [15]),
    .B(_7608__bF$buf7),
    .Y(_8316_)
);

AOI21X1 _19292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [15]),
    .B(\datapath.idinstr_20_bF$buf28 ),
    .C(\datapath.idinstr_21_bF$buf25 ),
    .Y(_8317_)
);

AOI21X1 _19293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8317_),
    .B(_8316_),
    .C(_7611__bF$buf4),
    .Y(_8318_)
);

OAI21X1 _19294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8314_),
    .B(_8315_),
    .C(_8318_),
    .Y(_8319_)
);

AOI21X1 _19295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8319_),
    .B(_8313_),
    .C(_7612__bF$buf7),
    .Y(_8320_)
);

MUX2X1 _19296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [15]),
    .B(\datapath.registers.1226[4] [15]),
    .S(\datapath.idinstr_20_bF$buf27 ),
    .Y(_8321_)
);

MUX2X1 _19297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [15]),
    .B(\datapath.registers.1226[6] [15]),
    .S(\datapath.idinstr_20_bF$buf26 ),
    .Y(_8322_)
);

MUX2X1 _19298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8322_),
    .B(_8321_),
    .S(\datapath.idinstr_21_bF$buf24 ),
    .Y(_8323_)
);

NAND2X1 _19299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf13 ),
    .B(_8323_),
    .Y(_8324_)
);

MUX2X1 _19300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [15]),
    .B(\datapath.registers.1226[0] [15]),
    .S(\datapath.idinstr_20_bF$buf25 ),
    .Y(_8325_)
);

MUX2X1 _19301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [15]),
    .B(\datapath.registers.1226[2] [15]),
    .S(\datapath.idinstr_20_bF$buf24 ),
    .Y(_8326_)
);

MUX2X1 _19302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8326_),
    .B(_8325_),
    .S(\datapath.idinstr_21_bF$buf23 ),
    .Y(_8327_)
);

NAND2X1 _19303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf3),
    .B(_8327_),
    .Y(_8328_)
);

AOI21X1 _19304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8324_),
    .B(_8328_),
    .C(\datapath.idinstr_23_bF$buf2 ),
    .Y(_8329_)
);

OAI21X1 _19305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8329_),
    .B(_8320_),
    .C(_7607__bF$buf3),
    .Y(_8330_)
);

AOI21X1 _19306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8309_),
    .B(_8330_),
    .C(_7614__bF$buf4),
    .Y(\datapath.registers.regb_data [15])
);

MUX2X1 _19307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [16]),
    .B(\datapath.registers.1226[8] [16]),
    .S(\datapath.idinstr_20_bF$buf23 ),
    .Y(_8331_)
);

MUX2X1 _19308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [16]),
    .B(\datapath.registers.1226[10] [16]),
    .S(\datapath.idinstr_20_bF$buf22 ),
    .Y(_8332_)
);

MUX2X1 _19309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8332_),
    .B(_8331_),
    .S(\datapath.idinstr_21_bF$buf22 ),
    .Y(_8333_)
);

NAND2X1 _19310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf2),
    .B(_8333_),
    .Y(_8334_)
);

NOR2X1 _19311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6883_),
    .B(_7608__bF$buf6),
    .Y(_8335_)
);

OAI21X1 _19312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6885_),
    .B(\datapath.idinstr_20_bF$buf21 ),
    .C(\datapath.idinstr_21_bF$buf21 ),
    .Y(_8336_)
);

NAND2X1 _19313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [16]),
    .B(_7608__bF$buf5),
    .Y(_8337_)
);

AOI21X1 _19314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [16]),
    .B(\datapath.idinstr_20_bF$buf20 ),
    .C(\datapath.idinstr_21_bF$buf20 ),
    .Y(_8338_)
);

AOI21X1 _19315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8338_),
    .B(_8337_),
    .C(_7611__bF$buf1),
    .Y(_8339_)
);

OAI21X1 _19316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8335_),
    .B(_8336_),
    .C(_8339_),
    .Y(_8340_)
);

AOI21X1 _19317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8340_),
    .B(_8334_),
    .C(_7612__bF$buf6),
    .Y(_8341_)
);

MUX2X1 _19318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [16]),
    .B(\datapath.registers.1226[4] [16]),
    .S(\datapath.idinstr_20_bF$buf19 ),
    .Y(_8342_)
);

MUX2X1 _19319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [16]),
    .B(\datapath.registers.1226[6] [16]),
    .S(\datapath.idinstr_20_bF$buf18 ),
    .Y(_8343_)
);

MUX2X1 _19320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8343_),
    .B(_8342_),
    .S(\datapath.idinstr_21_bF$buf19 ),
    .Y(_8344_)
);

NAND2X1 _19321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf12 ),
    .B(_8344_),
    .Y(_8345_)
);

MUX2X1 _19322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [16]),
    .B(\datapath.registers.1226[0] [16]),
    .S(\datapath.idinstr_20_bF$buf17 ),
    .Y(_8346_)
);

MUX2X1 _19323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [16]),
    .B(\datapath.registers.1226[2] [16]),
    .S(\datapath.idinstr_20_bF$buf16 ),
    .Y(_8347_)
);

MUX2X1 _19324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8347_),
    .B(_8346_),
    .S(\datapath.idinstr_21_bF$buf18 ),
    .Y(_8348_)
);

NAND2X1 _19325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf0),
    .B(_8348_),
    .Y(_8349_)
);

AOI21X1 _19326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8345_),
    .B(_8349_),
    .C(\datapath.idinstr_23_bF$buf1 ),
    .Y(_8350_)
);

OAI21X1 _19327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8350_),
    .B(_8341_),
    .C(_7607__bF$buf2),
    .Y(_8351_)
);

INVX1 _19328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [16]),
    .Y(_8352_)
);

AOI21X1 _19329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [16]),
    .B(\datapath.idinstr_22_bF$buf11 ),
    .C(_7608__bF$buf4),
    .Y(_8353_)
);

OAI21X1 _19330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8352_),
    .B(\datapath.idinstr_22_bF$buf10 ),
    .C(_8353_),
    .Y(_8354_)
);

NAND2X1 _19331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [16]),
    .B(_7611__bF$buf10),
    .Y(_8355_)
);

AOI21X1 _19332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [16]),
    .B(\datapath.idinstr_22_bF$buf9 ),
    .C(\datapath.idinstr_20_bF$buf15 ),
    .Y(_8356_)
);

AOI21X1 _19333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8356_),
    .B(_8355_),
    .C(_7610__bF$buf0),
    .Y(_8357_)
);

NAND2X1 _19334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8354_),
    .B(_8357_),
    .Y(_8358_)
);

INVX1 _19335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [16]),
    .Y(_8359_)
);

AOI21X1 _19336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [16]),
    .B(\datapath.idinstr_22_bF$buf8 ),
    .C(_7608__bF$buf3),
    .Y(_8360_)
);

OAI21X1 _19337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8359_),
    .B(\datapath.idinstr_22_bF$buf7 ),
    .C(_8360_),
    .Y(_8361_)
);

AOI21X1 _19338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[28] [16]),
    .B(\datapath.idinstr_22_bF$buf6 ),
    .C(\datapath.idinstr_20_bF$buf14 ),
    .Y(_8362_)
);

OAI21X1 _19339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5734_),
    .B(\datapath.idinstr_22_bF$buf5 ),
    .C(_8362_),
    .Y(_8363_)
);

NAND3X1 _19340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf4),
    .B(_8363_),
    .C(_8361_),
    .Y(_8364_)
);

AOI21X1 _19341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8358_),
    .B(_8364_),
    .C(_7612__bF$buf5),
    .Y(_8365_)
);

MUX2X1 _19342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [16]),
    .B(\datapath.registers.1226[16] [16]),
    .S(\datapath.idinstr_20_bF$buf13 ),
    .Y(_8366_)
);

MUX2X1 _19343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [16]),
    .B(\datapath.registers.1226[18] [16]),
    .S(\datapath.idinstr_20_bF$buf12 ),
    .Y(_8367_)
);

MUX2X1 _19344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8367_),
    .B(_8366_),
    .S(\datapath.idinstr_21_bF$buf17 ),
    .Y(_8368_)
);

NAND2X1 _19345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf9),
    .B(_8368_),
    .Y(_8369_)
);

MUX2X1 _19346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [16]),
    .B(\datapath.registers.1226[20] [16]),
    .S(\datapath.idinstr_20_bF$buf11 ),
    .Y(_8370_)
);

MUX2X1 _19347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [16]),
    .B(\datapath.registers.1226[22] [16]),
    .S(\datapath.idinstr_20_bF$buf10 ),
    .Y(_8371_)
);

MUX2X1 _19348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8371_),
    .B(_8370_),
    .S(\datapath.idinstr_21_bF$buf16 ),
    .Y(_8372_)
);

NAND2X1 _19349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf4 ),
    .B(_8372_),
    .Y(_8373_)
);

AOI21X1 _19350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8369_),
    .B(_8373_),
    .C(\datapath.idinstr_23_bF$buf0 ),
    .Y(_8374_)
);

OAI21X1 _19351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8374_),
    .B(_8365_),
    .C(\datapath.idinstr_24_bF$buf2 ),
    .Y(_8375_)
);

AOI21X1 _19352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8375_),
    .B(_8351_),
    .C(_7614__bF$buf3),
    .Y(\datapath.registers.regb_data [16])
);

MUX2X1 _19353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [17]),
    .B(\datapath.registers.1226[8] [17]),
    .S(\datapath.idinstr_20_bF$buf9 ),
    .Y(_8376_)
);

MUX2X1 _19354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [17]),
    .B(\datapath.registers.1226[10] [17]),
    .S(\datapath.idinstr_20_bF$buf8 ),
    .Y(_8377_)
);

MUX2X1 _19355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8377_),
    .B(_8376_),
    .S(\datapath.idinstr_21_bF$buf15 ),
    .Y(_8378_)
);

NAND2X1 _19356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf8),
    .B(_8378_),
    .Y(_8379_)
);

AND2X2 _19357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [17]),
    .B(\datapath.idinstr_20_bF$buf7 ),
    .Y(_8380_)
);

INVX1 _19358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [17]),
    .Y(_8381_)
);

OAI21X1 _19359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8381_),
    .B(\datapath.idinstr_20_bF$buf6 ),
    .C(\datapath.idinstr_21_bF$buf14 ),
    .Y(_8382_)
);

NAND2X1 _19360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [17]),
    .B(_7608__bF$buf2),
    .Y(_8383_)
);

AOI21X1 _19361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [17]),
    .B(\datapath.idinstr_20_bF$buf5 ),
    .C(\datapath.idinstr_21_bF$buf13 ),
    .Y(_8384_)
);

AOI21X1 _19362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8384_),
    .B(_8383_),
    .C(_7611__bF$buf7),
    .Y(_8385_)
);

OAI21X1 _19363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8380_),
    .B(_8382_),
    .C(_8385_),
    .Y(_8386_)
);

AOI21X1 _19364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8386_),
    .B(_8379_),
    .C(_7612__bF$buf4),
    .Y(_8387_)
);

MUX2X1 _19365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [17]),
    .B(\datapath.registers.1226[4] [17]),
    .S(\datapath.idinstr_20_bF$buf4 ),
    .Y(_8388_)
);

MUX2X1 _19366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [17]),
    .B(\datapath.registers.1226[6] [17]),
    .S(\datapath.idinstr_20_bF$buf3 ),
    .Y(_8389_)
);

MUX2X1 _19367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8389_),
    .B(_8388_),
    .S(\datapath.idinstr_21_bF$buf12 ),
    .Y(_8390_)
);

NAND2X1 _19368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf3 ),
    .B(_8390_),
    .Y(_8391_)
);

MUX2X1 _19369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [17]),
    .B(\datapath.registers.1226[0] [17]),
    .S(\datapath.idinstr_20_bF$buf2 ),
    .Y(_8392_)
);

MUX2X1 _19370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [17]),
    .B(\datapath.registers.1226[2] [17]),
    .S(\datapath.idinstr_20_bF$buf1 ),
    .Y(_8393_)
);

MUX2X1 _19371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8393_),
    .B(_8392_),
    .S(\datapath.idinstr_21_bF$buf11 ),
    .Y(_8394_)
);

NAND2X1 _19372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf6),
    .B(_8394_),
    .Y(_8395_)
);

AOI21X1 _19373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8391_),
    .B(_8395_),
    .C(\datapath.idinstr_23_bF$buf7 ),
    .Y(_8396_)
);

OAI21X1 _19374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8396_),
    .B(_8387_),
    .C(_7607__bF$buf1),
    .Y(_8397_)
);

INVX1 _19375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [17]),
    .Y(_8398_)
);

AOI21X1 _19376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [17]),
    .B(\datapath.idinstr_22_bF$buf2 ),
    .C(_7608__bF$buf1),
    .Y(_8399_)
);

OAI21X1 _19377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8398_),
    .B(\datapath.idinstr_22_bF$buf1 ),
    .C(_8399_),
    .Y(_8400_)
);

NAND2X1 _19378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [17]),
    .B(_7611__bF$buf5),
    .Y(_8401_)
);

AOI21X1 _19379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [17]),
    .B(\datapath.idinstr_22_bF$buf0 ),
    .C(\datapath.idinstr_20_bF$buf0 ),
    .Y(_8402_)
);

AOI21X1 _19380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8402_),
    .B(_8401_),
    .C(_7610__bF$buf3),
    .Y(_8403_)
);

NAND2X1 _19381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8400_),
    .B(_8403_),
    .Y(_8404_)
);

INVX1 _19382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [17]),
    .Y(_8405_)
);

AOI21X1 _19383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [17]),
    .B(\datapath.idinstr_22_bF$buf43 ),
    .C(_7608__bF$buf0),
    .Y(_8406_)
);

OAI21X1 _19384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8405_),
    .B(\datapath.idinstr_22_bF$buf42 ),
    .C(_8406_),
    .Y(_8407_)
);

AOI21X1 _19385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[28] [17]),
    .B(\datapath.idinstr_22_bF$buf41 ),
    .C(\datapath.idinstr_20_bF$buf55 ),
    .Y(_8408_)
);

OAI21X1 _19386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5736_),
    .B(\datapath.idinstr_22_bF$buf40 ),
    .C(_8408_),
    .Y(_8409_)
);

NAND3X1 _19387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf2),
    .B(_8409_),
    .C(_8407_),
    .Y(_8410_)
);

AOI21X1 _19388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8404_),
    .B(_8410_),
    .C(_7612__bF$buf3),
    .Y(_8411_)
);

MUX2X1 _19389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [17]),
    .B(\datapath.registers.1226[16] [17]),
    .S(\datapath.idinstr_20_bF$buf54 ),
    .Y(_8412_)
);

MUX2X1 _19390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [17]),
    .B(\datapath.registers.1226[18] [17]),
    .S(\datapath.idinstr_20_bF$buf53 ),
    .Y(_8413_)
);

MUX2X1 _19391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8413_),
    .B(_8412_),
    .S(\datapath.idinstr_21_bF$buf10 ),
    .Y(_8414_)
);

NAND2X1 _19392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf4),
    .B(_8414_),
    .Y(_8415_)
);

MUX2X1 _19393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [17]),
    .B(\datapath.registers.1226[20] [17]),
    .S(\datapath.idinstr_20_bF$buf52 ),
    .Y(_8416_)
);

MUX2X1 _19394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [17]),
    .B(\datapath.registers.1226[22] [17]),
    .S(\datapath.idinstr_20_bF$buf51 ),
    .Y(_8417_)
);

MUX2X1 _19395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8417_),
    .B(_8416_),
    .S(\datapath.idinstr_21_bF$buf9 ),
    .Y(_8418_)
);

NAND2X1 _19396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf39 ),
    .B(_8418_),
    .Y(_8419_)
);

AOI21X1 _19397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8415_),
    .B(_8419_),
    .C(\datapath.idinstr_23_bF$buf6 ),
    .Y(_8420_)
);

OAI21X1 _19398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8420_),
    .B(_8411_),
    .C(\datapath.idinstr_24_bF$buf1 ),
    .Y(_8421_)
);

AOI21X1 _19399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8421_),
    .B(_8397_),
    .C(_7614__bF$buf2),
    .Y(\datapath.registers.regb_data [17])
);

MUX2X1 _19400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [18]),
    .B(\datapath.registers.1226[24] [18]),
    .S(\datapath.idinstr_20_bF$buf50 ),
    .Y(_8422_)
);

MUX2X1 _19401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [18]),
    .B(\datapath.registers.1226[26] [18]),
    .S(\datapath.idinstr_20_bF$buf49 ),
    .Y(_8423_)
);

MUX2X1 _19402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8423_),
    .B(_8422_),
    .S(\datapath.idinstr_21_bF$buf8 ),
    .Y(_8424_)
);

NAND2X1 _19403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf3),
    .B(_8424_),
    .Y(_8425_)
);

MUX2X1 _19404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [18]),
    .B(\datapath.registers.1226[28] [18]),
    .S(\datapath.idinstr_20_bF$buf48 ),
    .Y(_8426_)
);

MUX2X1 _19405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [18]),
    .B(\datapath.registers.1226[30] [18]),
    .S(\datapath.idinstr_20_bF$buf47 ),
    .Y(_8427_)
);

MUX2X1 _19406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8427_),
    .B(_8426_),
    .S(\datapath.idinstr_21_bF$buf7 ),
    .Y(_8428_)
);

NAND2X1 _19407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf38 ),
    .B(_8428_),
    .Y(_8429_)
);

AOI21X1 _19408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8425_),
    .B(_8429_),
    .C(_7612__bF$buf2),
    .Y(_8430_)
);

MUX2X1 _19409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [18]),
    .B(\datapath.registers.1226[16] [18]),
    .S(\datapath.idinstr_21_bF$buf6 ),
    .Y(_8431_)
);

NAND2X1 _19410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf10),
    .B(_8431_),
    .Y(_8432_)
);

MUX2X1 _19411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [18]),
    .B(\datapath.registers.1226[17] [18]),
    .S(\datapath.idinstr_21_bF$buf5 ),
    .Y(_8433_)
);

AOI21X1 _19412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf46 ),
    .B(_8433_),
    .C(\datapath.idinstr_22_bF$buf37 ),
    .Y(_8434_)
);

NAND2X1 _19413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8432_),
    .B(_8434_),
    .Y(_8435_)
);

MUX2X1 _19414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [18]),
    .B(\datapath.registers.1226[20] [18]),
    .S(\datapath.idinstr_21_bF$buf4 ),
    .Y(_8436_)
);

NAND2X1 _19415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf9),
    .B(_8436_),
    .Y(_8437_)
);

MUX2X1 _19416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [18]),
    .B(\datapath.registers.1226[21] [18]),
    .S(\datapath.idinstr_21_bF$buf3 ),
    .Y(_8438_)
);

AOI21X1 _19417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf45 ),
    .B(_8438_),
    .C(_7611__bF$buf2),
    .Y(_8439_)
);

NAND2X1 _19418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8437_),
    .B(_8439_),
    .Y(_8440_)
);

AOI21X1 _19419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8435_),
    .B(_8440_),
    .C(\datapath.idinstr_23_bF$buf5 ),
    .Y(_8441_)
);

OAI21X1 _19420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8430_),
    .B(_8441_),
    .C(\datapath.idinstr_24_bF$buf0 ),
    .Y(_8442_)
);

INVX1 _19421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [18]),
    .Y(_8443_)
);

AOI21X1 _19422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [18]),
    .B(\datapath.idinstr_22_bF$buf36 ),
    .C(_7608__bF$buf8),
    .Y(_8444_)
);

OAI21X1 _19423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8443_),
    .B(\datapath.idinstr_22_bF$buf35 ),
    .C(_8444_),
    .Y(_8445_)
);

INVX1 _19424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [18]),
    .Y(_8446_)
);

AOI21X1 _19425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [18]),
    .B(\datapath.idinstr_22_bF$buf34 ),
    .C(\datapath.idinstr_20_bF$buf44 ),
    .Y(_8447_)
);

OAI21X1 _19426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8446_),
    .B(\datapath.idinstr_22_bF$buf33 ),
    .C(_8447_),
    .Y(_8448_)
);

NAND3X1 _19427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf1),
    .B(_8448_),
    .C(_8445_),
    .Y(_8449_)
);

INVX1 _19428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [18]),
    .Y(_8450_)
);

AOI21X1 _19429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [18]),
    .B(\datapath.idinstr_22_bF$buf32 ),
    .C(_7608__bF$buf7),
    .Y(_8451_)
);

OAI21X1 _19430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8450_),
    .B(\datapath.idinstr_22_bF$buf31 ),
    .C(_8451_),
    .Y(_8452_)
);

INVX1 _19431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[10] [18]),
    .Y(_8453_)
);

AOI21X1 _19432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [18]),
    .B(\datapath.idinstr_22_bF$buf30 ),
    .C(\datapath.idinstr_20_bF$buf43 ),
    .Y(_8454_)
);

OAI21X1 _19433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8453_),
    .B(\datapath.idinstr_22_bF$buf29 ),
    .C(_8454_),
    .Y(_8455_)
);

NAND3X1 _19434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf2 ),
    .B(_8455_),
    .C(_8452_),
    .Y(_8456_)
);

AOI21X1 _19435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8449_),
    .B(_8456_),
    .C(_7612__bF$buf1),
    .Y(_8457_)
);

MUX2X1 _19436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [18]),
    .B(\datapath.registers.1226[0] [18]),
    .S(\datapath.idinstr_20_bF$buf42 ),
    .Y(_8458_)
);

MUX2X1 _19437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [18]),
    .B(\datapath.registers.1226[2] [18]),
    .S(\datapath.idinstr_20_bF$buf41 ),
    .Y(_8459_)
);

MUX2X1 _19438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8459_),
    .B(_8458_),
    .S(\datapath.idinstr_21_bF$buf1 ),
    .Y(_8460_)
);

NAND2X1 _19439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf1),
    .B(_8460_),
    .Y(_8461_)
);

MUX2X1 _19440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [18]),
    .B(\datapath.registers.1226[4] [18]),
    .S(\datapath.idinstr_20_bF$buf40 ),
    .Y(_8462_)
);

MUX2X1 _19441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [18]),
    .B(\datapath.registers.1226[6] [18]),
    .S(\datapath.idinstr_20_bF$buf39 ),
    .Y(_8463_)
);

MUX2X1 _19442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8463_),
    .B(_8462_),
    .S(\datapath.idinstr_21_bF$buf0 ),
    .Y(_8464_)
);

NAND2X1 _19443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf28 ),
    .B(_8464_),
    .Y(_8465_)
);

AOI21X1 _19444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8461_),
    .B(_8465_),
    .C(\datapath.idinstr_23_bF$buf4 ),
    .Y(_8466_)
);

OAI21X1 _19445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8466_),
    .B(_8457_),
    .C(_7607__bF$buf0),
    .Y(_8467_)
);

AOI21X1 _19446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8442_),
    .B(_8467_),
    .C(_7614__bF$buf1),
    .Y(\datapath.registers.regb_data [18])
);

MUX2X1 _19447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [19]),
    .B(\datapath.registers.1226[24] [19]),
    .S(\datapath.idinstr_20_bF$buf38 ),
    .Y(_8468_)
);

MUX2X1 _19448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [19]),
    .B(\datapath.registers.1226[26] [19]),
    .S(\datapath.idinstr_20_bF$buf37 ),
    .Y(_8469_)
);

MUX2X1 _19449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8469_),
    .B(_8468_),
    .S(\datapath.idinstr_21_bF$buf44 ),
    .Y(_8470_)
);

NAND2X1 _19450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf0),
    .B(_8470_),
    .Y(_8471_)
);

MUX2X1 _19451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [19]),
    .B(\datapath.registers.1226[28] [19]),
    .S(\datapath.idinstr_20_bF$buf36 ),
    .Y(_8472_)
);

MUX2X1 _19452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [19]),
    .B(\datapath.registers.1226[30] [19]),
    .S(\datapath.idinstr_20_bF$buf35 ),
    .Y(_8473_)
);

MUX2X1 _19453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8473_),
    .B(_8472_),
    .S(\datapath.idinstr_21_bF$buf43 ),
    .Y(_8474_)
);

NAND2X1 _19454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf27 ),
    .B(_8474_),
    .Y(_8475_)
);

AOI21X1 _19455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8471_),
    .B(_8475_),
    .C(_7612__bF$buf0),
    .Y(_8476_)
);

MUX2X1 _19456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [19]),
    .B(\datapath.registers.1226[16] [19]),
    .S(\datapath.idinstr_21_bF$buf42 ),
    .Y(_8477_)
);

NAND2X1 _19457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf6),
    .B(_8477_),
    .Y(_8478_)
);

MUX2X1 _19458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [19]),
    .B(\datapath.registers.1226[17] [19]),
    .S(\datapath.idinstr_21_bF$buf41 ),
    .Y(_8479_)
);

AOI21X1 _19459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf34 ),
    .B(_8479_),
    .C(\datapath.idinstr_22_bF$buf26 ),
    .Y(_8480_)
);

NAND2X1 _19460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8478_),
    .B(_8480_),
    .Y(_8481_)
);

MUX2X1 _19461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [19]),
    .B(\datapath.registers.1226[20] [19]),
    .S(\datapath.idinstr_21_bF$buf40 ),
    .Y(_8482_)
);

NAND2X1 _19462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf5),
    .B(_8482_),
    .Y(_8483_)
);

MUX2X1 _19463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [19]),
    .B(\datapath.registers.1226[21] [19]),
    .S(\datapath.idinstr_21_bF$buf39 ),
    .Y(_8484_)
);

AOI21X1 _19464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf33 ),
    .B(_8484_),
    .C(_7611__bF$buf10),
    .Y(_8485_)
);

NAND2X1 _19465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8483_),
    .B(_8485_),
    .Y(_8486_)
);

AOI21X1 _19466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8481_),
    .B(_8486_),
    .C(\datapath.idinstr_23_bF$buf3 ),
    .Y(_8487_)
);

OAI21X1 _19467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8476_),
    .B(_8487_),
    .C(\datapath.idinstr_24_bF$buf5 ),
    .Y(_8488_)
);

MUX2X1 _19468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [19]),
    .B(\datapath.registers.1226[8] [19]),
    .S(\datapath.idinstr_20_bF$buf32 ),
    .Y(_8489_)
);

MUX2X1 _19469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [19]),
    .B(\datapath.registers.1226[10] [19]),
    .S(\datapath.idinstr_20_bF$buf31 ),
    .Y(_8490_)
);

MUX2X1 _19470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8490_),
    .B(_8489_),
    .S(\datapath.idinstr_21_bF$buf38 ),
    .Y(_8491_)
);

NAND2X1 _19471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf9),
    .B(_8491_),
    .Y(_8492_)
);

MUX2X1 _19472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [19]),
    .B(\datapath.registers.1226[12] [19]),
    .S(\datapath.idinstr_20_bF$buf30 ),
    .Y(_8493_)
);

MUX2X1 _19473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [19]),
    .B(\datapath.registers.1226[14] [19]),
    .S(\datapath.idinstr_20_bF$buf29 ),
    .Y(_8494_)
);

MUX2X1 _19474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8494_),
    .B(_8493_),
    .S(\datapath.idinstr_21_bF$buf37 ),
    .Y(_8495_)
);

NAND2X1 _19475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf25 ),
    .B(_8495_),
    .Y(_8496_)
);

AOI21X1 _19476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8492_),
    .B(_8496_),
    .C(_7612__bF$buf7),
    .Y(_8497_)
);

AOI21X1 _19477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [19]),
    .B(\datapath.idinstr_22_bF$buf24 ),
    .C(_7608__bF$buf4),
    .Y(_8498_)
);

OAI21X1 _19478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7045_),
    .B(\datapath.idinstr_22_bF$buf23 ),
    .C(_8498_),
    .Y(_8499_)
);

AOI21X1 _19479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [19]),
    .B(\datapath.idinstr_22_bF$buf22 ),
    .C(\datapath.idinstr_20_bF$buf28 ),
    .Y(_8500_)
);

OAI21X1 _19480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7048_),
    .B(\datapath.idinstr_22_bF$buf21 ),
    .C(_8500_),
    .Y(_8501_)
);

NAND3X1 _19481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf0),
    .B(_8501_),
    .C(_8499_),
    .Y(_8502_)
);

AOI21X1 _19482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [19]),
    .B(\datapath.idinstr_22_bF$buf20 ),
    .C(_7608__bF$buf3),
    .Y(_8503_)
);

OAI21X1 _19483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7052_),
    .B(\datapath.idinstr_22_bF$buf19 ),
    .C(_8503_),
    .Y(_8504_)
);

AOI21X1 _19484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[6] [19]),
    .B(\datapath.idinstr_22_bF$buf18 ),
    .C(\datapath.idinstr_20_bF$buf27 ),
    .Y(_8505_)
);

OAI21X1 _19485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7055_),
    .B(\datapath.idinstr_22_bF$buf17 ),
    .C(_8505_),
    .Y(_8506_)
);

NAND3X1 _19486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf36 ),
    .B(_8506_),
    .C(_8504_),
    .Y(_8507_)
);

AOI21X1 _19487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8502_),
    .B(_8507_),
    .C(\datapath.idinstr_23_bF$buf2 ),
    .Y(_8508_)
);

OAI21X1 _19488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8497_),
    .B(_8508_),
    .C(_7607__bF$buf4),
    .Y(_8509_)
);

AOI21X1 _19489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8488_),
    .B(_8509_),
    .C(_7614__bF$buf0),
    .Y(\datapath.registers.regb_data [19])
);

MUX2X1 _19490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [20]),
    .B(\datapath.registers.1226[24] [20]),
    .S(\datapath.idinstr_20_bF$buf26 ),
    .Y(_8510_)
);

MUX2X1 _19491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [20]),
    .B(\datapath.registers.1226[26] [20]),
    .S(\datapath.idinstr_20_bF$buf25 ),
    .Y(_8511_)
);

MUX2X1 _19492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8511_),
    .B(_8510_),
    .S(\datapath.idinstr_21_bF$buf35 ),
    .Y(_8512_)
);

NAND2X1 _19493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf8),
    .B(_8512_),
    .Y(_8513_)
);

MUX2X1 _19494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [20]),
    .B(\datapath.registers.1226[28] [20]),
    .S(\datapath.idinstr_20_bF$buf24 ),
    .Y(_8514_)
);

MUX2X1 _19495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [20]),
    .B(\datapath.registers.1226[30] [20]),
    .S(\datapath.idinstr_20_bF$buf23 ),
    .Y(_8515_)
);

MUX2X1 _19496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8515_),
    .B(_8514_),
    .S(\datapath.idinstr_21_bF$buf34 ),
    .Y(_8516_)
);

NAND2X1 _19497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf16 ),
    .B(_8516_),
    .Y(_8517_)
);

AOI21X1 _19498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8513_),
    .B(_8517_),
    .C(_7612__bF$buf6),
    .Y(_8518_)
);

MUX2X1 _19499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [20]),
    .B(\datapath.registers.1226[16] [20]),
    .S(\datapath.idinstr_21_bF$buf33 ),
    .Y(_8519_)
);

NAND2X1 _19500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf2),
    .B(_8519_),
    .Y(_8520_)
);

MUX2X1 _19501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [20]),
    .B(\datapath.registers.1226[17] [20]),
    .S(\datapath.idinstr_21_bF$buf32 ),
    .Y(_8521_)
);

AOI21X1 _19502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf22 ),
    .B(_8521_),
    .C(\datapath.idinstr_22_bF$buf15 ),
    .Y(_8522_)
);

NAND2X1 _19503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8520_),
    .B(_8522_),
    .Y(_8523_)
);

MUX2X1 _19504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [20]),
    .B(\datapath.registers.1226[20] [20]),
    .S(\datapath.idinstr_21_bF$buf31 ),
    .Y(_8524_)
);

NAND2X1 _19505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf1),
    .B(_8524_),
    .Y(_8525_)
);

MUX2X1 _19506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [20]),
    .B(\datapath.registers.1226[21] [20]),
    .S(\datapath.idinstr_21_bF$buf30 ),
    .Y(_8526_)
);

AOI21X1 _19507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf21 ),
    .B(_8526_),
    .C(_7611__bF$buf7),
    .Y(_8527_)
);

NAND2X1 _19508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8525_),
    .B(_8527_),
    .Y(_8528_)
);

AOI21X1 _19509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8523_),
    .B(_8528_),
    .C(\datapath.idinstr_23_bF$buf1 ),
    .Y(_8529_)
);

OAI21X1 _19510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8518_),
    .B(_8529_),
    .C(\datapath.idinstr_24_bF$buf4 ),
    .Y(_8530_)
);

MUX2X1 _19511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [20]),
    .B(\datapath.registers.1226[8] [20]),
    .S(\datapath.idinstr_20_bF$buf20 ),
    .Y(_8531_)
);

MUX2X1 _19512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [20]),
    .B(\datapath.registers.1226[10] [20]),
    .S(\datapath.idinstr_20_bF$buf19 ),
    .Y(_8532_)
);

MUX2X1 _19513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8532_),
    .B(_8531_),
    .S(\datapath.idinstr_21_bF$buf29 ),
    .Y(_8533_)
);

NAND2X1 _19514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf6),
    .B(_8533_),
    .Y(_8534_)
);

NOR2X1 _19515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7065_),
    .B(_7608__bF$buf0),
    .Y(_8535_)
);

OAI21X1 _19516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7067_),
    .B(\datapath.idinstr_20_bF$buf18 ),
    .C(\datapath.idinstr_21_bF$buf28 ),
    .Y(_8536_)
);

NAND2X1 _19517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [20]),
    .B(_7608__bF$buf10),
    .Y(_8537_)
);

AOI21X1 _19518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [20]),
    .B(\datapath.idinstr_20_bF$buf17 ),
    .C(\datapath.idinstr_21_bF$buf27 ),
    .Y(_8538_)
);

AOI21X1 _19519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8538_),
    .B(_8537_),
    .C(_7611__bF$buf5),
    .Y(_8539_)
);

OAI21X1 _19520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8535_),
    .B(_8536_),
    .C(_8539_),
    .Y(_8540_)
);

AOI21X1 _19521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8540_),
    .B(_8534_),
    .C(_7612__bF$buf5),
    .Y(_8541_)
);

MUX2X1 _19522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [20]),
    .B(\datapath.registers.1226[4] [20]),
    .S(\datapath.idinstr_20_bF$buf16 ),
    .Y(_8542_)
);

MUX2X1 _19523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [20]),
    .B(\datapath.registers.1226[6] [20]),
    .S(\datapath.idinstr_20_bF$buf15 ),
    .Y(_8543_)
);

MUX2X1 _19524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8543_),
    .B(_8542_),
    .S(\datapath.idinstr_21_bF$buf26 ),
    .Y(_8544_)
);

NAND2X1 _19525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf14 ),
    .B(_8544_),
    .Y(_8545_)
);

MUX2X1 _19526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [20]),
    .B(\datapath.registers.1226[0] [20]),
    .S(\datapath.idinstr_20_bF$buf14 ),
    .Y(_8546_)
);

MUX2X1 _19527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [20]),
    .B(\datapath.registers.1226[2] [20]),
    .S(\datapath.idinstr_20_bF$buf13 ),
    .Y(_8547_)
);

MUX2X1 _19528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8547_),
    .B(_8546_),
    .S(\datapath.idinstr_21_bF$buf25 ),
    .Y(_8548_)
);

NAND2X1 _19529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf4),
    .B(_8548_),
    .Y(_8549_)
);

AOI21X1 _19530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8545_),
    .B(_8549_),
    .C(\datapath.idinstr_23_bF$buf0 ),
    .Y(_8550_)
);

OAI21X1 _19531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8550_),
    .B(_8541_),
    .C(_7607__bF$buf3),
    .Y(_8551_)
);

AOI21X1 _19532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8530_),
    .B(_8551_),
    .C(_7614__bF$buf4),
    .Y(\datapath.registers.regb_data [20])
);

MUX2X1 _19533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [21]),
    .B(\datapath.registers.1226[8] [21]),
    .S(\datapath.idinstr_20_bF$buf12 ),
    .Y(_8552_)
);

MUX2X1 _19534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [21]),
    .B(\datapath.registers.1226[10] [21]),
    .S(\datapath.idinstr_20_bF$buf11 ),
    .Y(_8553_)
);

MUX2X1 _19535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8553_),
    .B(_8552_),
    .S(\datapath.idinstr_21_bF$buf24 ),
    .Y(_8554_)
);

NAND2X1 _19536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf3),
    .B(_8554_),
    .Y(_8555_)
);

NOR2X1 _19537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7112_),
    .B(_7608__bF$buf9),
    .Y(_8556_)
);

OAI21X1 _19538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7114_),
    .B(\datapath.idinstr_20_bF$buf10 ),
    .C(\datapath.idinstr_21_bF$buf23 ),
    .Y(_8557_)
);

NAND2X1 _19539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [21]),
    .B(_7608__bF$buf8),
    .Y(_8558_)
);

AOI21X1 _19540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [21]),
    .B(\datapath.idinstr_20_bF$buf9 ),
    .C(\datapath.idinstr_21_bF$buf22 ),
    .Y(_8559_)
);

AOI21X1 _19541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8559_),
    .B(_8558_),
    .C(_7611__bF$buf2),
    .Y(_8560_)
);

OAI21X1 _19542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8556_),
    .B(_8557_),
    .C(_8560_),
    .Y(_8561_)
);

AOI21X1 _19543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8561_),
    .B(_8555_),
    .C(_7612__bF$buf4),
    .Y(_8562_)
);

MUX2X1 _19544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [21]),
    .B(\datapath.registers.1226[4] [21]),
    .S(\datapath.idinstr_20_bF$buf8 ),
    .Y(_8563_)
);

MUX2X1 _19545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [21]),
    .B(\datapath.registers.1226[6] [21]),
    .S(\datapath.idinstr_20_bF$buf7 ),
    .Y(_8564_)
);

MUX2X1 _19546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8564_),
    .B(_8563_),
    .S(\datapath.idinstr_21_bF$buf21 ),
    .Y(_8565_)
);

NAND2X1 _19547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf13 ),
    .B(_8565_),
    .Y(_8566_)
);

MUX2X1 _19548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [21]),
    .B(\datapath.registers.1226[0] [21]),
    .S(\datapath.idinstr_20_bF$buf6 ),
    .Y(_8567_)
);

MUX2X1 _19549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [21]),
    .B(\datapath.registers.1226[2] [21]),
    .S(\datapath.idinstr_20_bF$buf5 ),
    .Y(_8568_)
);

MUX2X1 _19550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8568_),
    .B(_8567_),
    .S(\datapath.idinstr_21_bF$buf20 ),
    .Y(_8569_)
);

NAND2X1 _19551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf1),
    .B(_8569_),
    .Y(_8570_)
);

AOI21X1 _19552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8566_),
    .B(_8570_),
    .C(\datapath.idinstr_23_bF$buf7 ),
    .Y(_8571_)
);

OAI21X1 _19553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8571_),
    .B(_8562_),
    .C(_7607__bF$buf2),
    .Y(_8572_)
);

INVX1 _19554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [21]),
    .Y(_8573_)
);

AOI21X1 _19555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [21]),
    .B(\datapath.idinstr_22_bF$buf12 ),
    .C(_7608__bF$buf7),
    .Y(_8574_)
);

OAI21X1 _19556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8573_),
    .B(\datapath.idinstr_22_bF$buf11 ),
    .C(_8574_),
    .Y(_8575_)
);

NAND2X1 _19557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [21]),
    .B(_7611__bF$buf0),
    .Y(_8576_)
);

AOI21X1 _19558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [21]),
    .B(\datapath.idinstr_22_bF$buf10 ),
    .C(\datapath.idinstr_20_bF$buf4 ),
    .Y(_8577_)
);

AOI21X1 _19559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8577_),
    .B(_8576_),
    .C(_7610__bF$buf4),
    .Y(_8578_)
);

NAND2X1 _19560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8575_),
    .B(_8578_),
    .Y(_8579_)
);

INVX1 _19561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [21]),
    .Y(_8580_)
);

AOI21X1 _19562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [21]),
    .B(\datapath.idinstr_22_bF$buf9 ),
    .C(_7608__bF$buf6),
    .Y(_8581_)
);

OAI21X1 _19563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8580_),
    .B(\datapath.idinstr_22_bF$buf8 ),
    .C(_8581_),
    .Y(_8582_)
);

AOI21X1 _19564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[28] [21]),
    .B(\datapath.idinstr_22_bF$buf7 ),
    .C(\datapath.idinstr_20_bF$buf3 ),
    .Y(_8583_)
);

OAI21X1 _19565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5742_),
    .B(\datapath.idinstr_22_bF$buf6 ),
    .C(_8583_),
    .Y(_8584_)
);

NAND3X1 _19566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf3),
    .B(_8584_),
    .C(_8582_),
    .Y(_8585_)
);

AOI21X1 _19567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8579_),
    .B(_8585_),
    .C(_7612__bF$buf3),
    .Y(_8586_)
);

MUX2X1 _19568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [21]),
    .B(\datapath.registers.1226[16] [21]),
    .S(\datapath.idinstr_20_bF$buf2 ),
    .Y(_8587_)
);

MUX2X1 _19569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [21]),
    .B(\datapath.registers.1226[18] [21]),
    .S(\datapath.idinstr_20_bF$buf1 ),
    .Y(_8588_)
);

MUX2X1 _19570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8588_),
    .B(_8587_),
    .S(\datapath.idinstr_21_bF$buf19 ),
    .Y(_8589_)
);

NAND2X1 _19571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf10),
    .B(_8589_),
    .Y(_8590_)
);

MUX2X1 _19572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [21]),
    .B(\datapath.registers.1226[20] [21]),
    .S(\datapath.idinstr_20_bF$buf0 ),
    .Y(_8591_)
);

MUX2X1 _19573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [21]),
    .B(\datapath.registers.1226[22] [21]),
    .S(\datapath.idinstr_20_bF$buf55 ),
    .Y(_8592_)
);

MUX2X1 _19574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8592_),
    .B(_8591_),
    .S(\datapath.idinstr_21_bF$buf18 ),
    .Y(_8593_)
);

NAND2X1 _19575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf5 ),
    .B(_8593_),
    .Y(_8594_)
);

AOI21X1 _19576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8590_),
    .B(_8594_),
    .C(\datapath.idinstr_23_bF$buf6 ),
    .Y(_8595_)
);

OAI21X1 _19577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8595_),
    .B(_8586_),
    .C(\datapath.idinstr_24_bF$buf3 ),
    .Y(_8596_)
);

AOI21X1 _19578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8596_),
    .B(_8572_),
    .C(_7614__bF$buf3),
    .Y(\datapath.registers.regb_data [21])
);

MUX2X1 _19579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [22]),
    .B(\datapath.registers.1226[8] [22]),
    .S(\datapath.idinstr_20_bF$buf54 ),
    .Y(_8597_)
);

MUX2X1 _19580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [22]),
    .B(\datapath.registers.1226[10] [22]),
    .S(\datapath.idinstr_20_bF$buf53 ),
    .Y(_8598_)
);

MUX2X1 _19581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8598_),
    .B(_8597_),
    .S(\datapath.idinstr_21_bF$buf17 ),
    .Y(_8599_)
);

NAND2X1 _19582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf9),
    .B(_8599_),
    .Y(_8600_)
);

NOR2X1 _19583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7180_),
    .B(_7608__bF$buf5),
    .Y(_8601_)
);

OAI21X1 _19584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7182_),
    .B(\datapath.idinstr_20_bF$buf52 ),
    .C(\datapath.idinstr_21_bF$buf16 ),
    .Y(_8602_)
);

NAND2X1 _19585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [22]),
    .B(_7608__bF$buf4),
    .Y(_8603_)
);

AOI21X1 _19586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [22]),
    .B(\datapath.idinstr_20_bF$buf51 ),
    .C(\datapath.idinstr_21_bF$buf15 ),
    .Y(_8604_)
);

AOI21X1 _19587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8604_),
    .B(_8603_),
    .C(_7611__bF$buf8),
    .Y(_8605_)
);

OAI21X1 _19588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8601_),
    .B(_8602_),
    .C(_8605_),
    .Y(_8606_)
);

AOI21X1 _19589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8606_),
    .B(_8600_),
    .C(_7612__bF$buf2),
    .Y(_8607_)
);

MUX2X1 _19590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [22]),
    .B(\datapath.registers.1226[4] [22]),
    .S(\datapath.idinstr_20_bF$buf50 ),
    .Y(_8608_)
);

MUX2X1 _19591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [22]),
    .B(\datapath.registers.1226[6] [22]),
    .S(\datapath.idinstr_20_bF$buf49 ),
    .Y(_8609_)
);

MUX2X1 _19592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8609_),
    .B(_8608_),
    .S(\datapath.idinstr_21_bF$buf14 ),
    .Y(_8610_)
);

NAND2X1 _19593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf4 ),
    .B(_8610_),
    .Y(_8611_)
);

MUX2X1 _19594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [22]),
    .B(\datapath.registers.1226[0] [22]),
    .S(\datapath.idinstr_20_bF$buf48 ),
    .Y(_8612_)
);

MUX2X1 _19595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [22]),
    .B(\datapath.registers.1226[2] [22]),
    .S(\datapath.idinstr_20_bF$buf47 ),
    .Y(_8613_)
);

MUX2X1 _19596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8613_),
    .B(_8612_),
    .S(\datapath.idinstr_21_bF$buf13 ),
    .Y(_8614_)
);

NAND2X1 _19597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf7),
    .B(_8614_),
    .Y(_8615_)
);

AOI21X1 _19598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8611_),
    .B(_8615_),
    .C(\datapath.idinstr_23_bF$buf5 ),
    .Y(_8616_)
);

OAI21X1 _19599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8616_),
    .B(_8607_),
    .C(_7607__bF$buf1),
    .Y(_8617_)
);

INVX1 _19600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [22]),
    .Y(_8618_)
);

AOI21X1 _19601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [22]),
    .B(\datapath.idinstr_22_bF$buf3 ),
    .C(_7608__bF$buf3),
    .Y(_8619_)
);

OAI21X1 _19602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8618_),
    .B(\datapath.idinstr_22_bF$buf2 ),
    .C(_8619_),
    .Y(_8620_)
);

NAND2X1 _19603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [22]),
    .B(_7611__bF$buf6),
    .Y(_8621_)
);

AOI21X1 _19604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [22]),
    .B(\datapath.idinstr_22_bF$buf1 ),
    .C(\datapath.idinstr_20_bF$buf46 ),
    .Y(_8622_)
);

AOI21X1 _19605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8622_),
    .B(_8621_),
    .C(_7610__bF$buf2),
    .Y(_8623_)
);

NAND2X1 _19606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8620_),
    .B(_8623_),
    .Y(_8624_)
);

INVX1 _19607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [22]),
    .Y(_8625_)
);

AOI21X1 _19608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [22]),
    .B(\datapath.idinstr_22_bF$buf0 ),
    .C(_7608__bF$buf2),
    .Y(_8626_)
);

OAI21X1 _19609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8625_),
    .B(\datapath.idinstr_22_bF$buf43 ),
    .C(_8626_),
    .Y(_8627_)
);

AOI21X1 _19610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[20] [22]),
    .B(\datapath.idinstr_22_bF$buf42 ),
    .C(\datapath.idinstr_20_bF$buf45 ),
    .Y(_8628_)
);

OAI21X1 _19611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6026_),
    .B(\datapath.idinstr_22_bF$buf41 ),
    .C(_8628_),
    .Y(_8629_)
);

NAND3X1 _19612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf1),
    .B(_8629_),
    .C(_8627_),
    .Y(_8630_)
);

AOI21X1 _19613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8624_),
    .B(_8630_),
    .C(\datapath.idinstr_23_bF$buf4 ),
    .Y(_8631_)
);

MUX2X1 _19614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [22]),
    .B(\datapath.registers.1226[29] [22]),
    .S(\datapath.idinstr_21_bF$buf12 ),
    .Y(_8632_)
);

MUX2X1 _19615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [22]),
    .B(\datapath.registers.1226[28] [22]),
    .S(\datapath.idinstr_21_bF$buf11 ),
    .Y(_8633_)
);

MUX2X1 _19616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8633_),
    .B(_8632_),
    .S(_7608__bF$buf1),
    .Y(_8634_)
);

NAND2X1 _19617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf40 ),
    .B(_8634_),
    .Y(_8635_)
);

MUX2X1 _19618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [22]),
    .B(\datapath.registers.1226[25] [22]),
    .S(\datapath.idinstr_21_bF$buf10 ),
    .Y(_8636_)
);

MUX2X1 _19619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [22]),
    .B(\datapath.registers.1226[24] [22]),
    .S(\datapath.idinstr_21_bF$buf9 ),
    .Y(_8637_)
);

MUX2X1 _19620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8637_),
    .B(_8636_),
    .S(_7608__bF$buf0),
    .Y(_8638_)
);

NAND2X1 _19621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf5),
    .B(_8638_),
    .Y(_8639_)
);

AOI21X1 _19622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8635_),
    .B(_8639_),
    .C(_7612__bF$buf1),
    .Y(_8640_)
);

OAI21X1 _19623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8640_),
    .B(_8631_),
    .C(\datapath.idinstr_24_bF$buf2 ),
    .Y(_8641_)
);

AOI21X1 _19624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8641_),
    .B(_8617_),
    .C(_7614__bF$buf2),
    .Y(\datapath.registers.regb_data [22])
);

MUX2X1 _19625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [23]),
    .B(\datapath.registers.1226[24] [23]),
    .S(\datapath.idinstr_20_bF$buf44 ),
    .Y(_8642_)
);

MUX2X1 _19626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [23]),
    .B(\datapath.registers.1226[26] [23]),
    .S(\datapath.idinstr_20_bF$buf43 ),
    .Y(_8643_)
);

MUX2X1 _19627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8643_),
    .B(_8642_),
    .S(\datapath.idinstr_21_bF$buf8 ),
    .Y(_8644_)
);

NAND2X1 _19628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf4),
    .B(_8644_),
    .Y(_8645_)
);

MUX2X1 _19629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [23]),
    .B(\datapath.registers.1226[28] [23]),
    .S(\datapath.idinstr_20_bF$buf42 ),
    .Y(_8646_)
);

MUX2X1 _19630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [23]),
    .B(\datapath.registers.1226[30] [23]),
    .S(\datapath.idinstr_20_bF$buf41 ),
    .Y(_8647_)
);

MUX2X1 _19631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8647_),
    .B(_8646_),
    .S(\datapath.idinstr_21_bF$buf7 ),
    .Y(_8648_)
);

NAND2X1 _19632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf39 ),
    .B(_8648_),
    .Y(_8649_)
);

AOI21X1 _19633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8645_),
    .B(_8649_),
    .C(_7612__bF$buf0),
    .Y(_8650_)
);

MUX2X1 _19634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [23]),
    .B(\datapath.registers.1226[16] [23]),
    .S(\datapath.idinstr_21_bF$buf6 ),
    .Y(_8651_)
);

NAND2X1 _19635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf10),
    .B(_8651_),
    .Y(_8652_)
);

MUX2X1 _19636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [23]),
    .B(\datapath.registers.1226[17] [23]),
    .S(\datapath.idinstr_21_bF$buf5 ),
    .Y(_8653_)
);

AOI21X1 _19637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf40 ),
    .B(_8653_),
    .C(\datapath.idinstr_22_bF$buf38 ),
    .Y(_8654_)
);

NAND2X1 _19638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8652_),
    .B(_8654_),
    .Y(_8655_)
);

MUX2X1 _19639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [23]),
    .B(\datapath.registers.1226[20] [23]),
    .S(\datapath.idinstr_21_bF$buf4 ),
    .Y(_8656_)
);

NAND2X1 _19640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf9),
    .B(_8656_),
    .Y(_8657_)
);

MUX2X1 _19641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [23]),
    .B(\datapath.registers.1226[21] [23]),
    .S(\datapath.idinstr_21_bF$buf3 ),
    .Y(_8658_)
);

AOI21X1 _19642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf39 ),
    .B(_8658_),
    .C(_7611__bF$buf3),
    .Y(_8659_)
);

NAND2X1 _19643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8657_),
    .B(_8659_),
    .Y(_8660_)
);

AOI21X1 _19644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8655_),
    .B(_8660_),
    .C(\datapath.idinstr_23_bF$buf3 ),
    .Y(_8661_)
);

OAI21X1 _19645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8650_),
    .B(_8661_),
    .C(\datapath.idinstr_24_bF$buf1 ),
    .Y(_8662_)
);

MUX2X1 _19646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [23]),
    .B(\datapath.registers.1226[8] [23]),
    .S(\datapath.idinstr_20_bF$buf38 ),
    .Y(_8663_)
);

MUX2X1 _19647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [23]),
    .B(\datapath.registers.1226[10] [23]),
    .S(\datapath.idinstr_20_bF$buf37 ),
    .Y(_8664_)
);

MUX2X1 _19648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8664_),
    .B(_8663_),
    .S(\datapath.idinstr_21_bF$buf2 ),
    .Y(_8665_)
);

NAND2X1 _19649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf2),
    .B(_8665_),
    .Y(_8666_)
);

NOR2X1 _19650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7224_),
    .B(_7608__bF$buf8),
    .Y(_8667_)
);

OAI21X1 _19651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7226_),
    .B(\datapath.idinstr_20_bF$buf36 ),
    .C(\datapath.idinstr_21_bF$buf1 ),
    .Y(_8668_)
);

NAND2X1 _19652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [23]),
    .B(_7608__bF$buf7),
    .Y(_8669_)
);

AOI21X1 _19653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [23]),
    .B(\datapath.idinstr_20_bF$buf35 ),
    .C(\datapath.idinstr_21_bF$buf0 ),
    .Y(_8670_)
);

AOI21X1 _19654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8670_),
    .B(_8669_),
    .C(_7611__bF$buf1),
    .Y(_8671_)
);

OAI21X1 _19655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8667_),
    .B(_8668_),
    .C(_8671_),
    .Y(_8672_)
);

AOI21X1 _19656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8672_),
    .B(_8666_),
    .C(_7612__bF$buf7),
    .Y(_8673_)
);

MUX2X1 _19657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [23]),
    .B(\datapath.registers.1226[4] [23]),
    .S(\datapath.idinstr_20_bF$buf34 ),
    .Y(_8674_)
);

MUX2X1 _19658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [23]),
    .B(\datapath.registers.1226[6] [23]),
    .S(\datapath.idinstr_20_bF$buf33 ),
    .Y(_8675_)
);

MUX2X1 _19659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8675_),
    .B(_8674_),
    .S(\datapath.idinstr_21_bF$buf44 ),
    .Y(_8676_)
);

NAND2X1 _19660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf37 ),
    .B(_8676_),
    .Y(_8677_)
);

MUX2X1 _19661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [23]),
    .B(\datapath.registers.1226[0] [23]),
    .S(\datapath.idinstr_20_bF$buf32 ),
    .Y(_8678_)
);

MUX2X1 _19662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [23]),
    .B(\datapath.registers.1226[2] [23]),
    .S(\datapath.idinstr_20_bF$buf31 ),
    .Y(_8679_)
);

MUX2X1 _19663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8679_),
    .B(_8678_),
    .S(\datapath.idinstr_21_bF$buf43 ),
    .Y(_8680_)
);

NAND2X1 _19664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf0),
    .B(_8680_),
    .Y(_8681_)
);

AOI21X1 _19665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8677_),
    .B(_8681_),
    .C(\datapath.idinstr_23_bF$buf2 ),
    .Y(_8682_)
);

OAI21X1 _19666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8682_),
    .B(_8673_),
    .C(_7607__bF$buf0),
    .Y(_8683_)
);

AOI21X1 _19667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8662_),
    .B(_8683_),
    .C(_7614__bF$buf1),
    .Y(\datapath.registers.regb_data [23])
);

MUX2X1 _19668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [24]),
    .B(\datapath.registers.1226[24] [24]),
    .S(\datapath.idinstr_20_bF$buf30 ),
    .Y(_8684_)
);

MUX2X1 _19669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [24]),
    .B(\datapath.registers.1226[26] [24]),
    .S(\datapath.idinstr_20_bF$buf29 ),
    .Y(_8685_)
);

MUX2X1 _19670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8685_),
    .B(_8684_),
    .S(\datapath.idinstr_21_bF$buf42 ),
    .Y(_8686_)
);

NAND2X1 _19671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf10),
    .B(_8686_),
    .Y(_8687_)
);

MUX2X1 _19672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [24]),
    .B(\datapath.registers.1226[28] [24]),
    .S(\datapath.idinstr_20_bF$buf28 ),
    .Y(_8688_)
);

MUX2X1 _19673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [24]),
    .B(\datapath.registers.1226[30] [24]),
    .S(\datapath.idinstr_20_bF$buf27 ),
    .Y(_8689_)
);

MUX2X1 _19674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8689_),
    .B(_8688_),
    .S(\datapath.idinstr_21_bF$buf41 ),
    .Y(_8690_)
);

NAND2X1 _19675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf36 ),
    .B(_8690_),
    .Y(_8691_)
);

AOI21X1 _19676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8687_),
    .B(_8691_),
    .C(_7612__bF$buf6),
    .Y(_8692_)
);

MUX2X1 _19677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [24]),
    .B(\datapath.registers.1226[16] [24]),
    .S(\datapath.idinstr_21_bF$buf40 ),
    .Y(_8693_)
);

NAND2X1 _19678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf6),
    .B(_8693_),
    .Y(_8694_)
);

MUX2X1 _19679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [24]),
    .B(\datapath.registers.1226[17] [24]),
    .S(\datapath.idinstr_21_bF$buf39 ),
    .Y(_8695_)
);

AOI21X1 _19680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf26 ),
    .B(_8695_),
    .C(\datapath.idinstr_22_bF$buf35 ),
    .Y(_8696_)
);

NAND2X1 _19681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8694_),
    .B(_8696_),
    .Y(_8697_)
);

MUX2X1 _19682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [24]),
    .B(\datapath.registers.1226[20] [24]),
    .S(\datapath.idinstr_21_bF$buf38 ),
    .Y(_8698_)
);

NAND2X1 _19683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf5),
    .B(_8698_),
    .Y(_8699_)
);

MUX2X1 _19684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [24]),
    .B(\datapath.registers.1226[21] [24]),
    .S(\datapath.idinstr_21_bF$buf37 ),
    .Y(_8700_)
);

AOI21X1 _19685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf25 ),
    .B(_8700_),
    .C(_7611__bF$buf9),
    .Y(_8701_)
);

NAND2X1 _19686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8699_),
    .B(_8701_),
    .Y(_8702_)
);

AOI21X1 _19687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8697_),
    .B(_8702_),
    .C(\datapath.idinstr_23_bF$buf1 ),
    .Y(_8703_)
);

OAI21X1 _19688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8692_),
    .B(_8703_),
    .C(\datapath.idinstr_24_bF$buf0 ),
    .Y(_8704_)
);

MUX2X1 _19689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [24]),
    .B(\datapath.registers.1226[8] [24]),
    .S(\datapath.idinstr_20_bF$buf24 ),
    .Y(_8705_)
);

MUX2X1 _19690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [24]),
    .B(\datapath.registers.1226[10] [24]),
    .S(\datapath.idinstr_20_bF$buf23 ),
    .Y(_8706_)
);

MUX2X1 _19691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8706_),
    .B(_8705_),
    .S(\datapath.idinstr_21_bF$buf36 ),
    .Y(_8707_)
);

NAND2X1 _19692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf8),
    .B(_8707_),
    .Y(_8708_)
);

MUX2X1 _19693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [24]),
    .B(\datapath.registers.1226[12] [24]),
    .S(\datapath.idinstr_20_bF$buf22 ),
    .Y(_8709_)
);

MUX2X1 _19694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [24]),
    .B(\datapath.registers.1226[14] [24]),
    .S(\datapath.idinstr_20_bF$buf21 ),
    .Y(_8710_)
);

MUX2X1 _19695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8710_),
    .B(_8709_),
    .S(\datapath.idinstr_21_bF$buf35 ),
    .Y(_8711_)
);

NAND2X1 _19696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf34 ),
    .B(_8711_),
    .Y(_8712_)
);

AOI21X1 _19697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8708_),
    .B(_8712_),
    .C(_7612__bF$buf5),
    .Y(_8713_)
);

INVX1 _19698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [24]),
    .Y(_8714_)
);

AOI21X1 _19699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [24]),
    .B(\datapath.idinstr_22_bF$buf33 ),
    .C(_7608__bF$buf4),
    .Y(_8715_)
);

OAI21X1 _19700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8714_),
    .B(\datapath.idinstr_22_bF$buf32 ),
    .C(_8715_),
    .Y(_8716_)
);

INVX1 _19701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [24]),
    .Y(_8717_)
);

AOI21X1 _19702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [24]),
    .B(\datapath.idinstr_22_bF$buf31 ),
    .C(\datapath.idinstr_20_bF$buf20 ),
    .Y(_8718_)
);

OAI21X1 _19703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8717_),
    .B(\datapath.idinstr_22_bF$buf30 ),
    .C(_8718_),
    .Y(_8719_)
);

NAND3X1 _19704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf0),
    .B(_8719_),
    .C(_8716_),
    .Y(_8720_)
);

INVX1 _19705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [24]),
    .Y(_8721_)
);

AOI21X1 _19706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [24]),
    .B(\datapath.idinstr_22_bF$buf29 ),
    .C(_7608__bF$buf3),
    .Y(_8722_)
);

OAI21X1 _19707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8721_),
    .B(\datapath.idinstr_22_bF$buf28 ),
    .C(_8722_),
    .Y(_8723_)
);

INVX1 _19708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[2] [24]),
    .Y(_8724_)
);

AOI21X1 _19709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[6] [24]),
    .B(\datapath.idinstr_22_bF$buf27 ),
    .C(\datapath.idinstr_20_bF$buf19 ),
    .Y(_8725_)
);

OAI21X1 _19710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8724_),
    .B(\datapath.idinstr_22_bF$buf26 ),
    .C(_8725_),
    .Y(_8726_)
);

NAND3X1 _19711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf34 ),
    .B(_8726_),
    .C(_8723_),
    .Y(_8727_)
);

AOI21X1 _19712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8720_),
    .B(_8727_),
    .C(\datapath.idinstr_23_bF$buf0 ),
    .Y(_8728_)
);

OAI21X1 _19713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8713_),
    .B(_8728_),
    .C(_7607__bF$buf4),
    .Y(_8729_)
);

AOI21X1 _19714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8704_),
    .B(_8729_),
    .C(_7614__bF$buf0),
    .Y(\datapath.registers.regb_data [24])
);

MUX2X1 _19715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [25]),
    .B(\datapath.registers.1226[24] [25]),
    .S(\datapath.idinstr_20_bF$buf18 ),
    .Y(_8730_)
);

MUX2X1 _19716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [25]),
    .B(\datapath.registers.1226[26] [25]),
    .S(\datapath.idinstr_20_bF$buf17 ),
    .Y(_8731_)
);

MUX2X1 _19717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8731_),
    .B(_8730_),
    .S(\datapath.idinstr_21_bF$buf33 ),
    .Y(_8732_)
);

NAND2X1 _19718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf7),
    .B(_8732_),
    .Y(_8733_)
);

MUX2X1 _19719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [25]),
    .B(\datapath.registers.1226[28] [25]),
    .S(\datapath.idinstr_20_bF$buf16 ),
    .Y(_8734_)
);

MUX2X1 _19720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [25]),
    .B(\datapath.registers.1226[30] [25]),
    .S(\datapath.idinstr_20_bF$buf15 ),
    .Y(_8735_)
);

MUX2X1 _19721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8735_),
    .B(_8734_),
    .S(\datapath.idinstr_21_bF$buf32 ),
    .Y(_8736_)
);

NAND2X1 _19722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf25 ),
    .B(_8736_),
    .Y(_8737_)
);

AOI21X1 _19723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8733_),
    .B(_8737_),
    .C(_7612__bF$buf4),
    .Y(_8738_)
);

MUX2X1 _19724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [25]),
    .B(\datapath.registers.1226[16] [25]),
    .S(\datapath.idinstr_21_bF$buf31 ),
    .Y(_8739_)
);

NAND2X1 _19725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf2),
    .B(_8739_),
    .Y(_8740_)
);

MUX2X1 _19726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [25]),
    .B(\datapath.registers.1226[17] [25]),
    .S(\datapath.idinstr_21_bF$buf30 ),
    .Y(_8741_)
);

AOI21X1 _19727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf14 ),
    .B(_8741_),
    .C(\datapath.idinstr_22_bF$buf24 ),
    .Y(_8742_)
);

NAND2X1 _19728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8740_),
    .B(_8742_),
    .Y(_8743_)
);

MUX2X1 _19729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [25]),
    .B(\datapath.registers.1226[20] [25]),
    .S(\datapath.idinstr_21_bF$buf29 ),
    .Y(_8744_)
);

NAND2X1 _19730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf1),
    .B(_8744_),
    .Y(_8745_)
);

MUX2X1 _19731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [25]),
    .B(\datapath.registers.1226[21] [25]),
    .S(\datapath.idinstr_21_bF$buf28 ),
    .Y(_8746_)
);

AOI21X1 _19732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf13 ),
    .B(_8746_),
    .C(_7611__bF$buf6),
    .Y(_8747_)
);

NAND2X1 _19733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8745_),
    .B(_8747_),
    .Y(_8748_)
);

AOI21X1 _19734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8743_),
    .B(_8748_),
    .C(\datapath.idinstr_23_bF$buf7 ),
    .Y(_8749_)
);

OAI21X1 _19735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8738_),
    .B(_8749_),
    .C(\datapath.idinstr_24_bF$buf5 ),
    .Y(_8750_)
);

INVX1 _19736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [25]),
    .Y(_8751_)
);

AOI21X1 _19737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [25]),
    .B(\datapath.idinstr_22_bF$buf23 ),
    .C(_7608__bF$buf0),
    .Y(_8752_)
);

OAI21X1 _19738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8751_),
    .B(\datapath.idinstr_22_bF$buf22 ),
    .C(_8752_),
    .Y(_8753_)
);

INVX1 _19739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [25]),
    .Y(_8754_)
);

AOI21X1 _19740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [25]),
    .B(\datapath.idinstr_22_bF$buf21 ),
    .C(\datapath.idinstr_20_bF$buf12 ),
    .Y(_8755_)
);

OAI21X1 _19741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8754_),
    .B(\datapath.idinstr_22_bF$buf20 ),
    .C(_8755_),
    .Y(_8756_)
);

NAND3X1 _19742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf4),
    .B(_8756_),
    .C(_8753_),
    .Y(_8757_)
);

INVX1 _19743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [25]),
    .Y(_8758_)
);

AOI21X1 _19744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [25]),
    .B(\datapath.idinstr_22_bF$buf19 ),
    .C(_7608__bF$buf10),
    .Y(_8759_)
);

OAI21X1 _19745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8758_),
    .B(\datapath.idinstr_22_bF$buf18 ),
    .C(_8759_),
    .Y(_8760_)
);

INVX1 _19746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[10] [25]),
    .Y(_8761_)
);

AOI21X1 _19747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [25]),
    .B(\datapath.idinstr_22_bF$buf17 ),
    .C(\datapath.idinstr_20_bF$buf11 ),
    .Y(_8762_)
);

OAI21X1 _19748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8761_),
    .B(\datapath.idinstr_22_bF$buf16 ),
    .C(_8762_),
    .Y(_8763_)
);

NAND3X1 _19749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf27 ),
    .B(_8763_),
    .C(_8760_),
    .Y(_8764_)
);

AOI21X1 _19750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8757_),
    .B(_8764_),
    .C(_7612__bF$buf3),
    .Y(_8765_)
);

MUX2X1 _19751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [25]),
    .B(\datapath.registers.1226[0] [25]),
    .S(\datapath.idinstr_20_bF$buf10 ),
    .Y(_8766_)
);

MUX2X1 _19752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [25]),
    .B(\datapath.registers.1226[2] [25]),
    .S(\datapath.idinstr_20_bF$buf9 ),
    .Y(_8767_)
);

MUX2X1 _19753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8767_),
    .B(_8766_),
    .S(\datapath.idinstr_21_bF$buf26 ),
    .Y(_8768_)
);

NAND2X1 _19754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf5),
    .B(_8768_),
    .Y(_8769_)
);

MUX2X1 _19755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [25]),
    .B(\datapath.registers.1226[4] [25]),
    .S(\datapath.idinstr_20_bF$buf8 ),
    .Y(_8770_)
);

MUX2X1 _19756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [25]),
    .B(\datapath.registers.1226[6] [25]),
    .S(\datapath.idinstr_20_bF$buf7 ),
    .Y(_8771_)
);

MUX2X1 _19757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8771_),
    .B(_8770_),
    .S(\datapath.idinstr_21_bF$buf25 ),
    .Y(_8772_)
);

NAND2X1 _19758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf15 ),
    .B(_8772_),
    .Y(_8773_)
);

AOI21X1 _19759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8769_),
    .B(_8773_),
    .C(\datapath.idinstr_23_bF$buf6 ),
    .Y(_8774_)
);

OAI21X1 _19760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8774_),
    .B(_8765_),
    .C(_7607__bF$buf3),
    .Y(_8775_)
);

AOI21X1 _19761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8750_),
    .B(_8775_),
    .C(_7614__bF$buf4),
    .Y(\datapath.registers.regb_data [25])
);

MUX2X1 _19762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [26]),
    .B(\datapath.registers.1226[24] [26]),
    .S(\datapath.idinstr_20_bF$buf6 ),
    .Y(_8776_)
);

MUX2X1 _19763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [26]),
    .B(\datapath.registers.1226[26] [26]),
    .S(\datapath.idinstr_20_bF$buf5 ),
    .Y(_8777_)
);

MUX2X1 _19764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8777_),
    .B(_8776_),
    .S(\datapath.idinstr_21_bF$buf24 ),
    .Y(_8778_)
);

NAND2X1 _19765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf4),
    .B(_8778_),
    .Y(_8779_)
);

MUX2X1 _19766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [26]),
    .B(\datapath.registers.1226[28] [26]),
    .S(\datapath.idinstr_20_bF$buf4 ),
    .Y(_8780_)
);

MUX2X1 _19767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [26]),
    .B(\datapath.registers.1226[30] [26]),
    .S(\datapath.idinstr_20_bF$buf3 ),
    .Y(_8781_)
);

MUX2X1 _19768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8781_),
    .B(_8780_),
    .S(\datapath.idinstr_21_bF$buf23 ),
    .Y(_8782_)
);

NAND2X1 _19769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf14 ),
    .B(_8782_),
    .Y(_8783_)
);

AOI21X1 _19770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8779_),
    .B(_8783_),
    .C(_7612__bF$buf2),
    .Y(_8784_)
);

MUX2X1 _19771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [26]),
    .B(\datapath.registers.1226[16] [26]),
    .S(\datapath.idinstr_21_bF$buf22 ),
    .Y(_8785_)
);

NAND2X1 _19772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf9),
    .B(_8785_),
    .Y(_8786_)
);

MUX2X1 _19773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [26]),
    .B(\datapath.registers.1226[17] [26]),
    .S(\datapath.idinstr_21_bF$buf21 ),
    .Y(_8787_)
);

AOI21X1 _19774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf2 ),
    .B(_8787_),
    .C(\datapath.idinstr_22_bF$buf13 ),
    .Y(_8788_)
);

NAND2X1 _19775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8786_),
    .B(_8788_),
    .Y(_8789_)
);

MUX2X1 _19776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [26]),
    .B(\datapath.registers.1226[20] [26]),
    .S(\datapath.idinstr_21_bF$buf20 ),
    .Y(_8790_)
);

NAND2X1 _19777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf8),
    .B(_8790_),
    .Y(_8791_)
);

MUX2X1 _19778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [26]),
    .B(\datapath.registers.1226[21] [26]),
    .S(\datapath.idinstr_21_bF$buf19 ),
    .Y(_8792_)
);

AOI21X1 _19779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf1 ),
    .B(_8792_),
    .C(_7611__bF$buf3),
    .Y(_8793_)
);

NAND2X1 _19780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8791_),
    .B(_8793_),
    .Y(_8794_)
);

AOI21X1 _19781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8789_),
    .B(_8794_),
    .C(\datapath.idinstr_23_bF$buf5 ),
    .Y(_8795_)
);

OAI21X1 _19782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8784_),
    .B(_8795_),
    .C(\datapath.idinstr_24_bF$buf4 ),
    .Y(_8796_)
);

MUX2X1 _19783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [26]),
    .B(\datapath.registers.1226[8] [26]),
    .S(\datapath.idinstr_20_bF$buf0 ),
    .Y(_8797_)
);

MUX2X1 _19784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [26]),
    .B(\datapath.registers.1226[10] [26]),
    .S(\datapath.idinstr_20_bF$buf55 ),
    .Y(_8798_)
);

MUX2X1 _19785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8798_),
    .B(_8797_),
    .S(\datapath.idinstr_21_bF$buf18 ),
    .Y(_8799_)
);

NAND2X1 _19786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf2),
    .B(_8799_),
    .Y(_8800_)
);

NOR2X1 _19787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7360_),
    .B(_7608__bF$buf7),
    .Y(_8801_)
);

OAI21X1 _19788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7362_),
    .B(\datapath.idinstr_20_bF$buf54 ),
    .C(\datapath.idinstr_21_bF$buf17 ),
    .Y(_8802_)
);

NAND2X1 _19789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [26]),
    .B(_7608__bF$buf6),
    .Y(_8803_)
);

AOI21X1 _19790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [26]),
    .B(\datapath.idinstr_20_bF$buf53 ),
    .C(\datapath.idinstr_21_bF$buf16 ),
    .Y(_8804_)
);

AOI21X1 _19791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8804_),
    .B(_8803_),
    .C(_7611__bF$buf1),
    .Y(_8805_)
);

OAI21X1 _19792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8801_),
    .B(_8802_),
    .C(_8805_),
    .Y(_8806_)
);

AOI21X1 _19793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8806_),
    .B(_8800_),
    .C(_7612__bF$buf1),
    .Y(_8807_)
);

MUX2X1 _19794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [26]),
    .B(\datapath.registers.1226[4] [26]),
    .S(\datapath.idinstr_20_bF$buf52 ),
    .Y(_8808_)
);

MUX2X1 _19795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [26]),
    .B(\datapath.registers.1226[6] [26]),
    .S(\datapath.idinstr_20_bF$buf51 ),
    .Y(_8809_)
);

MUX2X1 _19796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8809_),
    .B(_8808_),
    .S(\datapath.idinstr_21_bF$buf15 ),
    .Y(_8810_)
);

NAND2X1 _19797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf12 ),
    .B(_8810_),
    .Y(_8811_)
);

MUX2X1 _19798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [26]),
    .B(\datapath.registers.1226[0] [26]),
    .S(\datapath.idinstr_20_bF$buf50 ),
    .Y(_8812_)
);

MUX2X1 _19799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [26]),
    .B(\datapath.registers.1226[2] [26]),
    .S(\datapath.idinstr_20_bF$buf49 ),
    .Y(_8813_)
);

MUX2X1 _19800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8813_),
    .B(_8812_),
    .S(\datapath.idinstr_21_bF$buf14 ),
    .Y(_8814_)
);

NAND2X1 _19801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf0),
    .B(_8814_),
    .Y(_8815_)
);

AOI21X1 _19802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8811_),
    .B(_8815_),
    .C(\datapath.idinstr_23_bF$buf4 ),
    .Y(_8816_)
);

OAI21X1 _19803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8816_),
    .B(_8807_),
    .C(_7607__bF$buf2),
    .Y(_8817_)
);

AOI21X1 _19804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8796_),
    .B(_8817_),
    .C(_7614__bF$buf3),
    .Y(\datapath.registers.regb_data [26])
);

MUX2X1 _19805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [27]),
    .B(\datapath.registers.1226[24] [27]),
    .S(\datapath.idinstr_20_bF$buf48 ),
    .Y(_8818_)
);

MUX2X1 _19806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [27]),
    .B(\datapath.registers.1226[26] [27]),
    .S(\datapath.idinstr_20_bF$buf47 ),
    .Y(_8819_)
);

MUX2X1 _19807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8819_),
    .B(_8818_),
    .S(\datapath.idinstr_21_bF$buf13 ),
    .Y(_8820_)
);

NAND2X1 _19808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf10),
    .B(_8820_),
    .Y(_8821_)
);

MUX2X1 _19809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [27]),
    .B(\datapath.registers.1226[28] [27]),
    .S(\datapath.idinstr_20_bF$buf46 ),
    .Y(_8822_)
);

MUX2X1 _19810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [27]),
    .B(\datapath.registers.1226[30] [27]),
    .S(\datapath.idinstr_20_bF$buf45 ),
    .Y(_8823_)
);

MUX2X1 _19811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8823_),
    .B(_8822_),
    .S(\datapath.idinstr_21_bF$buf12 ),
    .Y(_8824_)
);

NAND2X1 _19812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf11 ),
    .B(_8824_),
    .Y(_8825_)
);

AOI21X1 _19813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8821_),
    .B(_8825_),
    .C(_7612__bF$buf0),
    .Y(_8826_)
);

MUX2X1 _19814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [27]),
    .B(\datapath.registers.1226[16] [27]),
    .S(\datapath.idinstr_21_bF$buf11 ),
    .Y(_8827_)
);

NAND2X1 _19815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf5),
    .B(_8827_),
    .Y(_8828_)
);

MUX2X1 _19816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [27]),
    .B(\datapath.registers.1226[17] [27]),
    .S(\datapath.idinstr_21_bF$buf10 ),
    .Y(_8829_)
);

AOI21X1 _19817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf44 ),
    .B(_8829_),
    .C(\datapath.idinstr_22_bF$buf10 ),
    .Y(_8830_)
);

NAND2X1 _19818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8828_),
    .B(_8830_),
    .Y(_8831_)
);

MUX2X1 _19819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [27]),
    .B(\datapath.registers.1226[20] [27]),
    .S(\datapath.idinstr_21_bF$buf9 ),
    .Y(_8832_)
);

NAND2X1 _19820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf4),
    .B(_8832_),
    .Y(_8833_)
);

MUX2X1 _19821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [27]),
    .B(\datapath.registers.1226[21] [27]),
    .S(\datapath.idinstr_21_bF$buf8 ),
    .Y(_8834_)
);

AOI21X1 _19822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf43 ),
    .B(_8834_),
    .C(_7611__bF$buf9),
    .Y(_8835_)
);

NAND2X1 _19823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8833_),
    .B(_8835_),
    .Y(_8836_)
);

AOI21X1 _19824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8831_),
    .B(_8836_),
    .C(\datapath.idinstr_23_bF$buf3 ),
    .Y(_8837_)
);

OAI21X1 _19825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8826_),
    .B(_8837_),
    .C(\datapath.idinstr_24_bF$buf3 ),
    .Y(_8838_)
);

MUX2X1 _19826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [27]),
    .B(\datapath.registers.1226[8] [27]),
    .S(\datapath.idinstr_20_bF$buf42 ),
    .Y(_8839_)
);

MUX2X1 _19827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [27]),
    .B(\datapath.registers.1226[10] [27]),
    .S(\datapath.idinstr_20_bF$buf41 ),
    .Y(_8840_)
);

MUX2X1 _19828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8840_),
    .B(_8839_),
    .S(\datapath.idinstr_21_bF$buf7 ),
    .Y(_8841_)
);

NAND2X1 _19829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf8),
    .B(_8841_),
    .Y(_8842_)
);

AND2X2 _19830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [27]),
    .B(\datapath.idinstr_20_bF$buf40 ),
    .Y(_8843_)
);

INVX1 _19831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [27]),
    .Y(_8844_)
);

OAI21X1 _19832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8844_),
    .B(\datapath.idinstr_20_bF$buf39 ),
    .C(\datapath.idinstr_21_bF$buf6 ),
    .Y(_8845_)
);

NAND2X1 _19833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [27]),
    .B(_7608__bF$buf3),
    .Y(_8846_)
);

AOI21X1 _19834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [27]),
    .B(\datapath.idinstr_20_bF$buf38 ),
    .C(\datapath.idinstr_21_bF$buf5 ),
    .Y(_8847_)
);

AOI21X1 _19835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8847_),
    .B(_8846_),
    .C(_7611__bF$buf7),
    .Y(_8848_)
);

OAI21X1 _19836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8843_),
    .B(_8845_),
    .C(_8848_),
    .Y(_8849_)
);

AOI21X1 _19837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8849_),
    .B(_8842_),
    .C(_7612__bF$buf7),
    .Y(_8850_)
);

MUX2X1 _19838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [27]),
    .B(\datapath.registers.1226[4] [27]),
    .S(\datapath.idinstr_20_bF$buf37 ),
    .Y(_8851_)
);

MUX2X1 _19839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [27]),
    .B(\datapath.registers.1226[6] [27]),
    .S(\datapath.idinstr_20_bF$buf36 ),
    .Y(_8852_)
);

MUX2X1 _19840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8852_),
    .B(_8851_),
    .S(\datapath.idinstr_21_bF$buf4 ),
    .Y(_8853_)
);

NAND2X1 _19841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf9 ),
    .B(_8853_),
    .Y(_8854_)
);

MUX2X1 _19842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [27]),
    .B(\datapath.registers.1226[0] [27]),
    .S(\datapath.idinstr_20_bF$buf35 ),
    .Y(_8855_)
);

MUX2X1 _19843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [27]),
    .B(\datapath.registers.1226[2] [27]),
    .S(\datapath.idinstr_20_bF$buf34 ),
    .Y(_8856_)
);

MUX2X1 _19844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8856_),
    .B(_8855_),
    .S(\datapath.idinstr_21_bF$buf3 ),
    .Y(_8857_)
);

NAND2X1 _19845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf6),
    .B(_8857_),
    .Y(_8858_)
);

AOI21X1 _19846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8854_),
    .B(_8858_),
    .C(\datapath.idinstr_23_bF$buf2 ),
    .Y(_8859_)
);

OAI21X1 _19847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8859_),
    .B(_8850_),
    .C(_7607__bF$buf1),
    .Y(_8860_)
);

AOI21X1 _19848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8838_),
    .B(_8860_),
    .C(_7614__bF$buf2),
    .Y(\datapath.registers.regb_data [27])
);

MUX2X1 _19849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [28]),
    .B(\datapath.registers.1226[8] [28]),
    .S(\datapath.idinstr_20_bF$buf33 ),
    .Y(_8861_)
);

MUX2X1 _19850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [28]),
    .B(\datapath.registers.1226[10] [28]),
    .S(\datapath.idinstr_20_bF$buf32 ),
    .Y(_8862_)
);

MUX2X1 _19851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8862_),
    .B(_8861_),
    .S(\datapath.idinstr_21_bF$buf2 ),
    .Y(_8863_)
);

NAND2X1 _19852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf5),
    .B(_8863_),
    .Y(_8864_)
);

AND2X2 _19853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [28]),
    .B(\datapath.idinstr_20_bF$buf31 ),
    .Y(_8865_)
);

INVX1 _19854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [28]),
    .Y(_8866_)
);

OAI21X1 _19855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8866_),
    .B(\datapath.idinstr_20_bF$buf30 ),
    .C(\datapath.idinstr_21_bF$buf1 ),
    .Y(_8867_)
);

NAND2X1 _19856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [28]),
    .B(_7608__bF$buf2),
    .Y(_8868_)
);

AOI21X1 _19857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [28]),
    .B(\datapath.idinstr_20_bF$buf29 ),
    .C(\datapath.idinstr_21_bF$buf0 ),
    .Y(_8869_)
);

AOI21X1 _19858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8869_),
    .B(_8868_),
    .C(_7611__bF$buf4),
    .Y(_8870_)
);

OAI21X1 _19859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8865_),
    .B(_8867_),
    .C(_8870_),
    .Y(_8871_)
);

AOI21X1 _19860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8871_),
    .B(_8864_),
    .C(_7612__bF$buf6),
    .Y(_8872_)
);

MUX2X1 _19861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [28]),
    .B(\datapath.registers.1226[4] [28]),
    .S(\datapath.idinstr_20_bF$buf28 ),
    .Y(_8873_)
);

MUX2X1 _19862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [28]),
    .B(\datapath.registers.1226[6] [28]),
    .S(\datapath.idinstr_20_bF$buf27 ),
    .Y(_8874_)
);

MUX2X1 _19863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8874_),
    .B(_8873_),
    .S(\datapath.idinstr_21_bF$buf44 ),
    .Y(_8875_)
);

NAND2X1 _19864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf8 ),
    .B(_8875_),
    .Y(_8876_)
);

MUX2X1 _19865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [28]),
    .B(\datapath.registers.1226[0] [28]),
    .S(\datapath.idinstr_20_bF$buf26 ),
    .Y(_8877_)
);

MUX2X1 _19866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [28]),
    .B(\datapath.registers.1226[2] [28]),
    .S(\datapath.idinstr_20_bF$buf25 ),
    .Y(_8878_)
);

MUX2X1 _19867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8878_),
    .B(_8877_),
    .S(\datapath.idinstr_21_bF$buf43 ),
    .Y(_8879_)
);

NAND2X1 _19868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf3),
    .B(_8879_),
    .Y(_8880_)
);

AOI21X1 _19869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8876_),
    .B(_8880_),
    .C(\datapath.idinstr_23_bF$buf1 ),
    .Y(_8881_)
);

OAI21X1 _19870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8881_),
    .B(_8872_),
    .C(_7607__bF$buf0),
    .Y(_8882_)
);

INVX1 _19871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [28]),
    .Y(_8883_)
);

AOI21X1 _19872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [28]),
    .B(\datapath.idinstr_22_bF$buf7 ),
    .C(_7608__bF$buf1),
    .Y(_8884_)
);

OAI21X1 _19873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8883_),
    .B(\datapath.idinstr_22_bF$buf6 ),
    .C(_8884_),
    .Y(_8885_)
);

NAND2X1 _19874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [28]),
    .B(_7611__bF$buf2),
    .Y(_8886_)
);

AOI21X1 _19875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [28]),
    .B(\datapath.idinstr_22_bF$buf5 ),
    .C(\datapath.idinstr_20_bF$buf24 ),
    .Y(_8887_)
);

AOI21X1 _19876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8887_),
    .B(_8886_),
    .C(_7610__bF$buf3),
    .Y(_8888_)
);

NAND2X1 _19877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8885_),
    .B(_8888_),
    .Y(_8889_)
);

INVX1 _19878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [28]),
    .Y(_8890_)
);

AOI21X1 _19879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [28]),
    .B(\datapath.idinstr_22_bF$buf4 ),
    .C(_7608__bF$buf0),
    .Y(_8891_)
);

OAI21X1 _19880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8890_),
    .B(\datapath.idinstr_22_bF$buf3 ),
    .C(_8891_),
    .Y(_8892_)
);

AOI21X1 _19881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[28] [28]),
    .B(\datapath.idinstr_22_bF$buf2 ),
    .C(\datapath.idinstr_20_bF$buf23 ),
    .Y(_8893_)
);

OAI21X1 _19882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5751_),
    .B(\datapath.idinstr_22_bF$buf1 ),
    .C(_8893_),
    .Y(_8894_)
);

NAND3X1 _19883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf2),
    .B(_8894_),
    .C(_8892_),
    .Y(_8895_)
);

AOI21X1 _19884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8889_),
    .B(_8895_),
    .C(_7612__bF$buf5),
    .Y(_8896_)
);

MUX2X1 _19885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [28]),
    .B(\datapath.registers.1226[16] [28]),
    .S(\datapath.idinstr_20_bF$buf22 ),
    .Y(_8897_)
);

MUX2X1 _19886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [28]),
    .B(\datapath.registers.1226[18] [28]),
    .S(\datapath.idinstr_20_bF$buf21 ),
    .Y(_8898_)
);

MUX2X1 _19887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8898_),
    .B(_8897_),
    .S(\datapath.idinstr_21_bF$buf42 ),
    .Y(_8899_)
);

NAND2X1 _19888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf1),
    .B(_8899_),
    .Y(_8900_)
);

MUX2X1 _19889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [28]),
    .B(\datapath.registers.1226[20] [28]),
    .S(\datapath.idinstr_20_bF$buf20 ),
    .Y(_8901_)
);

MUX2X1 _19890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [28]),
    .B(\datapath.registers.1226[22] [28]),
    .S(\datapath.idinstr_20_bF$buf19 ),
    .Y(_8902_)
);

MUX2X1 _19891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8902_),
    .B(_8901_),
    .S(\datapath.idinstr_21_bF$buf41 ),
    .Y(_8903_)
);

NAND2X1 _19892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf0 ),
    .B(_8903_),
    .Y(_8904_)
);

AOI21X1 _19893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8900_),
    .B(_8904_),
    .C(\datapath.idinstr_23_bF$buf0 ),
    .Y(_8905_)
);

OAI21X1 _19894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8905_),
    .B(_8896_),
    .C(\datapath.idinstr_24_bF$buf2 ),
    .Y(_8906_)
);

AOI21X1 _19895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8906_),
    .B(_8882_),
    .C(_7614__bF$buf1),
    .Y(\datapath.registers.regb_data [28])
);

MUX2X1 _19896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [29]),
    .B(\datapath.registers.1226[24] [29]),
    .S(\datapath.idinstr_20_bF$buf18 ),
    .Y(_8907_)
);

MUX2X1 _19897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [29]),
    .B(\datapath.registers.1226[26] [29]),
    .S(\datapath.idinstr_20_bF$buf17 ),
    .Y(_8908_)
);

MUX2X1 _19898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8908_),
    .B(_8907_),
    .S(\datapath.idinstr_21_bF$buf40 ),
    .Y(_8909_)
);

NAND2X1 _19899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf0),
    .B(_8909_),
    .Y(_8910_)
);

MUX2X1 _19900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [29]),
    .B(\datapath.registers.1226[28] [29]),
    .S(\datapath.idinstr_20_bF$buf16 ),
    .Y(_8911_)
);

MUX2X1 _19901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [29]),
    .B(\datapath.registers.1226[30] [29]),
    .S(\datapath.idinstr_20_bF$buf15 ),
    .Y(_8912_)
);

MUX2X1 _19902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8912_),
    .B(_8911_),
    .S(\datapath.idinstr_21_bF$buf39 ),
    .Y(_8913_)
);

NAND2X1 _19903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf43 ),
    .B(_8913_),
    .Y(_8914_)
);

AOI21X1 _19904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8910_),
    .B(_8914_),
    .C(_7612__bF$buf4),
    .Y(_8915_)
);

MUX2X1 _19905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [29]),
    .B(\datapath.registers.1226[16] [29]),
    .S(\datapath.idinstr_21_bF$buf38 ),
    .Y(_8916_)
);

NAND2X1 _19906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf10),
    .B(_8916_),
    .Y(_8917_)
);

MUX2X1 _19907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [29]),
    .B(\datapath.registers.1226[17] [29]),
    .S(\datapath.idinstr_21_bF$buf37 ),
    .Y(_8918_)
);

AOI21X1 _19908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf14 ),
    .B(_8918_),
    .C(\datapath.idinstr_22_bF$buf42 ),
    .Y(_8919_)
);

NAND2X1 _19909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8917_),
    .B(_8919_),
    .Y(_8920_)
);

MUX2X1 _19910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [29]),
    .B(\datapath.registers.1226[20] [29]),
    .S(\datapath.idinstr_21_bF$buf36 ),
    .Y(_8921_)
);

NAND2X1 _19911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf9),
    .B(_8921_),
    .Y(_8922_)
);

MUX2X1 _19912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [29]),
    .B(\datapath.registers.1226[21] [29]),
    .S(\datapath.idinstr_21_bF$buf35 ),
    .Y(_8923_)
);

AOI21X1 _19913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf13 ),
    .B(_8923_),
    .C(_7611__bF$buf10),
    .Y(_8924_)
);

NAND2X1 _19914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8922_),
    .B(_8924_),
    .Y(_8925_)
);

AOI21X1 _19915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8920_),
    .B(_8925_),
    .C(\datapath.idinstr_23_bF$buf7 ),
    .Y(_8926_)
);

OAI21X1 _19916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8915_),
    .B(_8926_),
    .C(\datapath.idinstr_24_bF$buf1 ),
    .Y(_8927_)
);

MUX2X1 _19917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [29]),
    .B(\datapath.registers.1226[8] [29]),
    .S(\datapath.idinstr_20_bF$buf12 ),
    .Y(_8928_)
);

MUX2X1 _19918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [29]),
    .B(\datapath.registers.1226[10] [29]),
    .S(\datapath.idinstr_20_bF$buf11 ),
    .Y(_8929_)
);

MUX2X1 _19919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8929_),
    .B(_8928_),
    .S(\datapath.idinstr_21_bF$buf34 ),
    .Y(_8930_)
);

NAND2X1 _19920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf9),
    .B(_8930_),
    .Y(_8931_)
);

MUX2X1 _19921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [29]),
    .B(\datapath.registers.1226[12] [29]),
    .S(\datapath.idinstr_20_bF$buf10 ),
    .Y(_8932_)
);

MUX2X1 _19922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [29]),
    .B(\datapath.registers.1226[14] [29]),
    .S(\datapath.idinstr_20_bF$buf9 ),
    .Y(_8933_)
);

MUX2X1 _19923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8933_),
    .B(_8932_),
    .S(\datapath.idinstr_21_bF$buf33 ),
    .Y(_8934_)
);

NAND2X1 _19924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf41 ),
    .B(_8934_),
    .Y(_8935_)
);

AOI21X1 _19925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8931_),
    .B(_8935_),
    .C(_7612__bF$buf3),
    .Y(_8936_)
);

INVX1 _19926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [29]),
    .Y(_8937_)
);

AOI21X1 _19927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [29]),
    .B(\datapath.idinstr_22_bF$buf40 ),
    .C(_7608__bF$buf8),
    .Y(_8938_)
);

OAI21X1 _19928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8937_),
    .B(\datapath.idinstr_22_bF$buf39 ),
    .C(_8938_),
    .Y(_8939_)
);

INVX1 _19929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [29]),
    .Y(_8940_)
);

AOI21X1 _19930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [29]),
    .B(\datapath.idinstr_22_bF$buf38 ),
    .C(\datapath.idinstr_20_bF$buf8 ),
    .Y(_8941_)
);

OAI21X1 _19931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8940_),
    .B(\datapath.idinstr_22_bF$buf37 ),
    .C(_8941_),
    .Y(_8942_)
);

NAND3X1 _19932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf1),
    .B(_8942_),
    .C(_8939_),
    .Y(_8943_)
);

INVX1 _19933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [29]),
    .Y(_8944_)
);

AOI21X1 _19934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [29]),
    .B(\datapath.idinstr_22_bF$buf36 ),
    .C(_7608__bF$buf7),
    .Y(_8945_)
);

OAI21X1 _19935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8944_),
    .B(\datapath.idinstr_22_bF$buf35 ),
    .C(_8945_),
    .Y(_8946_)
);

INVX1 _19936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[2] [29]),
    .Y(_8947_)
);

AOI21X1 _19937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[6] [29]),
    .B(\datapath.idinstr_22_bF$buf34 ),
    .C(\datapath.idinstr_20_bF$buf7 ),
    .Y(_8948_)
);

OAI21X1 _19938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8947_),
    .B(\datapath.idinstr_22_bF$buf33 ),
    .C(_8948_),
    .Y(_8949_)
);

NAND3X1 _19939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf32 ),
    .B(_8949_),
    .C(_8946_),
    .Y(_8950_)
);

AOI21X1 _19940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8943_),
    .B(_8950_),
    .C(\datapath.idinstr_23_bF$buf6 ),
    .Y(_8951_)
);

OAI21X1 _19941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8936_),
    .B(_8951_),
    .C(_7607__bF$buf4),
    .Y(_8952_)
);

AOI21X1 _19942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8927_),
    .B(_8952_),
    .C(_7614__bF$buf0),
    .Y(\datapath.registers.regb_data [29])
);

MUX2X1 _19943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [30]),
    .B(\datapath.registers.1226[24] [30]),
    .S(\datapath.idinstr_20_bF$buf6 ),
    .Y(_8953_)
);

MUX2X1 _19944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [30]),
    .B(\datapath.registers.1226[26] [30]),
    .S(\datapath.idinstr_20_bF$buf5 ),
    .Y(_8954_)
);

MUX2X1 _19945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8954_),
    .B(_8953_),
    .S(\datapath.idinstr_21_bF$buf31 ),
    .Y(_8955_)
);

NAND2X1 _19946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf8),
    .B(_8955_),
    .Y(_8956_)
);

MUX2X1 _19947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [30]),
    .B(\datapath.registers.1226[28] [30]),
    .S(\datapath.idinstr_20_bF$buf4 ),
    .Y(_8957_)
);

MUX2X1 _19948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [30]),
    .B(\datapath.registers.1226[30] [30]),
    .S(\datapath.idinstr_20_bF$buf3 ),
    .Y(_8958_)
);

MUX2X1 _19949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8958_),
    .B(_8957_),
    .S(\datapath.idinstr_21_bF$buf30 ),
    .Y(_8959_)
);

NAND2X1 _19950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf32 ),
    .B(_8959_),
    .Y(_8960_)
);

AOI21X1 _19951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8956_),
    .B(_8960_),
    .C(_7612__bF$buf2),
    .Y(_8961_)
);

MUX2X1 _19952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[18] [30]),
    .B(\datapath.registers.1226[16] [30]),
    .S(\datapath.idinstr_21_bF$buf29 ),
    .Y(_8962_)
);

NAND2X1 _19953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf6),
    .B(_8962_),
    .Y(_8963_)
);

MUX2X1 _19954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [30]),
    .B(\datapath.registers.1226[17] [30]),
    .S(\datapath.idinstr_21_bF$buf28 ),
    .Y(_8964_)
);

AOI21X1 _19955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf2 ),
    .B(_8964_),
    .C(\datapath.idinstr_22_bF$buf31 ),
    .Y(_8965_)
);

NAND2X1 _19956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8963_),
    .B(_8965_),
    .Y(_8966_)
);

MUX2X1 _19957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[22] [30]),
    .B(\datapath.registers.1226[20] [30]),
    .S(\datapath.idinstr_21_bF$buf27 ),
    .Y(_8967_)
);

NAND2X1 _19958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7608__bF$buf5),
    .B(_8967_),
    .Y(_8968_)
);

MUX2X1 _19959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [30]),
    .B(\datapath.registers.1226[21] [30]),
    .S(\datapath.idinstr_21_bF$buf26 ),
    .Y(_8969_)
);

AOI21X1 _19960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf1 ),
    .B(_8969_),
    .C(_7611__bF$buf7),
    .Y(_8970_)
);

NAND2X1 _19961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8968_),
    .B(_8970_),
    .Y(_8971_)
);

AOI21X1 _19962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8966_),
    .B(_8971_),
    .C(\datapath.idinstr_23_bF$buf5 ),
    .Y(_8972_)
);

OAI21X1 _19963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8961_),
    .B(_8972_),
    .C(\datapath.idinstr_24_bF$buf0 ),
    .Y(_8973_)
);

MUX2X1 _19964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [30]),
    .B(\datapath.registers.1226[8] [30]),
    .S(\datapath.idinstr_20_bF$buf0 ),
    .Y(_8974_)
);

MUX2X1 _19965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [30]),
    .B(\datapath.registers.1226[10] [30]),
    .S(\datapath.idinstr_20_bF$buf55 ),
    .Y(_8975_)
);

MUX2X1 _19966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8975_),
    .B(_8974_),
    .S(\datapath.idinstr_21_bF$buf25 ),
    .Y(_8976_)
);

NAND2X1 _19967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf6),
    .B(_8976_),
    .Y(_8977_)
);

AND2X2 _19968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[15] [30]),
    .B(\datapath.idinstr_20_bF$buf54 ),
    .Y(_8978_)
);

INVX1 _19969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[14] [30]),
    .Y(_8979_)
);

OAI21X1 _19970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8979_),
    .B(\datapath.idinstr_20_bF$buf53 ),
    .C(\datapath.idinstr_21_bF$buf24 ),
    .Y(_8980_)
);

NAND2X1 _19971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [30]),
    .B(_7608__bF$buf4),
    .Y(_8981_)
);

AOI21X1 _19972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [30]),
    .B(\datapath.idinstr_20_bF$buf52 ),
    .C(\datapath.idinstr_21_bF$buf23 ),
    .Y(_8982_)
);

AOI21X1 _19973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8982_),
    .B(_8981_),
    .C(_7611__bF$buf5),
    .Y(_8983_)
);

OAI21X1 _19974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8978_),
    .B(_8980_),
    .C(_8983_),
    .Y(_8984_)
);

AOI21X1 _19975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8984_),
    .B(_8977_),
    .C(_7612__bF$buf1),
    .Y(_8985_)
);

MUX2X1 _19976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [30]),
    .B(\datapath.registers.1226[4] [30]),
    .S(\datapath.idinstr_20_bF$buf51 ),
    .Y(_8986_)
);

MUX2X1 _19977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [30]),
    .B(\datapath.registers.1226[6] [30]),
    .S(\datapath.idinstr_20_bF$buf50 ),
    .Y(_8987_)
);

MUX2X1 _19978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8987_),
    .B(_8986_),
    .S(\datapath.idinstr_21_bF$buf22 ),
    .Y(_8988_)
);

NAND2X1 _19979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf30 ),
    .B(_8988_),
    .Y(_8989_)
);

MUX2X1 _19980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [30]),
    .B(\datapath.registers.1226[0] [30]),
    .S(\datapath.idinstr_20_bF$buf49 ),
    .Y(_8990_)
);

MUX2X1 _19981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [30]),
    .B(\datapath.registers.1226[2] [30]),
    .S(\datapath.idinstr_20_bF$buf48 ),
    .Y(_8991_)
);

MUX2X1 _19982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8991_),
    .B(_8990_),
    .S(\datapath.idinstr_21_bF$buf21 ),
    .Y(_8992_)
);

NAND2X1 _19983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf4),
    .B(_8992_),
    .Y(_8993_)
);

AOI21X1 _19984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8989_),
    .B(_8993_),
    .C(\datapath.idinstr_23_bF$buf4 ),
    .Y(_8994_)
);

OAI21X1 _19985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8994_),
    .B(_8985_),
    .C(_7607__bF$buf3),
    .Y(_8995_)
);

AOI21X1 _19986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8973_),
    .B(_8995_),
    .C(_7614__bF$buf4),
    .Y(\datapath.registers.regb_data [30])
);

MUX2X1 _19987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[9] [31]),
    .B(\datapath.registers.1226[8] [31]),
    .S(\datapath.idinstr_20_bF$buf47 ),
    .Y(_8996_)
);

MUX2X1 _19988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[11] [31]),
    .B(\datapath.registers.1226[10] [31]),
    .S(\datapath.idinstr_20_bF$buf46 ),
    .Y(_8997_)
);

MUX2X1 _19989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8997_),
    .B(_8996_),
    .S(\datapath.idinstr_21_bF$buf20 ),
    .Y(_8998_)
);

NAND2X1 _19990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf3),
    .B(_8998_),
    .Y(_8999_)
);

NOR2X1 _19991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7588_),
    .B(_7608__bF$buf3),
    .Y(_9000_)
);

OAI21X1 _19992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7590_),
    .B(\datapath.idinstr_20_bF$buf45 ),
    .C(\datapath.idinstr_21_bF$buf19 ),
    .Y(_9001_)
);

NAND2X1 _19993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [31]),
    .B(_7608__bF$buf2),
    .Y(_9002_)
);

AOI21X1 _19994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[13] [31]),
    .B(\datapath.idinstr_20_bF$buf44 ),
    .C(\datapath.idinstr_21_bF$buf18 ),
    .Y(_9003_)
);

AOI21X1 _19995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9003_),
    .B(_9002_),
    .C(_7611__bF$buf2),
    .Y(_9004_)
);

OAI21X1 _19996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9000_),
    .B(_9001_),
    .C(_9004_),
    .Y(_9005_)
);

AOI21X1 _19997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9005_),
    .B(_8999_),
    .C(_7612__bF$buf0),
    .Y(_9006_)
);

MUX2X1 _19998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[5] [31]),
    .B(\datapath.registers.1226[4] [31]),
    .S(\datapath.idinstr_20_bF$buf43 ),
    .Y(_9007_)
);

MUX2X1 _19999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[7] [31]),
    .B(\datapath.registers.1226[6] [31]),
    .S(\datapath.idinstr_20_bF$buf42 ),
    .Y(_9008_)
);

MUX2X1 _20000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9008_),
    .B(_9007_),
    .S(\datapath.idinstr_21_bF$buf17 ),
    .Y(_9009_)
);

NAND2X1 _20001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf29 ),
    .B(_9009_),
    .Y(_9010_)
);

MUX2X1 _20002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[1] [31]),
    .B(\datapath.registers.1226[0] [31]),
    .S(\datapath.idinstr_20_bF$buf41 ),
    .Y(_9011_)
);

MUX2X1 _20003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [31]),
    .B(\datapath.registers.1226[2] [31]),
    .S(\datapath.idinstr_20_bF$buf40 ),
    .Y(_9012_)
);

MUX2X1 _20004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9012_),
    .B(_9011_),
    .S(\datapath.idinstr_21_bF$buf16 ),
    .Y(_9013_)
);

NAND2X1 _20005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf1),
    .B(_9013_),
    .Y(_9014_)
);

AOI21X1 _20006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9010_),
    .B(_9014_),
    .C(\datapath.idinstr_23_bF$buf3 ),
    .Y(_9015_)
);

OAI21X1 _20007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9015_),
    .B(_9006_),
    .C(_7607__bF$buf2),
    .Y(_9016_)
);

INVX1 _20008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[27] [31]),
    .Y(_9017_)
);

AOI21X1 _20009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[31] [31]),
    .B(\datapath.idinstr_22_bF$buf28 ),
    .C(_7608__bF$buf1),
    .Y(_9018_)
);

OAI21X1 _20010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9017_),
    .B(\datapath.idinstr_22_bF$buf27 ),
    .C(_9018_),
    .Y(_9019_)
);

NAND2X1 _20011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[26] [31]),
    .B(_7611__bF$buf0),
    .Y(_9020_)
);

AOI21X1 _20012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[30] [31]),
    .B(\datapath.idinstr_22_bF$buf26 ),
    .C(\datapath.idinstr_20_bF$buf39 ),
    .Y(_9021_)
);

AOI21X1 _20013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9021_),
    .B(_9020_),
    .C(_7610__bF$buf0),
    .Y(_9022_)
);

NAND2X1 _20014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9019_),
    .B(_9022_),
    .Y(_9023_)
);

INVX1 _20015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[25] [31]),
    .Y(_9024_)
);

AOI21X1 _20016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[29] [31]),
    .B(\datapath.idinstr_22_bF$buf25 ),
    .C(_7608__bF$buf0),
    .Y(_9025_)
);

OAI21X1 _20017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9024_),
    .B(\datapath.idinstr_22_bF$buf24 ),
    .C(_9025_),
    .Y(_9026_)
);

AOI21X1 _20018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[28] [31]),
    .B(\datapath.idinstr_22_bF$buf23 ),
    .C(\datapath.idinstr_20_bF$buf38 ),
    .Y(_9027_)
);

OAI21X1 _20019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5755_),
    .B(\datapath.idinstr_22_bF$buf22 ),
    .C(_9027_),
    .Y(_9028_)
);

NAND3X1 _20020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7610__bF$buf4),
    .B(_9028_),
    .C(_9026_),
    .Y(_9029_)
);

AOI21X1 _20021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9023_),
    .B(_9029_),
    .C(_7612__bF$buf7),
    .Y(_9030_)
);

MUX2X1 _20022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[17] [31]),
    .B(\datapath.registers.1226[16] [31]),
    .S(\datapath.idinstr_20_bF$buf37 ),
    .Y(_9031_)
);

MUX2X1 _20023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[19] [31]),
    .B(\datapath.registers.1226[18] [31]),
    .S(\datapath.idinstr_20_bF$buf36 ),
    .Y(_9032_)
);

MUX2X1 _20024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9032_),
    .B(_9031_),
    .S(\datapath.idinstr_21_bF$buf15 ),
    .Y(_9033_)
);

NAND2X1 _20025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611__bF$buf10),
    .B(_9033_),
    .Y(_9034_)
);

MUX2X1 _20026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[21] [31]),
    .B(\datapath.registers.1226[20] [31]),
    .S(\datapath.idinstr_20_bF$buf35 ),
    .Y(_9035_)
);

MUX2X1 _20027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[23] [31]),
    .B(\datapath.registers.1226[22] [31]),
    .S(\datapath.idinstr_20_bF$buf34 ),
    .Y(_9036_)
);

MUX2X1 _20028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9036_),
    .B(_9035_),
    .S(\datapath.idinstr_21_bF$buf14 ),
    .Y(_9037_)
);

NAND2X1 _20029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf21 ),
    .B(_9037_),
    .Y(_9038_)
);

AOI21X1 _20030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9034_),
    .B(_9038_),
    .C(\datapath.idinstr_23_bF$buf2 ),
    .Y(_9039_)
);

OAI21X1 _20031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9039_),
    .B(_9030_),
    .C(\datapath.idinstr_24_bF$buf5 ),
    .Y(_9040_)
);

AOI21X1 _20032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9040_),
    .B(_9016_),
    .C(_7614__bF$buf3),
    .Y(\datapath.registers.regb_data [31])
);

NOR2X1 _20033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf5),
    .B(_6041__bF$buf2),
    .Y(_9041_)
);

NOR2X1 _20034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [0]),
    .B(_9041__bF$buf7),
    .Y(_9042_)
);

AOI21X1 _20035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf1),
    .B(_9041__bF$buf6),
    .C(_9042_),
    .Y(_4501_)
);

NOR2X1 _20036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [1]),
    .B(_9041__bF$buf5),
    .Y(_9043_)
);

AOI21X1 _20037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf1),
    .B(_9041__bF$buf4),
    .C(_9043_),
    .Y(_4512_)
);

NOR2X1 _20038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [2]),
    .B(_9041__bF$buf3),
    .Y(_9044_)
);

AOI21X1 _20039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf0),
    .B(_9041__bF$buf2),
    .C(_9044_),
    .Y(_4523_)
);

NOR2X1 _20040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [3]),
    .B(_9041__bF$buf1),
    .Y(_9045_)
);

AOI21X1 _20041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf2),
    .B(_9041__bF$buf0),
    .C(_9045_),
    .Y(_4526_)
);

NOR2X1 _20042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [4]),
    .B(_9041__bF$buf7),
    .Y(_9046_)
);

AOI21X1 _20043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf0),
    .B(_9041__bF$buf6),
    .C(_9046_),
    .Y(_4527_)
);

NOR2X1 _20044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [5]),
    .B(_9041__bF$buf5),
    .Y(_9047_)
);

AOI21X1 _20045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf0),
    .B(_9041__bF$buf4),
    .C(_9047_),
    .Y(_4528_)
);

NOR2X1 _20046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [6]),
    .B(_9041__bF$buf3),
    .Y(_9048_)
);

AOI21X1 _20047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf1),
    .B(_9041__bF$buf2),
    .C(_9048_),
    .Y(_4529_)
);

NOR2X1 _20048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [7]),
    .B(_9041__bF$buf1),
    .Y(_9049_)
);

AOI21X1 _20049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf1),
    .B(_9041__bF$buf0),
    .C(_9049_),
    .Y(_4530_)
);

NOR2X1 _20050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [8]),
    .B(_9041__bF$buf7),
    .Y(_9050_)
);

AOI21X1 _20051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf1),
    .B(_9041__bF$buf6),
    .C(_9050_),
    .Y(_4531_)
);

NOR2X1 _20052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [9]),
    .B(_9041__bF$buf5),
    .Y(_9051_)
);

AOI21X1 _20053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf0),
    .B(_9041__bF$buf4),
    .C(_9051_),
    .Y(_4532_)
);

NOR2X1 _20054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [10]),
    .B(_9041__bF$buf3),
    .Y(_9052_)
);

AOI21X1 _20055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf2),
    .B(_9041__bF$buf2),
    .C(_9052_),
    .Y(_4502_)
);

NOR2X1 _20056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [11]),
    .B(_9041__bF$buf1),
    .Y(_9053_)
);

AOI21X1 _20057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf0),
    .B(_9041__bF$buf0),
    .C(_9053_),
    .Y(_4503_)
);

NOR2X1 _20058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [12]),
    .B(_9041__bF$buf7),
    .Y(_9054_)
);

AOI21X1 _20059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf1),
    .B(_9041__bF$buf6),
    .C(_9054_),
    .Y(_4504_)
);

NOR2X1 _20060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [13]),
    .B(_9041__bF$buf5),
    .Y(_9055_)
);

AOI21X1 _20061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf1),
    .B(_9041__bF$buf4),
    .C(_9055_),
    .Y(_4505_)
);

NOR2X1 _20062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [14]),
    .B(_9041__bF$buf3),
    .Y(_9056_)
);

AOI21X1 _20063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf0),
    .B(_9041__bF$buf2),
    .C(_9056_),
    .Y(_4506_)
);

NOR2X1 _20064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [15]),
    .B(_9041__bF$buf1),
    .Y(_9057_)
);

AOI21X1 _20065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf0),
    .B(_9041__bF$buf0),
    .C(_9057_),
    .Y(_4507_)
);

NOR2X1 _20066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [16]),
    .B(_9041__bF$buf7),
    .Y(_9058_)
);

AOI21X1 _20067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf2),
    .B(_9041__bF$buf6),
    .C(_9058_),
    .Y(_4508_)
);

NOR2X1 _20068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [17]),
    .B(_9041__bF$buf5),
    .Y(_9059_)
);

AOI21X1 _20069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf1),
    .B(_9041__bF$buf4),
    .C(_9059_),
    .Y(_4509_)
);

NOR2X1 _20070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [18]),
    .B(_9041__bF$buf3),
    .Y(_9060_)
);

AOI21X1 _20071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf0),
    .B(_9041__bF$buf2),
    .C(_9060_),
    .Y(_4510_)
);

NOR2X1 _20072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [19]),
    .B(_9041__bF$buf1),
    .Y(_9061_)
);

AOI21X1 _20073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf0),
    .B(_9041__bF$buf0),
    .C(_9061_),
    .Y(_4511_)
);

NOR2X1 _20074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [20]),
    .B(_9041__bF$buf7),
    .Y(_9062_)
);

AOI21X1 _20075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf1),
    .B(_9041__bF$buf6),
    .C(_9062_),
    .Y(_4513_)
);

NOR2X1 _20076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [21]),
    .B(_9041__bF$buf5),
    .Y(_9063_)
);

AOI21X1 _20077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf2),
    .B(_9041__bF$buf4),
    .C(_9063_),
    .Y(_4514_)
);

NOR2X1 _20078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [22]),
    .B(_9041__bF$buf3),
    .Y(_9064_)
);

AOI21X1 _20079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf1),
    .B(_9041__bF$buf2),
    .C(_9064_),
    .Y(_4515_)
);

NOR2X1 _20080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [23]),
    .B(_9041__bF$buf1),
    .Y(_9065_)
);

AOI21X1 _20081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf0),
    .B(_9041__bF$buf0),
    .C(_9065_),
    .Y(_4516_)
);

NOR2X1 _20082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [24]),
    .B(_9041__bF$buf7),
    .Y(_9066_)
);

AOI21X1 _20083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf0),
    .B(_9041__bF$buf6),
    .C(_9066_),
    .Y(_4517_)
);

NOR2X1 _20084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [25]),
    .B(_9041__bF$buf5),
    .Y(_9067_)
);

AOI21X1 _20085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486__bF$buf1),
    .B(_9041__bF$buf4),
    .C(_9067_),
    .Y(_4518_)
);

NOR2X1 _20086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [26]),
    .B(_9041__bF$buf3),
    .Y(_9068_)
);

AOI21X1 _20087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf0),
    .B(_9041__bF$buf2),
    .C(_9068_),
    .Y(_4519_)
);

NOR2X1 _20088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [27]),
    .B(_9041__bF$buf1),
    .Y(_9069_)
);

AOI21X1 _20089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf1),
    .B(_9041__bF$buf0),
    .C(_9069_),
    .Y(_4520_)
);

NOR2X1 _20090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [28]),
    .B(_9041__bF$buf7),
    .Y(_9070_)
);

AOI21X1 _20091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf1),
    .B(_9041__bF$buf6),
    .C(_9070_),
    .Y(_4521_)
);

NOR2X1 _20092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [29]),
    .B(_9041__bF$buf5),
    .Y(_9071_)
);

AOI21X1 _20093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf0),
    .B(_9041__bF$buf4),
    .C(_9071_),
    .Y(_4522_)
);

NOR2X1 _20094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [30]),
    .B(_9041__bF$buf3),
    .Y(_9072_)
);

AOI21X1 _20095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf0),
    .B(_9041__bF$buf2),
    .C(_9072_),
    .Y(_4524_)
);

NOR2X1 _20096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[12] [31]),
    .B(_9041__bF$buf1),
    .Y(_9073_)
);

AOI21X1 _20097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf1),
    .B(_9041__bF$buf0),
    .C(_9073_),
    .Y(_4525_)
);

NOR2X1 _20098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [9]),
    .B(_6038_),
    .Y(_9074_)
);

NAND2X1 _20099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5435_),
    .B(_9074_),
    .Y(_9075_)
);

INVX8 _20100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9074_),
    .Y(_9076_)
);

OAI21X1 _20101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf8),
    .B(_5434__bF$buf3),
    .C(\datapath.registers.1226[11] [0]),
    .Y(_9077_)
);

OAI21X1 _20102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf4),
    .B(_5429__bF$buf0),
    .C(_9077_),
    .Y(_4469_)
);

OAI21X1 _20103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf7),
    .B(_5434__bF$buf2),
    .C(\datapath.registers.1226[11] [1]),
    .Y(_9078_)
);

OAI21X1 _20104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf3),
    .B(_5438__bF$buf0),
    .C(_9078_),
    .Y(_4480_)
);

OAI21X1 _20105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf6),
    .B(_5434__bF$buf1),
    .C(\datapath.registers.1226[11] [2]),
    .Y(_9079_)
);

OAI21X1 _20106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf2),
    .B(_5440__bF$buf4),
    .C(_9079_),
    .Y(_4491_)
);

OAI21X1 _20107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf5),
    .B(_5434__bF$buf0),
    .C(\datapath.registers.1226[11] [3]),
    .Y(_9080_)
);

OAI21X1 _20108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf1),
    .B(_5442__bF$buf1),
    .C(_9080_),
    .Y(_4494_)
);

OAI21X1 _20109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf4),
    .B(_5434__bF$buf14),
    .C(\datapath.registers.1226[11] [4]),
    .Y(_9081_)
);

OAI21X1 _20110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf0),
    .B(_5444__bF$buf4),
    .C(_9081_),
    .Y(_4495_)
);

OAI21X1 _20111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf3),
    .B(_5434__bF$buf13),
    .C(\datapath.registers.1226[11] [5]),
    .Y(_9082_)
);

OAI21X1 _20112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf4),
    .B(_5446__bF$buf4),
    .C(_9082_),
    .Y(_4496_)
);

OAI21X1 _20113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf2),
    .B(_5434__bF$buf12),
    .C(\datapath.registers.1226[11] [6]),
    .Y(_9083_)
);

OAI21X1 _20114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf3),
    .B(_5448__bF$buf0),
    .C(_9083_),
    .Y(_4497_)
);

OAI21X1 _20115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf1),
    .B(_5434__bF$buf11),
    .C(\datapath.registers.1226[11] [7]),
    .Y(_9084_)
);

OAI21X1 _20116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf2),
    .B(_5450__bF$buf0),
    .C(_9084_),
    .Y(_4498_)
);

OAI21X1 _20117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf0),
    .B(_5434__bF$buf10),
    .C(\datapath.registers.1226[11] [8]),
    .Y(_9085_)
);

OAI21X1 _20118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf1),
    .B(_5452__bF$buf0),
    .C(_9085_),
    .Y(_4499_)
);

OAI21X1 _20119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf8),
    .B(_5434__bF$buf9),
    .C(\datapath.registers.1226[11] [9]),
    .Y(_9086_)
);

OAI21X1 _20120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf0),
    .B(_5454__bF$buf4),
    .C(_9086_),
    .Y(_4500_)
);

OAI21X1 _20121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf7),
    .B(_5434__bF$buf8),
    .C(\datapath.registers.1226[11] [10]),
    .Y(_9087_)
);

OAI21X1 _20122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf4),
    .B(_5456__bF$buf1),
    .C(_9087_),
    .Y(_4470_)
);

OAI21X1 _20123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf6),
    .B(_5434__bF$buf7),
    .C(\datapath.registers.1226[11] [11]),
    .Y(_9088_)
);

OAI21X1 _20124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf3),
    .B(_5458__bF$buf4),
    .C(_9088_),
    .Y(_4471_)
);

OAI21X1 _20125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf5),
    .B(_5434__bF$buf6),
    .C(\datapath.registers.1226[11] [12]),
    .Y(_9089_)
);

OAI21X1 _20126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf2),
    .B(_5460__bF$buf0),
    .C(_9089_),
    .Y(_4472_)
);

OAI21X1 _20127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf4),
    .B(_5434__bF$buf5),
    .C(\datapath.registers.1226[11] [13]),
    .Y(_9090_)
);

OAI21X1 _20128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf1),
    .B(_5462__bF$buf0),
    .C(_9090_),
    .Y(_4473_)
);

OAI21X1 _20129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf3),
    .B(_5434__bF$buf4),
    .C(\datapath.registers.1226[11] [14]),
    .Y(_9091_)
);

OAI21X1 _20130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf0),
    .B(_5464__bF$buf4),
    .C(_9091_),
    .Y(_4474_)
);

OAI21X1 _20131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf2),
    .B(_5434__bF$buf3),
    .C(\datapath.registers.1226[11] [15]),
    .Y(_9092_)
);

OAI21X1 _20132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf4),
    .B(_5466__bF$buf4),
    .C(_9092_),
    .Y(_4475_)
);

OAI21X1 _20133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf1),
    .B(_5434__bF$buf2),
    .C(\datapath.registers.1226[11] [16]),
    .Y(_9093_)
);

OAI21X1 _20134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf3),
    .B(_5468__bF$buf1),
    .C(_9093_),
    .Y(_4476_)
);

OAI21X1 _20135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf0),
    .B(_5434__bF$buf1),
    .C(\datapath.registers.1226[11] [17]),
    .Y(_9094_)
);

OAI21X1 _20136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf2),
    .B(_5470__bF$buf0),
    .C(_9094_),
    .Y(_4477_)
);

OAI21X1 _20137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf8),
    .B(_5434__bF$buf0),
    .C(\datapath.registers.1226[11] [18]),
    .Y(_9095_)
);

OAI21X1 _20138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf1),
    .B(_5472__bF$buf4),
    .C(_9095_),
    .Y(_4478_)
);

OAI21X1 _20139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf7),
    .B(_5434__bF$buf14),
    .C(\datapath.registers.1226[11] [19]),
    .Y(_9096_)
);

OAI21X1 _20140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf0),
    .B(_5474__bF$buf4),
    .C(_9096_),
    .Y(_4479_)
);

OAI21X1 _20141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf6),
    .B(_5434__bF$buf13),
    .C(\datapath.registers.1226[11] [20]),
    .Y(_9097_)
);

OAI21X1 _20142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf4),
    .B(_5476__bF$buf0),
    .C(_9097_),
    .Y(_4481_)
);

OAI21X1 _20143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf5),
    .B(_5434__bF$buf12),
    .C(\datapath.registers.1226[11] [21]),
    .Y(_9098_)
);

OAI21X1 _20144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf3),
    .B(_5478__bF$buf1),
    .C(_9098_),
    .Y(_4482_)
);

OAI21X1 _20145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf4),
    .B(_5434__bF$buf11),
    .C(\datapath.registers.1226[11] [22]),
    .Y(_9099_)
);

OAI21X1 _20146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf2),
    .B(_5480__bF$buf0),
    .C(_9099_),
    .Y(_4483_)
);

OAI21X1 _20147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf3),
    .B(_5434__bF$buf10),
    .C(\datapath.registers.1226[11] [23]),
    .Y(_9100_)
);

OAI21X1 _20148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf1),
    .B(_5482__bF$buf4),
    .C(_9100_),
    .Y(_4484_)
);

OAI21X1 _20149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf2),
    .B(_5434__bF$buf9),
    .C(\datapath.registers.1226[11] [24]),
    .Y(_9101_)
);

OAI21X1 _20150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf0),
    .B(_5484__bF$buf4),
    .C(_9101_),
    .Y(_4485_)
);

OAI21X1 _20151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf1),
    .B(_5434__bF$buf8),
    .C(\datapath.registers.1226[11] [25]),
    .Y(_9102_)
);

OAI21X1 _20152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf4),
    .B(_5486__bF$buf0),
    .C(_9102_),
    .Y(_4486_)
);

OAI21X1 _20153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf0),
    .B(_5434__bF$buf7),
    .C(\datapath.registers.1226[11] [26]),
    .Y(_9103_)
);

OAI21X1 _20154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf3),
    .B(_5488__bF$buf4),
    .C(_9103_),
    .Y(_4487_)
);

OAI21X1 _20155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf8),
    .B(_5434__bF$buf6),
    .C(\datapath.registers.1226[11] [27]),
    .Y(_9104_)
);

OAI21X1 _20156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf2),
    .B(_5490__bF$buf0),
    .C(_9104_),
    .Y(_4488_)
);

OAI21X1 _20157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf7),
    .B(_5434__bF$buf5),
    .C(\datapath.registers.1226[11] [28]),
    .Y(_9105_)
);

OAI21X1 _20158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf1),
    .B(_5492__bF$buf0),
    .C(_9105_),
    .Y(_4489_)
);

OAI21X1 _20159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf6),
    .B(_5434__bF$buf4),
    .C(\datapath.registers.1226[11] [29]),
    .Y(_9106_)
);

OAI21X1 _20160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf0),
    .B(_5494__bF$buf4),
    .C(_9106_),
    .Y(_4490_)
);

OAI21X1 _20161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf5),
    .B(_5434__bF$buf3),
    .C(\datapath.registers.1226[11] [30]),
    .Y(_9107_)
);

OAI21X1 _20162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf4),
    .B(_5496__bF$buf4),
    .C(_9107_),
    .Y(_4492_)
);

OAI21X1 _20163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9076__bF$buf4),
    .B(_5434__bF$buf2),
    .C(\datapath.registers.1226[11] [31]),
    .Y(_9108_)
);

OAI21X1 _20164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075__bF$buf3),
    .B(_5498__bF$buf0),
    .C(_9108_),
    .Y(_4493_)
);

NAND2X1 _20165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9074_),
    .B(_5508_),
    .Y(_9109_)
);

OAI21X1 _20166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf15),
    .B(_9076__bF$buf3),
    .C(\datapath.registers.1226[10] [0]),
    .Y(_9110_)
);

OAI21X1 _20167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf4),
    .B(_9109__bF$buf4),
    .C(_9110_),
    .Y(_4437_)
);

OAI21X1 _20168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf14),
    .B(_9076__bF$buf2),
    .C(\datapath.registers.1226[10] [1]),
    .Y(_9111_)
);

OAI21X1 _20169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf4),
    .B(_9109__bF$buf3),
    .C(_9111_),
    .Y(_4448_)
);

OAI21X1 _20170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf13),
    .B(_9076__bF$buf1),
    .C(\datapath.registers.1226[10] [2]),
    .Y(_9112_)
);

OAI21X1 _20171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf3),
    .B(_9109__bF$buf2),
    .C(_9112_),
    .Y(_4459_)
);

OAI21X1 _20172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf12),
    .B(_9076__bF$buf0),
    .C(\datapath.registers.1226[10] [3]),
    .Y(_9113_)
);

OAI21X1 _20173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf0),
    .B(_9109__bF$buf1),
    .C(_9113_),
    .Y(_4462_)
);

OAI21X1 _20174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf11),
    .B(_9076__bF$buf8),
    .C(\datapath.registers.1226[10] [4]),
    .Y(_9114_)
);

OAI21X1 _20175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf3),
    .B(_9109__bF$buf0),
    .C(_9114_),
    .Y(_4463_)
);

OAI21X1 _20176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf10),
    .B(_9076__bF$buf7),
    .C(\datapath.registers.1226[10] [5]),
    .Y(_9115_)
);

OAI21X1 _20177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf3),
    .B(_9109__bF$buf4),
    .C(_9115_),
    .Y(_4464_)
);

OAI21X1 _20178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf9),
    .B(_9076__bF$buf6),
    .C(\datapath.registers.1226[10] [6]),
    .Y(_9116_)
);

OAI21X1 _20179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf4),
    .B(_9109__bF$buf3),
    .C(_9116_),
    .Y(_4465_)
);

OAI21X1 _20180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf8),
    .B(_9076__bF$buf5),
    .C(\datapath.registers.1226[10] [7]),
    .Y(_9117_)
);

OAI21X1 _20181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf4),
    .B(_9109__bF$buf2),
    .C(_9117_),
    .Y(_4466_)
);

OAI21X1 _20182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf7),
    .B(_9076__bF$buf4),
    .C(\datapath.registers.1226[10] [8]),
    .Y(_9118_)
);

OAI21X1 _20183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf4),
    .B(_9109__bF$buf1),
    .C(_9118_),
    .Y(_4467_)
);

OAI21X1 _20184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf6),
    .B(_9076__bF$buf3),
    .C(\datapath.registers.1226[10] [9]),
    .Y(_9119_)
);

OAI21X1 _20185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf3),
    .B(_9109__bF$buf0),
    .C(_9119_),
    .Y(_4468_)
);

OAI21X1 _20186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf5),
    .B(_9076__bF$buf2),
    .C(\datapath.registers.1226[10] [10]),
    .Y(_9120_)
);

OAI21X1 _20187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf0),
    .B(_9109__bF$buf4),
    .C(_9120_),
    .Y(_4438_)
);

OAI21X1 _20188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf4),
    .B(_9076__bF$buf1),
    .C(\datapath.registers.1226[10] [11]),
    .Y(_9121_)
);

OAI21X1 _20189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf3),
    .B(_9109__bF$buf3),
    .C(_9121_),
    .Y(_4439_)
);

OAI21X1 _20190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf3),
    .B(_9076__bF$buf0),
    .C(\datapath.registers.1226[10] [12]),
    .Y(_9122_)
);

OAI21X1 _20191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf4),
    .B(_9109__bF$buf2),
    .C(_9122_),
    .Y(_4440_)
);

OAI21X1 _20192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf2),
    .B(_9076__bF$buf8),
    .C(\datapath.registers.1226[10] [13]),
    .Y(_9123_)
);

OAI21X1 _20193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf4),
    .B(_9109__bF$buf1),
    .C(_9123_),
    .Y(_4441_)
);

OAI21X1 _20194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf1),
    .B(_9076__bF$buf7),
    .C(\datapath.registers.1226[10] [14]),
    .Y(_9124_)
);

OAI21X1 _20195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf3),
    .B(_9109__bF$buf0),
    .C(_9124_),
    .Y(_4442_)
);

OAI21X1 _20196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf0),
    .B(_9076__bF$buf6),
    .C(\datapath.registers.1226[10] [15]),
    .Y(_9125_)
);

OAI21X1 _20197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf3),
    .B(_9109__bF$buf4),
    .C(_9125_),
    .Y(_4443_)
);

OAI21X1 _20198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf15),
    .B(_9076__bF$buf5),
    .C(\datapath.registers.1226[10] [16]),
    .Y(_9126_)
);

OAI21X1 _20199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf0),
    .B(_9109__bF$buf3),
    .C(_9126_),
    .Y(_4444_)
);

OAI21X1 _20200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf14),
    .B(_9076__bF$buf4),
    .C(\datapath.registers.1226[10] [17]),
    .Y(_9127_)
);

OAI21X1 _20201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf4),
    .B(_9109__bF$buf2),
    .C(_9127_),
    .Y(_4445_)
);

OAI21X1 _20202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf13),
    .B(_9076__bF$buf3),
    .C(\datapath.registers.1226[10] [18]),
    .Y(_9128_)
);

OAI21X1 _20203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf3),
    .B(_9109__bF$buf1),
    .C(_9128_),
    .Y(_4446_)
);

OAI21X1 _20204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf12),
    .B(_9076__bF$buf2),
    .C(\datapath.registers.1226[10] [19]),
    .Y(_9129_)
);

OAI21X1 _20205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf3),
    .B(_9109__bF$buf0),
    .C(_9129_),
    .Y(_4447_)
);

OAI21X1 _20206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf11),
    .B(_9076__bF$buf1),
    .C(\datapath.registers.1226[10] [20]),
    .Y(_9130_)
);

OAI21X1 _20207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf4),
    .B(_9109__bF$buf4),
    .C(_9130_),
    .Y(_4449_)
);

OAI21X1 _20208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf10),
    .B(_9076__bF$buf0),
    .C(\datapath.registers.1226[10] [21]),
    .Y(_9131_)
);

OAI21X1 _20209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf0),
    .B(_9109__bF$buf3),
    .C(_9131_),
    .Y(_4450_)
);

OAI21X1 _20210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf9),
    .B(_9076__bF$buf8),
    .C(\datapath.registers.1226[10] [22]),
    .Y(_9132_)
);

OAI21X1 _20211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf4),
    .B(_9109__bF$buf2),
    .C(_9132_),
    .Y(_4451_)
);

OAI21X1 _20212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf8),
    .B(_9076__bF$buf7),
    .C(\datapath.registers.1226[10] [23]),
    .Y(_9133_)
);

OAI21X1 _20213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf3),
    .B(_9109__bF$buf1),
    .C(_9133_),
    .Y(_4452_)
);

OAI21X1 _20214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf7),
    .B(_9076__bF$buf6),
    .C(\datapath.registers.1226[10] [24]),
    .Y(_9134_)
);

OAI21X1 _20215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf3),
    .B(_9109__bF$buf0),
    .C(_9134_),
    .Y(_4453_)
);

OAI21X1 _20216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf6),
    .B(_9076__bF$buf5),
    .C(\datapath.registers.1226[10] [25]),
    .Y(_9135_)
);

OAI21X1 _20217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486__bF$buf4),
    .B(_9109__bF$buf4),
    .C(_9135_),
    .Y(_4454_)
);

OAI21X1 _20218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf5),
    .B(_9076__bF$buf4),
    .C(\datapath.registers.1226[10] [26]),
    .Y(_9136_)
);

OAI21X1 _20219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf3),
    .B(_9109__bF$buf3),
    .C(_9136_),
    .Y(_4455_)
);

OAI21X1 _20220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf4),
    .B(_9076__bF$buf3),
    .C(\datapath.registers.1226[10] [27]),
    .Y(_9137_)
);

OAI21X1 _20221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf4),
    .B(_9109__bF$buf2),
    .C(_9137_),
    .Y(_4456_)
);

OAI21X1 _20222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf3),
    .B(_9076__bF$buf2),
    .C(\datapath.registers.1226[10] [28]),
    .Y(_9138_)
);

OAI21X1 _20223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf4),
    .B(_9109__bF$buf1),
    .C(_9138_),
    .Y(_4457_)
);

OAI21X1 _20224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf2),
    .B(_9076__bF$buf1),
    .C(\datapath.registers.1226[10] [29]),
    .Y(_9139_)
);

OAI21X1 _20225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf3),
    .B(_9109__bF$buf0),
    .C(_9139_),
    .Y(_4458_)
);

OAI21X1 _20226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf1),
    .B(_9076__bF$buf0),
    .C(\datapath.registers.1226[10] [30]),
    .Y(_9140_)
);

OAI21X1 _20227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf3),
    .B(_9109__bF$buf4),
    .C(_9140_),
    .Y(_4460_)
);

OAI21X1 _20228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf0),
    .B(_9076__bF$buf8),
    .C(\datapath.registers.1226[10] [31]),
    .Y(_9141_)
);

OAI21X1 _20229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf4),
    .B(_9109__bF$buf3),
    .C(_9141_),
    .Y(_4461_)
);

NAND2X1 _20230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9074_),
    .B(_5544_),
    .Y(_9142_)
);

OAI21X1 _20231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf15),
    .B(_9076__bF$buf7),
    .C(\datapath.registers.1226[9] [0]),
    .Y(_9143_)
);

OAI21X1 _20232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf3),
    .B(_9142__bF$buf4),
    .C(_9143_),
    .Y(_5397_)
);

OAI21X1 _20233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf14),
    .B(_9076__bF$buf6),
    .C(\datapath.registers.1226[9] [1]),
    .Y(_9144_)
);

OAI21X1 _20234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf3),
    .B(_9142__bF$buf3),
    .C(_9144_),
    .Y(_5408_)
);

OAI21X1 _20235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf13),
    .B(_9076__bF$buf5),
    .C(\datapath.registers.1226[9] [2]),
    .Y(_9145_)
);

OAI21X1 _20236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf2),
    .B(_9142__bF$buf2),
    .C(_9145_),
    .Y(_5419_)
);

OAI21X1 _20237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf12),
    .B(_9076__bF$buf4),
    .C(\datapath.registers.1226[9] [3]),
    .Y(_9146_)
);

OAI21X1 _20238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf4),
    .B(_9142__bF$buf1),
    .C(_9146_),
    .Y(_5422_)
);

OAI21X1 _20239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf11),
    .B(_9076__bF$buf3),
    .C(\datapath.registers.1226[9] [4]),
    .Y(_9147_)
);

OAI21X1 _20240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf2),
    .B(_9142__bF$buf0),
    .C(_9147_),
    .Y(_5423_)
);

OAI21X1 _20241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf10),
    .B(_9076__bF$buf2),
    .C(\datapath.registers.1226[9] [5]),
    .Y(_9148_)
);

OAI21X1 _20242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf2),
    .B(_9142__bF$buf4),
    .C(_9148_),
    .Y(_5424_)
);

OAI21X1 _20243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf9),
    .B(_9076__bF$buf1),
    .C(\datapath.registers.1226[9] [6]),
    .Y(_9149_)
);

OAI21X1 _20244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf3),
    .B(_9142__bF$buf3),
    .C(_9149_),
    .Y(_5425_)
);

OAI21X1 _20245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf8),
    .B(_9076__bF$buf0),
    .C(\datapath.registers.1226[9] [7]),
    .Y(_9150_)
);

OAI21X1 _20246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf3),
    .B(_9142__bF$buf2),
    .C(_9150_),
    .Y(_5426_)
);

OAI21X1 _20247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf7),
    .B(_9076__bF$buf8),
    .C(\datapath.registers.1226[9] [8]),
    .Y(_9151_)
);

OAI21X1 _20248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf3),
    .B(_9142__bF$buf1),
    .C(_9151_),
    .Y(_5427_)
);

OAI21X1 _20249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf6),
    .B(_9076__bF$buf7),
    .C(\datapath.registers.1226[9] [9]),
    .Y(_9152_)
);

OAI21X1 _20250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf2),
    .B(_9142__bF$buf0),
    .C(_9152_),
    .Y(_5428_)
);

OAI21X1 _20251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf5),
    .B(_9076__bF$buf6),
    .C(\datapath.registers.1226[9] [10]),
    .Y(_9153_)
);

OAI21X1 _20252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf4),
    .B(_9142__bF$buf4),
    .C(_9153_),
    .Y(_5398_)
);

OAI21X1 _20253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf4),
    .B(_9076__bF$buf5),
    .C(\datapath.registers.1226[9] [11]),
    .Y(_9154_)
);

OAI21X1 _20254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf2),
    .B(_9142__bF$buf3),
    .C(_9154_),
    .Y(_5399_)
);

OAI21X1 _20255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf3),
    .B(_9076__bF$buf4),
    .C(\datapath.registers.1226[9] [12]),
    .Y(_9155_)
);

OAI21X1 _20256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf3),
    .B(_9142__bF$buf2),
    .C(_9155_),
    .Y(_5400_)
);

OAI21X1 _20257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf2),
    .B(_9076__bF$buf3),
    .C(\datapath.registers.1226[9] [13]),
    .Y(_9156_)
);

OAI21X1 _20258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf3),
    .B(_9142__bF$buf1),
    .C(_9156_),
    .Y(_5401_)
);

OAI21X1 _20259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf1),
    .B(_9076__bF$buf2),
    .C(\datapath.registers.1226[9] [14]),
    .Y(_9157_)
);

OAI21X1 _20260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf2),
    .B(_9142__bF$buf0),
    .C(_9157_),
    .Y(_5402_)
);

OAI21X1 _20261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf0),
    .B(_9076__bF$buf1),
    .C(\datapath.registers.1226[9] [15]),
    .Y(_9158_)
);

OAI21X1 _20262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf2),
    .B(_9142__bF$buf4),
    .C(_9158_),
    .Y(_5403_)
);

OAI21X1 _20263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf15),
    .B(_9076__bF$buf0),
    .C(\datapath.registers.1226[9] [16]),
    .Y(_9159_)
);

OAI21X1 _20264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf4),
    .B(_9142__bF$buf3),
    .C(_9159_),
    .Y(_5404_)
);

OAI21X1 _20265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf14),
    .B(_9076__bF$buf8),
    .C(\datapath.registers.1226[9] [17]),
    .Y(_9160_)
);

OAI21X1 _20266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf3),
    .B(_9142__bF$buf2),
    .C(_9160_),
    .Y(_5405_)
);

OAI21X1 _20267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf13),
    .B(_9076__bF$buf7),
    .C(\datapath.registers.1226[9] [18]),
    .Y(_9161_)
);

OAI21X1 _20268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf2),
    .B(_9142__bF$buf1),
    .C(_9161_),
    .Y(_5406_)
);

OAI21X1 _20269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf12),
    .B(_9076__bF$buf6),
    .C(\datapath.registers.1226[9] [19]),
    .Y(_9162_)
);

OAI21X1 _20270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf2),
    .B(_9142__bF$buf0),
    .C(_9162_),
    .Y(_5407_)
);

OAI21X1 _20271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf11),
    .B(_9076__bF$buf5),
    .C(\datapath.registers.1226[9] [20]),
    .Y(_9163_)
);

OAI21X1 _20272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf3),
    .B(_9142__bF$buf4),
    .C(_9163_),
    .Y(_5409_)
);

OAI21X1 _20273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf10),
    .B(_9076__bF$buf4),
    .C(\datapath.registers.1226[9] [21]),
    .Y(_9164_)
);

OAI21X1 _20274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf4),
    .B(_9142__bF$buf3),
    .C(_9164_),
    .Y(_5410_)
);

OAI21X1 _20275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf9),
    .B(_9076__bF$buf3),
    .C(\datapath.registers.1226[9] [22]),
    .Y(_9165_)
);

OAI21X1 _20276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf3),
    .B(_9142__bF$buf2),
    .C(_9165_),
    .Y(_5411_)
);

OAI21X1 _20277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf8),
    .B(_9076__bF$buf2),
    .C(\datapath.registers.1226[9] [23]),
    .Y(_9166_)
);

OAI21X1 _20278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf2),
    .B(_9142__bF$buf1),
    .C(_9166_),
    .Y(_5412_)
);

OAI21X1 _20279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf7),
    .B(_9076__bF$buf1),
    .C(\datapath.registers.1226[9] [24]),
    .Y(_9167_)
);

OAI21X1 _20280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf2),
    .B(_9142__bF$buf0),
    .C(_9167_),
    .Y(_5413_)
);

OAI21X1 _20281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf6),
    .B(_9076__bF$buf0),
    .C(\datapath.registers.1226[9] [25]),
    .Y(_9168_)
);

OAI21X1 _20282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486__bF$buf3),
    .B(_9142__bF$buf4),
    .C(_9168_),
    .Y(_5414_)
);

OAI21X1 _20283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf5),
    .B(_9076__bF$buf8),
    .C(\datapath.registers.1226[9] [26]),
    .Y(_9169_)
);

OAI21X1 _20284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf2),
    .B(_9142__bF$buf3),
    .C(_9169_),
    .Y(_5415_)
);

OAI21X1 _20285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf4),
    .B(_9076__bF$buf7),
    .C(\datapath.registers.1226[9] [27]),
    .Y(_9170_)
);

OAI21X1 _20286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf3),
    .B(_9142__bF$buf2),
    .C(_9170_),
    .Y(_5416_)
);

OAI21X1 _20287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf3),
    .B(_9076__bF$buf6),
    .C(\datapath.registers.1226[9] [28]),
    .Y(_9171_)
);

OAI21X1 _20288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf3),
    .B(_9142__bF$buf1),
    .C(_9171_),
    .Y(_5417_)
);

OAI21X1 _20289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf2),
    .B(_9076__bF$buf5),
    .C(\datapath.registers.1226[9] [29]),
    .Y(_9172_)
);

OAI21X1 _20290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf2),
    .B(_9142__bF$buf0),
    .C(_9172_),
    .Y(_5418_)
);

OAI21X1 _20291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf1),
    .B(_9076__bF$buf4),
    .C(\datapath.registers.1226[9] [30]),
    .Y(_9173_)
);

OAI21X1 _20292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf2),
    .B(_9142__bF$buf4),
    .C(_9173_),
    .Y(_5420_)
);

OAI21X1 _20293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf0),
    .B(_9076__bF$buf3),
    .C(\datapath.registers.1226[9] [31]),
    .Y(_9174_)
);

OAI21X1 _20294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf3),
    .B(_9142__bF$buf3),
    .C(_9174_),
    .Y(_5421_)
);

NOR2X1 _20295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf4),
    .B(_9076__bF$buf2),
    .Y(_9175_)
);

NOR2X1 _20296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [0]),
    .B(_9175__bF$buf7),
    .Y(_9176_)
);

AOI21X1 _20297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf2),
    .B(_9175__bF$buf6),
    .C(_9176_),
    .Y(_5365_)
);

NOR2X1 _20298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [1]),
    .B(_9175__bF$buf5),
    .Y(_9177_)
);

AOI21X1 _20299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf2),
    .B(_9175__bF$buf4),
    .C(_9177_),
    .Y(_5376_)
);

NOR2X1 _20300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [2]),
    .B(_9175__bF$buf3),
    .Y(_9178_)
);

AOI21X1 _20301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf1),
    .B(_9175__bF$buf2),
    .C(_9178_),
    .Y(_5387_)
);

NOR2X1 _20302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [3]),
    .B(_9175__bF$buf1),
    .Y(_9179_)
);

AOI21X1 _20303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf3),
    .B(_9175__bF$buf0),
    .C(_9179_),
    .Y(_5390_)
);

NOR2X1 _20304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [4]),
    .B(_9175__bF$buf7),
    .Y(_9180_)
);

AOI21X1 _20305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf1),
    .B(_9175__bF$buf6),
    .C(_9180_),
    .Y(_5391_)
);

NAND2X1 _20306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [5]),
    .B(_9175__bF$buf5),
    .Y(_9181_)
);

OAI21X1 _20307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6406_),
    .B(_9175__bF$buf4),
    .C(_9181_),
    .Y(_5392_)
);

NOR2X1 _20308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [6]),
    .B(_9175__bF$buf3),
    .Y(_9182_)
);

AOI21X1 _20309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf2),
    .B(_9175__bF$buf2),
    .C(_9182_),
    .Y(_5393_)
);

NOR2X1 _20310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [7]),
    .B(_9175__bF$buf1),
    .Y(_9183_)
);

AOI21X1 _20311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf2),
    .B(_9175__bF$buf0),
    .C(_9183_),
    .Y(_5394_)
);

NOR2X1 _20312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [8]),
    .B(_9175__bF$buf7),
    .Y(_9184_)
);

AOI21X1 _20313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf2),
    .B(_9175__bF$buf6),
    .C(_9184_),
    .Y(_5395_)
);

NOR2X1 _20314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [9]),
    .B(_9175__bF$buf5),
    .Y(_9185_)
);

AOI21X1 _20315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf1),
    .B(_9175__bF$buf4),
    .C(_9185_),
    .Y(_5396_)
);

NOR2X1 _20316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [10]),
    .B(_9175__bF$buf3),
    .Y(_9186_)
);

AOI21X1 _20317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf3),
    .B(_9175__bF$buf2),
    .C(_9186_),
    .Y(_5366_)
);

NAND2X1 _20318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [11]),
    .B(_9175__bF$buf1),
    .Y(_9187_)
);

OAI21X1 _20319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8129_),
    .B(_9175__bF$buf0),
    .C(_9187_),
    .Y(_5367_)
);

NAND2X1 _20320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [12]),
    .B(_9175__bF$buf7),
    .Y(_9188_)
);

OAI21X1 _20321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6724_),
    .B(_9175__bF$buf6),
    .C(_9188_),
    .Y(_5368_)
);

NAND2X1 _20322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [13]),
    .B(_9175__bF$buf5),
    .Y(_9189_)
);

OAI21X1 _20323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6770_),
    .B(_9175__bF$buf4),
    .C(_9189_),
    .Y(_5369_)
);

NOR2X1 _20324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [14]),
    .B(_9175__bF$buf3),
    .Y(_9190_)
);

AOI21X1 _20325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf1),
    .B(_9175__bF$buf2),
    .C(_9190_),
    .Y(_5370_)
);

NOR2X1 _20326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [15]),
    .B(_9175__bF$buf1),
    .Y(_9191_)
);

AOI21X1 _20327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf1),
    .B(_9175__bF$buf0),
    .C(_9191_),
    .Y(_5371_)
);

NOR2X1 _20328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [16]),
    .B(_9175__bF$buf7),
    .Y(_9192_)
);

AOI21X1 _20329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf3),
    .B(_9175__bF$buf6),
    .C(_9192_),
    .Y(_5372_)
);

NAND2X1 _20330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [17]),
    .B(_9175__bF$buf5),
    .Y(_9193_)
);

OAI21X1 _20331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6950_),
    .B(_9175__bF$buf4),
    .C(_9193_),
    .Y(_5373_)
);

NAND2X1 _20332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [18]),
    .B(_9175__bF$buf3),
    .Y(_9194_)
);

OAI21X1 _20333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8446_),
    .B(_9175__bF$buf2),
    .C(_9194_),
    .Y(_5374_)
);

NOR2X1 _20334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [19]),
    .B(_9175__bF$buf1),
    .Y(_9195_)
);

AOI21X1 _20335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf1),
    .B(_9175__bF$buf0),
    .C(_9195_),
    .Y(_5375_)
);

NOR2X1 _20336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [20]),
    .B(_9175__bF$buf7),
    .Y(_9196_)
);

AOI21X1 _20337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf2),
    .B(_9175__bF$buf6),
    .C(_9196_),
    .Y(_5377_)
);

NOR2X1 _20338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [21]),
    .B(_9175__bF$buf5),
    .Y(_9197_)
);

AOI21X1 _20339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf3),
    .B(_9175__bF$buf4),
    .C(_9197_),
    .Y(_5378_)
);

NOR2X1 _20340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [22]),
    .B(_9175__bF$buf3),
    .Y(_9198_)
);

AOI21X1 _20341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf2),
    .B(_9175__bF$buf2),
    .C(_9198_),
    .Y(_5379_)
);

NOR2X1 _20342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [23]),
    .B(_9175__bF$buf1),
    .Y(_9199_)
);

AOI21X1 _20343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf1),
    .B(_9175__bF$buf0),
    .C(_9199_),
    .Y(_5380_)
);

NOR2X1 _20344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [24]),
    .B(_9175__bF$buf7),
    .Y(_9200_)
);

AOI21X1 _20345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf1),
    .B(_9175__bF$buf6),
    .C(_9200_),
    .Y(_5381_)
);

NAND2X1 _20346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [25]),
    .B(_9175__bF$buf5),
    .Y(_9201_)
);

OAI21X1 _20347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8754_),
    .B(_9175__bF$buf4),
    .C(_9201_),
    .Y(_5382_)
);

NOR2X1 _20348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [26]),
    .B(_9175__bF$buf3),
    .Y(_9202_)
);

AOI21X1 _20349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf1),
    .B(_9175__bF$buf2),
    .C(_9202_),
    .Y(_5383_)
);

NOR2X1 _20350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [27]),
    .B(_9175__bF$buf1),
    .Y(_9203_)
);

AOI21X1 _20351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf2),
    .B(_9175__bF$buf0),
    .C(_9203_),
    .Y(_5384_)
);

NOR2X1 _20352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [28]),
    .B(_9175__bF$buf7),
    .Y(_9204_)
);

AOI21X1 _20353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf2),
    .B(_9175__bF$buf6),
    .C(_9204_),
    .Y(_5385_)
);

NOR2X1 _20354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [29]),
    .B(_9175__bF$buf5),
    .Y(_9205_)
);

AOI21X1 _20355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf1),
    .B(_9175__bF$buf4),
    .C(_9205_),
    .Y(_5386_)
);

NOR2X1 _20356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [30]),
    .B(_9175__bF$buf3),
    .Y(_9206_)
);

AOI21X1 _20357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf1),
    .B(_9175__bF$buf2),
    .C(_9206_),
    .Y(_5388_)
);

NOR2X1 _20358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[8] [31]),
    .B(_9175__bF$buf1),
    .Y(_9207_)
);

AOI21X1 _20359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf2),
    .B(_9175__bF$buf0),
    .C(_9207_),
    .Y(_5389_)
);

NAND2X1 _20360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5503_),
    .B(_5504_),
    .Y(_9208_)
);

NOR2X1 _20361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5430_),
    .B(_9208_),
    .Y(_9209_)
);

NAND2X1 _20362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5435_),
    .B(_9209_),
    .Y(_9210_)
);

INVX8 _20363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9209_),
    .Y(_9211_)
);

OAI21X1 _20364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf8),
    .B(_5434__bF$buf1),
    .C(\datapath.registers.1226[7] [0]),
    .Y(_9212_)
);

OAI21X1 _20365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf4),
    .B(_5429__bF$buf1),
    .C(_9212_),
    .Y(_5333_)
);

OAI21X1 _20366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf7),
    .B(_5434__bF$buf0),
    .C(\datapath.registers.1226[7] [1]),
    .Y(_9213_)
);

OAI21X1 _20367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf3),
    .B(_5438__bF$buf1),
    .C(_9213_),
    .Y(_5344_)
);

OAI21X1 _20368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf6),
    .B(_5434__bF$buf14),
    .C(\datapath.registers.1226[7] [2]),
    .Y(_9214_)
);

OAI21X1 _20369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf2),
    .B(_5440__bF$buf0),
    .C(_9214_),
    .Y(_5355_)
);

OAI21X1 _20370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf5),
    .B(_5434__bF$buf13),
    .C(\datapath.registers.1226[7] [3]),
    .Y(_9215_)
);

OAI21X1 _20371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf1),
    .B(_5442__bF$buf2),
    .C(_9215_),
    .Y(_5358_)
);

OAI21X1 _20372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf4),
    .B(_5434__bF$buf12),
    .C(\datapath.registers.1226[7] [4]),
    .Y(_9216_)
);

OAI21X1 _20373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf0),
    .B(_5444__bF$buf0),
    .C(_9216_),
    .Y(_5359_)
);

OAI21X1 _20374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf3),
    .B(_5434__bF$buf11),
    .C(\datapath.registers.1226[7] [5]),
    .Y(_9217_)
);

OAI21X1 _20375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf4),
    .B(_5446__bF$buf1),
    .C(_9217_),
    .Y(_5360_)
);

OAI21X1 _20376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf2),
    .B(_5434__bF$buf10),
    .C(\datapath.registers.1226[7] [6]),
    .Y(_9218_)
);

OAI21X1 _20377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf3),
    .B(_5448__bF$buf1),
    .C(_9218_),
    .Y(_5361_)
);

OAI21X1 _20378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf1),
    .B(_5434__bF$buf9),
    .C(\datapath.registers.1226[7] [7]),
    .Y(_9219_)
);

OAI21X1 _20379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf2),
    .B(_5450__bF$buf1),
    .C(_9219_),
    .Y(_5362_)
);

OAI21X1 _20380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf0),
    .B(_5434__bF$buf8),
    .C(\datapath.registers.1226[7] [8]),
    .Y(_9220_)
);

OAI21X1 _20381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf1),
    .B(_5452__bF$buf1),
    .C(_9220_),
    .Y(_5363_)
);

OAI21X1 _20382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf8),
    .B(_5434__bF$buf7),
    .C(\datapath.registers.1226[7] [9]),
    .Y(_9221_)
);

OAI21X1 _20383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf0),
    .B(_5454__bF$buf0),
    .C(_9221_),
    .Y(_5364_)
);

OAI21X1 _20384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf7),
    .B(_5434__bF$buf6),
    .C(\datapath.registers.1226[7] [10]),
    .Y(_9222_)
);

OAI21X1 _20385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf4),
    .B(_5456__bF$buf2),
    .C(_9222_),
    .Y(_5334_)
);

OAI21X1 _20386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf6),
    .B(_5434__bF$buf5),
    .C(\datapath.registers.1226[7] [11]),
    .Y(_9223_)
);

OAI21X1 _20387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf3),
    .B(_5458__bF$buf1),
    .C(_9223_),
    .Y(_5335_)
);

OAI21X1 _20388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf5),
    .B(_5434__bF$buf4),
    .C(\datapath.registers.1226[7] [12]),
    .Y(_9224_)
);

OAI21X1 _20389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf2),
    .B(_5460__bF$buf2),
    .C(_9224_),
    .Y(_5336_)
);

OAI21X1 _20390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf4),
    .B(_5434__bF$buf3),
    .C(\datapath.registers.1226[7] [13]),
    .Y(_9225_)
);

OAI21X1 _20391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf1),
    .B(_5462__bF$buf2),
    .C(_9225_),
    .Y(_5337_)
);

OAI21X1 _20392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf3),
    .B(_5434__bF$buf2),
    .C(\datapath.registers.1226[7] [14]),
    .Y(_9226_)
);

OAI21X1 _20393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf0),
    .B(_5464__bF$buf0),
    .C(_9226_),
    .Y(_5338_)
);

OAI21X1 _20394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf2),
    .B(_5434__bF$buf1),
    .C(\datapath.registers.1226[7] [15]),
    .Y(_9227_)
);

OAI21X1 _20395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf4),
    .B(_5466__bF$buf0),
    .C(_9227_),
    .Y(_5339_)
);

OAI21X1 _20396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf1),
    .B(_5434__bF$buf0),
    .C(\datapath.registers.1226[7] [16]),
    .Y(_9228_)
);

OAI21X1 _20397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf3),
    .B(_5468__bF$buf2),
    .C(_9228_),
    .Y(_5340_)
);

OAI21X1 _20398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf0),
    .B(_5434__bF$buf14),
    .C(\datapath.registers.1226[7] [17]),
    .Y(_9229_)
);

OAI21X1 _20399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf2),
    .B(_5470__bF$buf2),
    .C(_9229_),
    .Y(_5341_)
);

OAI21X1 _20400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf8),
    .B(_5434__bF$buf13),
    .C(\datapath.registers.1226[7] [18]),
    .Y(_9230_)
);

OAI21X1 _20401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf1),
    .B(_5472__bF$buf1),
    .C(_9230_),
    .Y(_5342_)
);

OAI21X1 _20402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf7),
    .B(_5434__bF$buf12),
    .C(\datapath.registers.1226[7] [19]),
    .Y(_9231_)
);

OAI21X1 _20403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf0),
    .B(_5474__bF$buf0),
    .C(_9231_),
    .Y(_5343_)
);

OAI21X1 _20404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf6),
    .B(_5434__bF$buf11),
    .C(\datapath.registers.1226[7] [20]),
    .Y(_9232_)
);

OAI21X1 _20405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf4),
    .B(_5476__bF$buf1),
    .C(_9232_),
    .Y(_5345_)
);

OAI21X1 _20406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf5),
    .B(_5434__bF$buf10),
    .C(\datapath.registers.1226[7] [21]),
    .Y(_9233_)
);

OAI21X1 _20407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf3),
    .B(_5478__bF$buf2),
    .C(_9233_),
    .Y(_5346_)
);

OAI21X1 _20408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf4),
    .B(_5434__bF$buf9),
    .C(\datapath.registers.1226[7] [22]),
    .Y(_9234_)
);

OAI21X1 _20409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf2),
    .B(_5480__bF$buf1),
    .C(_9234_),
    .Y(_5347_)
);

OAI21X1 _20410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf3),
    .B(_5434__bF$buf8),
    .C(\datapath.registers.1226[7] [23]),
    .Y(_9235_)
);

OAI21X1 _20411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf1),
    .B(_5482__bF$buf0),
    .C(_9235_),
    .Y(_5348_)
);

OAI21X1 _20412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf2),
    .B(_5434__bF$buf7),
    .C(\datapath.registers.1226[7] [24]),
    .Y(_9236_)
);

OAI21X1 _20413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf0),
    .B(_5484__bF$buf0),
    .C(_9236_),
    .Y(_5349_)
);

OAI21X1 _20414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf1),
    .B(_5434__bF$buf6),
    .C(\datapath.registers.1226[7] [25]),
    .Y(_9237_)
);

OAI21X1 _20415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf4),
    .B(_5486__bF$buf2),
    .C(_9237_),
    .Y(_5350_)
);

OAI21X1 _20416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf0),
    .B(_5434__bF$buf5),
    .C(\datapath.registers.1226[7] [26]),
    .Y(_9238_)
);

OAI21X1 _20417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf3),
    .B(_5488__bF$buf0),
    .C(_9238_),
    .Y(_5351_)
);

OAI21X1 _20418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf8),
    .B(_5434__bF$buf4),
    .C(\datapath.registers.1226[7] [27]),
    .Y(_9239_)
);

OAI21X1 _20419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf2),
    .B(_5490__bF$buf1),
    .C(_9239_),
    .Y(_5352_)
);

OAI21X1 _20420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf7),
    .B(_5434__bF$buf3),
    .C(\datapath.registers.1226[7] [28]),
    .Y(_9240_)
);

OAI21X1 _20421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf1),
    .B(_5492__bF$buf1),
    .C(_9240_),
    .Y(_5353_)
);

OAI21X1 _20422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf6),
    .B(_5434__bF$buf2),
    .C(\datapath.registers.1226[7] [29]),
    .Y(_9241_)
);

OAI21X1 _20423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf0),
    .B(_5494__bF$buf0),
    .C(_9241_),
    .Y(_5354_)
);

OAI21X1 _20424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf5),
    .B(_5434__bF$buf1),
    .C(\datapath.registers.1226[7] [30]),
    .Y(_9242_)
);

OAI21X1 _20425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf4),
    .B(_5496__bF$buf0),
    .C(_9242_),
    .Y(_5356_)
);

OAI21X1 _20426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf4),
    .B(_5434__bF$buf0),
    .C(\datapath.registers.1226[7] [31]),
    .Y(_9243_)
);

OAI21X1 _20427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210__bF$buf3),
    .B(_5498__bF$buf1),
    .C(_9243_),
    .Y(_5357_)
);

NAND2X1 _20428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9209_),
    .B(_5508_),
    .Y(_9244_)
);

OAI21X1 _20429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf15),
    .B(_9211__bF$buf3),
    .C(\datapath.registers.1226[6] [0]),
    .Y(_9245_)
);

OAI21X1 _20430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf0),
    .B(_9244__bF$buf4),
    .C(_9245_),
    .Y(_5301_)
);

OAI21X1 _20431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf14),
    .B(_9211__bF$buf2),
    .C(\datapath.registers.1226[6] [1]),
    .Y(_9246_)
);

OAI21X1 _20432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf0),
    .B(_9244__bF$buf3),
    .C(_9246_),
    .Y(_5312_)
);

OAI21X1 _20433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf13),
    .B(_9211__bF$buf1),
    .C(\datapath.registers.1226[6] [2]),
    .Y(_9247_)
);

OAI21X1 _20434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf4),
    .B(_9244__bF$buf2),
    .C(_9247_),
    .Y(_5323_)
);

OAI21X1 _20435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf12),
    .B(_9211__bF$buf0),
    .C(\datapath.registers.1226[6] [3]),
    .Y(_9248_)
);

OAI21X1 _20436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf1),
    .B(_9244__bF$buf1),
    .C(_9248_),
    .Y(_5326_)
);

OAI21X1 _20437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf11),
    .B(_9211__bF$buf8),
    .C(\datapath.registers.1226[6] [4]),
    .Y(_9249_)
);

OAI21X1 _20438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf4),
    .B(_9244__bF$buf0),
    .C(_9249_),
    .Y(_5327_)
);

OAI21X1 _20439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf10),
    .B(_9211__bF$buf7),
    .C(\datapath.registers.1226[6] [5]),
    .Y(_9250_)
);

OAI21X1 _20440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf0),
    .B(_9244__bF$buf4),
    .C(_9250_),
    .Y(_5328_)
);

OAI21X1 _20441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf9),
    .B(_9211__bF$buf6),
    .C(\datapath.registers.1226[6] [6]),
    .Y(_9251_)
);

OAI21X1 _20442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf0),
    .B(_9244__bF$buf3),
    .C(_9251_),
    .Y(_5329_)
);

OAI21X1 _20443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf8),
    .B(_9211__bF$buf5),
    .C(\datapath.registers.1226[6] [7]),
    .Y(_9252_)
);

OAI21X1 _20444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf0),
    .B(_9244__bF$buf2),
    .C(_9252_),
    .Y(_5330_)
);

OAI21X1 _20445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf7),
    .B(_9211__bF$buf4),
    .C(\datapath.registers.1226[6] [8]),
    .Y(_9253_)
);

OAI21X1 _20446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf0),
    .B(_9244__bF$buf1),
    .C(_9253_),
    .Y(_5331_)
);

OAI21X1 _20447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf6),
    .B(_9211__bF$buf3),
    .C(\datapath.registers.1226[6] [9]),
    .Y(_9254_)
);

OAI21X1 _20448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf4),
    .B(_9244__bF$buf0),
    .C(_9254_),
    .Y(_5332_)
);

OAI21X1 _20449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf5),
    .B(_9211__bF$buf2),
    .C(\datapath.registers.1226[6] [10]),
    .Y(_9255_)
);

OAI21X1 _20450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf1),
    .B(_9244__bF$buf4),
    .C(_9255_),
    .Y(_5302_)
);

OAI21X1 _20451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf4),
    .B(_9211__bF$buf1),
    .C(\datapath.registers.1226[6] [11]),
    .Y(_9256_)
);

OAI21X1 _20452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf0),
    .B(_9244__bF$buf3),
    .C(_9256_),
    .Y(_5303_)
);

OAI21X1 _20453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf3),
    .B(_9211__bF$buf0),
    .C(\datapath.registers.1226[6] [12]),
    .Y(_9257_)
);

OAI21X1 _20454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf1),
    .B(_9244__bF$buf2),
    .C(_9257_),
    .Y(_5304_)
);

OAI21X1 _20455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf2),
    .B(_9211__bF$buf8),
    .C(\datapath.registers.1226[6] [13]),
    .Y(_9258_)
);

OAI21X1 _20456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf1),
    .B(_9244__bF$buf1),
    .C(_9258_),
    .Y(_5305_)
);

OAI21X1 _20457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf1),
    .B(_9211__bF$buf7),
    .C(\datapath.registers.1226[6] [14]),
    .Y(_9259_)
);

OAI21X1 _20458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf4),
    .B(_9244__bF$buf0),
    .C(_9259_),
    .Y(_5306_)
);

OAI21X1 _20459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf0),
    .B(_9211__bF$buf6),
    .C(\datapath.registers.1226[6] [15]),
    .Y(_9260_)
);

OAI21X1 _20460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf4),
    .B(_9244__bF$buf4),
    .C(_9260_),
    .Y(_5307_)
);

OAI21X1 _20461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf15),
    .B(_9211__bF$buf5),
    .C(\datapath.registers.1226[6] [16]),
    .Y(_9261_)
);

OAI21X1 _20462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf1),
    .B(_9244__bF$buf3),
    .C(_9261_),
    .Y(_5308_)
);

OAI21X1 _20463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf14),
    .B(_9211__bF$buf4),
    .C(\datapath.registers.1226[6] [17]),
    .Y(_9262_)
);

OAI21X1 _20464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf1),
    .B(_9244__bF$buf2),
    .C(_9262_),
    .Y(_5309_)
);

OAI21X1 _20465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf13),
    .B(_9211__bF$buf3),
    .C(\datapath.registers.1226[6] [18]),
    .Y(_9263_)
);

OAI21X1 _20466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf0),
    .B(_9244__bF$buf1),
    .C(_9263_),
    .Y(_5310_)
);

OAI21X1 _20467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf12),
    .B(_9211__bF$buf2),
    .C(\datapath.registers.1226[6] [19]),
    .Y(_9264_)
);

OAI21X1 _20468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf4),
    .B(_9244__bF$buf0),
    .C(_9264_),
    .Y(_5311_)
);

OAI21X1 _20469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf11),
    .B(_9211__bF$buf1),
    .C(\datapath.registers.1226[6] [20]),
    .Y(_9265_)
);

OAI21X1 _20470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf0),
    .B(_9244__bF$buf4),
    .C(_9265_),
    .Y(_5313_)
);

OAI21X1 _20471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf10),
    .B(_9211__bF$buf0),
    .C(\datapath.registers.1226[6] [21]),
    .Y(_9266_)
);

OAI21X1 _20472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf1),
    .B(_9244__bF$buf3),
    .C(_9266_),
    .Y(_5314_)
);

OAI21X1 _20473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf9),
    .B(_9211__bF$buf8),
    .C(\datapath.registers.1226[6] [22]),
    .Y(_9267_)
);

OAI21X1 _20474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf0),
    .B(_9244__bF$buf2),
    .C(_9267_),
    .Y(_5315_)
);

OAI21X1 _20475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf8),
    .B(_9211__bF$buf7),
    .C(\datapath.registers.1226[6] [23]),
    .Y(_9268_)
);

OAI21X1 _20476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf4),
    .B(_9244__bF$buf1),
    .C(_9268_),
    .Y(_5316_)
);

OAI21X1 _20477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf7),
    .B(_9211__bF$buf6),
    .C(\datapath.registers.1226[6] [24]),
    .Y(_9269_)
);

OAI21X1 _20478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf4),
    .B(_9244__bF$buf0),
    .C(_9269_),
    .Y(_5317_)
);

OAI21X1 _20479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf6),
    .B(_9211__bF$buf5),
    .C(\datapath.registers.1226[6] [25]),
    .Y(_9270_)
);

OAI21X1 _20480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486__bF$buf1),
    .B(_9244__bF$buf4),
    .C(_9270_),
    .Y(_5318_)
);

OAI21X1 _20481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf5),
    .B(_9211__bF$buf4),
    .C(\datapath.registers.1226[6] [26]),
    .Y(_9271_)
);

OAI21X1 _20482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf4),
    .B(_9244__bF$buf3),
    .C(_9271_),
    .Y(_5319_)
);

OAI21X1 _20483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf4),
    .B(_9211__bF$buf3),
    .C(\datapath.registers.1226[6] [27]),
    .Y(_9272_)
);

OAI21X1 _20484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf0),
    .B(_9244__bF$buf2),
    .C(_9272_),
    .Y(_5320_)
);

OAI21X1 _20485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf3),
    .B(_9211__bF$buf2),
    .C(\datapath.registers.1226[6] [28]),
    .Y(_9273_)
);

OAI21X1 _20486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf0),
    .B(_9244__bF$buf1),
    .C(_9273_),
    .Y(_5321_)
);

OAI21X1 _20487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf2),
    .B(_9211__bF$buf1),
    .C(\datapath.registers.1226[6] [29]),
    .Y(_9274_)
);

OAI21X1 _20488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf4),
    .B(_9244__bF$buf0),
    .C(_9274_),
    .Y(_5322_)
);

OAI21X1 _20489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf1),
    .B(_9211__bF$buf0),
    .C(\datapath.registers.1226[6] [30]),
    .Y(_9275_)
);

OAI21X1 _20490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf4),
    .B(_9244__bF$buf4),
    .C(_9275_),
    .Y(_5324_)
);

OAI21X1 _20491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf0),
    .B(_9211__bF$buf8),
    .C(\datapath.registers.1226[6] [31]),
    .Y(_9276_)
);

OAI21X1 _20492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf0),
    .B(_9244__bF$buf3),
    .C(_9276_),
    .Y(_5325_)
);

NAND2X1 _20493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5544_),
    .B(_9209_),
    .Y(_9277_)
);

OAI21X1 _20494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf7),
    .B(_5546__bF$buf15),
    .C(\datapath.registers.1226[5] [0]),
    .Y(_9278_)
);

OAI21X1 _20495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf4),
    .B(_9277__bF$buf4),
    .C(_9278_),
    .Y(_5269_)
);

OAI21X1 _20496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf6),
    .B(_5546__bF$buf14),
    .C(\datapath.registers.1226[5] [1]),
    .Y(_9279_)
);

OAI21X1 _20497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf4),
    .B(_9277__bF$buf3),
    .C(_9279_),
    .Y(_5280_)
);

OAI21X1 _20498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf5),
    .B(_5546__bF$buf13),
    .C(\datapath.registers.1226[5] [2]),
    .Y(_9280_)
);

OAI21X1 _20499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf3),
    .B(_9277__bF$buf2),
    .C(_9280_),
    .Y(_5291_)
);

OAI21X1 _20500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf4),
    .B(_5546__bF$buf12),
    .C(\datapath.registers.1226[5] [3]),
    .Y(_9281_)
);

OAI21X1 _20501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf0),
    .B(_9277__bF$buf1),
    .C(_9281_),
    .Y(_5294_)
);

OAI21X1 _20502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf3),
    .B(_5546__bF$buf11),
    .C(\datapath.registers.1226[5] [4]),
    .Y(_9282_)
);

OAI21X1 _20503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf3),
    .B(_9277__bF$buf0),
    .C(_9282_),
    .Y(_5295_)
);

OAI21X1 _20504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf2),
    .B(_5546__bF$buf10),
    .C(\datapath.registers.1226[5] [5]),
    .Y(_9283_)
);

OAI21X1 _20505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf4),
    .B(_9277__bF$buf4),
    .C(_9283_),
    .Y(_5296_)
);

OAI21X1 _20506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf1),
    .B(_5546__bF$buf9),
    .C(\datapath.registers.1226[5] [6]),
    .Y(_9284_)
);

OAI21X1 _20507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf4),
    .B(_9277__bF$buf3),
    .C(_9284_),
    .Y(_5297_)
);

OAI21X1 _20508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf0),
    .B(_5546__bF$buf8),
    .C(\datapath.registers.1226[5] [7]),
    .Y(_9285_)
);

OAI21X1 _20509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf4),
    .B(_9277__bF$buf2),
    .C(_9285_),
    .Y(_5298_)
);

OAI21X1 _20510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf8),
    .B(_5546__bF$buf7),
    .C(\datapath.registers.1226[5] [8]),
    .Y(_9286_)
);

OAI21X1 _20511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf4),
    .B(_9277__bF$buf1),
    .C(_9286_),
    .Y(_5299_)
);

OAI21X1 _20512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf7),
    .B(_5546__bF$buf6),
    .C(\datapath.registers.1226[5] [9]),
    .Y(_9287_)
);

OAI21X1 _20513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf3),
    .B(_9277__bF$buf0),
    .C(_9287_),
    .Y(_5300_)
);

OAI21X1 _20514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf6),
    .B(_5546__bF$buf5),
    .C(\datapath.registers.1226[5] [10]),
    .Y(_9288_)
);

OAI21X1 _20515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf0),
    .B(_9277__bF$buf4),
    .C(_9288_),
    .Y(_5270_)
);

OAI21X1 _20516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf5),
    .B(_5546__bF$buf4),
    .C(\datapath.registers.1226[5] [11]),
    .Y(_9289_)
);

OAI21X1 _20517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf4),
    .B(_9277__bF$buf3),
    .C(_9289_),
    .Y(_5271_)
);

OAI21X1 _20518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf4),
    .B(_5546__bF$buf3),
    .C(\datapath.registers.1226[5] [12]),
    .Y(_9290_)
);

OAI21X1 _20519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf0),
    .B(_9277__bF$buf2),
    .C(_9290_),
    .Y(_5272_)
);

OAI21X1 _20520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf3),
    .B(_5546__bF$buf2),
    .C(\datapath.registers.1226[5] [13]),
    .Y(_9291_)
);

OAI21X1 _20521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf0),
    .B(_9277__bF$buf1),
    .C(_9291_),
    .Y(_5273_)
);

OAI21X1 _20522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf2),
    .B(_5546__bF$buf1),
    .C(\datapath.registers.1226[5] [14]),
    .Y(_9292_)
);

OAI21X1 _20523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf3),
    .B(_9277__bF$buf0),
    .C(_9292_),
    .Y(_5274_)
);

OAI21X1 _20524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf1),
    .B(_5546__bF$buf0),
    .C(\datapath.registers.1226[5] [15]),
    .Y(_9293_)
);

OAI21X1 _20525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf3),
    .B(_9277__bF$buf4),
    .C(_9293_),
    .Y(_5275_)
);

OAI21X1 _20526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf0),
    .B(_5546__bF$buf15),
    .C(\datapath.registers.1226[5] [16]),
    .Y(_9294_)
);

OAI21X1 _20527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf0),
    .B(_9277__bF$buf3),
    .C(_9294_),
    .Y(_5276_)
);

OAI21X1 _20528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf8),
    .B(_5546__bF$buf14),
    .C(\datapath.registers.1226[5] [17]),
    .Y(_9295_)
);

OAI21X1 _20529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf0),
    .B(_9277__bF$buf2),
    .C(_9295_),
    .Y(_5277_)
);

OAI21X1 _20530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf7),
    .B(_5546__bF$buf13),
    .C(\datapath.registers.1226[5] [18]),
    .Y(_9296_)
);

OAI21X1 _20531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf4),
    .B(_9277__bF$buf1),
    .C(_9296_),
    .Y(_5278_)
);

OAI21X1 _20532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf6),
    .B(_5546__bF$buf12),
    .C(\datapath.registers.1226[5] [19]),
    .Y(_9297_)
);

OAI21X1 _20533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf3),
    .B(_9277__bF$buf0),
    .C(_9297_),
    .Y(_5279_)
);

OAI21X1 _20534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf5),
    .B(_5546__bF$buf11),
    .C(\datapath.registers.1226[5] [20]),
    .Y(_9298_)
);

OAI21X1 _20535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf4),
    .B(_9277__bF$buf4),
    .C(_9298_),
    .Y(_5281_)
);

OAI21X1 _20536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf4),
    .B(_5546__bF$buf10),
    .C(\datapath.registers.1226[5] [21]),
    .Y(_9299_)
);

OAI21X1 _20537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf0),
    .B(_9277__bF$buf3),
    .C(_9299_),
    .Y(_5282_)
);

OAI21X1 _20538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf3),
    .B(_5546__bF$buf9),
    .C(\datapath.registers.1226[5] [22]),
    .Y(_9300_)
);

OAI21X1 _20539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf4),
    .B(_9277__bF$buf2),
    .C(_9300_),
    .Y(_5283_)
);

OAI21X1 _20540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf2),
    .B(_5546__bF$buf8),
    .C(\datapath.registers.1226[5] [23]),
    .Y(_9301_)
);

OAI21X1 _20541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf3),
    .B(_9277__bF$buf1),
    .C(_9301_),
    .Y(_5284_)
);

OAI21X1 _20542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf1),
    .B(_5546__bF$buf7),
    .C(\datapath.registers.1226[5] [24]),
    .Y(_9302_)
);

OAI21X1 _20543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf3),
    .B(_9277__bF$buf0),
    .C(_9302_),
    .Y(_5285_)
);

OAI21X1 _20544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf0),
    .B(_5546__bF$buf6),
    .C(\datapath.registers.1226[5] [25]),
    .Y(_9303_)
);

OAI21X1 _20545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486__bF$buf0),
    .B(_9277__bF$buf4),
    .C(_9303_),
    .Y(_5286_)
);

OAI21X1 _20546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf8),
    .B(_5546__bF$buf5),
    .C(\datapath.registers.1226[5] [26]),
    .Y(_9304_)
);

OAI21X1 _20547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf3),
    .B(_9277__bF$buf3),
    .C(_9304_),
    .Y(_5287_)
);

OAI21X1 _20548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf7),
    .B(_5546__bF$buf4),
    .C(\datapath.registers.1226[5] [27]),
    .Y(_9305_)
);

OAI21X1 _20549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf4),
    .B(_9277__bF$buf2),
    .C(_9305_),
    .Y(_5288_)
);

OAI21X1 _20550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf6),
    .B(_5546__bF$buf3),
    .C(\datapath.registers.1226[5] [28]),
    .Y(_9306_)
);

OAI21X1 _20551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf4),
    .B(_9277__bF$buf1),
    .C(_9306_),
    .Y(_5289_)
);

OAI21X1 _20552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf5),
    .B(_5546__bF$buf2),
    .C(\datapath.registers.1226[5] [29]),
    .Y(_9307_)
);

OAI21X1 _20553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf3),
    .B(_9277__bF$buf0),
    .C(_9307_),
    .Y(_5290_)
);

OAI21X1 _20554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf4),
    .B(_5546__bF$buf1),
    .C(\datapath.registers.1226[5] [30]),
    .Y(_9308_)
);

OAI21X1 _20555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf3),
    .B(_9277__bF$buf4),
    .C(_9308_),
    .Y(_5292_)
);

OAI21X1 _20556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9211__bF$buf3),
    .B(_5546__bF$buf0),
    .C(\datapath.registers.1226[5] [31]),
    .Y(_9309_)
);

OAI21X1 _20557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf4),
    .B(_9277__bF$buf3),
    .C(_9309_),
    .Y(_5293_)
);

NOR2X1 _20558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5579__bF$buf3),
    .B(_9211__bF$buf2),
    .Y(_9310_)
);

NOR2X1 _20559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [0]),
    .B(_9310__bF$buf7),
    .Y(_9311_)
);

AOI21X1 _20560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf3),
    .B(_9310__bF$buf6),
    .C(_9311_),
    .Y(_5237_)
);

NOR2X1 _20561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [1]),
    .B(_9310__bF$buf5),
    .Y(_9312_)
);

AOI21X1 _20562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf3),
    .B(_9310__bF$buf4),
    .C(_9312_),
    .Y(_5248_)
);

NOR2X1 _20563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [2]),
    .B(_9310__bF$buf3),
    .Y(_9313_)
);

AOI21X1 _20564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf2),
    .B(_9310__bF$buf2),
    .C(_9313_),
    .Y(_5259_)
);

NOR2X1 _20565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [3]),
    .B(_9310__bF$buf1),
    .Y(_9314_)
);

AOI21X1 _20566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf4),
    .B(_9310__bF$buf0),
    .C(_9314_),
    .Y(_5262_)
);

NOR2X1 _20567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [4]),
    .B(_9310__bF$buf7),
    .Y(_9315_)
);

AOI21X1 _20568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf2),
    .B(_9310__bF$buf6),
    .C(_9315_),
    .Y(_5263_)
);

NOR2X1 _20569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [5]),
    .B(_9310__bF$buf5),
    .Y(_9316_)
);

AOI21X1 _20570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf3),
    .B(_9310__bF$buf4),
    .C(_9316_),
    .Y(_5264_)
);

NOR2X1 _20571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [6]),
    .B(_9310__bF$buf3),
    .Y(_9317_)
);

AOI21X1 _20572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf3),
    .B(_9310__bF$buf2),
    .C(_9317_),
    .Y(_5265_)
);

NOR2X1 _20573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [7]),
    .B(_9310__bF$buf1),
    .Y(_9318_)
);

AOI21X1 _20574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf3),
    .B(_9310__bF$buf0),
    .C(_9318_),
    .Y(_5266_)
);

NOR2X1 _20575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [8]),
    .B(_9310__bF$buf7),
    .Y(_9319_)
);

AOI21X1 _20576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf3),
    .B(_9310__bF$buf6),
    .C(_9319_),
    .Y(_5267_)
);

NOR2X1 _20577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [9]),
    .B(_9310__bF$buf5),
    .Y(_9320_)
);

AOI21X1 _20578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf2),
    .B(_9310__bF$buf4),
    .C(_9320_),
    .Y(_5268_)
);

NOR2X1 _20579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [10]),
    .B(_9310__bF$buf3),
    .Y(_9321_)
);

AOI21X1 _20580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf4),
    .B(_9310__bF$buf2),
    .C(_9321_),
    .Y(_5238_)
);

NOR2X1 _20581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [11]),
    .B(_9310__bF$buf1),
    .Y(_9322_)
);

AOI21X1 _20582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf3),
    .B(_9310__bF$buf0),
    .C(_9322_),
    .Y(_5239_)
);

NOR2X1 _20583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [12]),
    .B(_9310__bF$buf7),
    .Y(_9323_)
);

AOI21X1 _20584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf4),
    .B(_9310__bF$buf6),
    .C(_9323_),
    .Y(_5240_)
);

NOR2X1 _20585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [13]),
    .B(_9310__bF$buf5),
    .Y(_9324_)
);

AOI21X1 _20586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf4),
    .B(_9310__bF$buf4),
    .C(_9324_),
    .Y(_5241_)
);

NOR2X1 _20587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [14]),
    .B(_9310__bF$buf3),
    .Y(_9325_)
);

AOI21X1 _20588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf2),
    .B(_9310__bF$buf2),
    .C(_9325_),
    .Y(_5242_)
);

NOR2X1 _20589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [15]),
    .B(_9310__bF$buf1),
    .Y(_9326_)
);

AOI21X1 _20590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf2),
    .B(_9310__bF$buf0),
    .C(_9326_),
    .Y(_5243_)
);

NOR2X1 _20591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [16]),
    .B(_9310__bF$buf7),
    .Y(_9327_)
);

AOI21X1 _20592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf4),
    .B(_9310__bF$buf6),
    .C(_9327_),
    .Y(_5244_)
);

NOR2X1 _20593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [17]),
    .B(_9310__bF$buf5),
    .Y(_9328_)
);

AOI21X1 _20594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf4),
    .B(_9310__bF$buf4),
    .C(_9328_),
    .Y(_5245_)
);

NOR2X1 _20595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [18]),
    .B(_9310__bF$buf3),
    .Y(_9329_)
);

AOI21X1 _20596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf3),
    .B(_9310__bF$buf2),
    .C(_9329_),
    .Y(_5246_)
);

NOR2X1 _20597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [19]),
    .B(_9310__bF$buf1),
    .Y(_9330_)
);

AOI21X1 _20598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf2),
    .B(_9310__bF$buf0),
    .C(_9330_),
    .Y(_5247_)
);

NOR2X1 _20599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [20]),
    .B(_9310__bF$buf7),
    .Y(_9331_)
);

AOI21X1 _20600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf3),
    .B(_9310__bF$buf6),
    .C(_9331_),
    .Y(_5249_)
);

NOR2X1 _20601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [21]),
    .B(_9310__bF$buf5),
    .Y(_9332_)
);

AOI21X1 _20602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf4),
    .B(_9310__bF$buf4),
    .C(_9332_),
    .Y(_5250_)
);

NOR2X1 _20603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [22]),
    .B(_9310__bF$buf3),
    .Y(_9333_)
);

AOI21X1 _20604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf3),
    .B(_9310__bF$buf2),
    .C(_9333_),
    .Y(_5251_)
);

NOR2X1 _20605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [23]),
    .B(_9310__bF$buf1),
    .Y(_9334_)
);

AOI21X1 _20606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf2),
    .B(_9310__bF$buf0),
    .C(_9334_),
    .Y(_5252_)
);

NOR2X1 _20607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [24]),
    .B(_9310__bF$buf7),
    .Y(_9335_)
);

AOI21X1 _20608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf2),
    .B(_9310__bF$buf6),
    .C(_9335_),
    .Y(_5253_)
);

NOR2X1 _20609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [25]),
    .B(_9310__bF$buf5),
    .Y(_9336_)
);

AOI21X1 _20610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486__bF$buf4),
    .B(_9310__bF$buf4),
    .C(_9336_),
    .Y(_5254_)
);

NOR2X1 _20611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [26]),
    .B(_9310__bF$buf3),
    .Y(_9337_)
);

AOI21X1 _20612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf2),
    .B(_9310__bF$buf2),
    .C(_9337_),
    .Y(_5255_)
);

NOR2X1 _20613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [27]),
    .B(_9310__bF$buf1),
    .Y(_9338_)
);

AOI21X1 _20614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf3),
    .B(_9310__bF$buf0),
    .C(_9338_),
    .Y(_5256_)
);

NOR2X1 _20615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [28]),
    .B(_9310__bF$buf7),
    .Y(_9339_)
);

AOI21X1 _20616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf3),
    .B(_9310__bF$buf6),
    .C(_9339_),
    .Y(_5257_)
);

NOR2X1 _20617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [29]),
    .B(_9310__bF$buf5),
    .Y(_9340_)
);

AOI21X1 _20618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf2),
    .B(_9310__bF$buf4),
    .C(_9340_),
    .Y(_5258_)
);

NOR2X1 _20619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [30]),
    .B(_9310__bF$buf3),
    .Y(_9341_)
);

AOI21X1 _20620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf2),
    .B(_9310__bF$buf2),
    .C(_9341_),
    .Y(_5260_)
);

NOR2X1 _20621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[4] [31]),
    .B(_9310__bF$buf1),
    .Y(_9342_)
);

AOI21X1 _20622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf3),
    .B(_9310__bF$buf0),
    .C(_9342_),
    .Y(_5261_)
);

NOR2X1 _20623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5434__bF$buf14),
    .B(_5505__bF$buf6),
    .Y(_9343_)
);

NAND2X1 _20624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [0]),
    .B(_9343__bF$buf7),
    .Y(_9344_)
);

OAI21X1 _20625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6155_),
    .B(_9343__bF$buf6),
    .C(_9344_),
    .Y(_5205_)
);

NAND2X1 _20626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [1]),
    .B(_9343__bF$buf5),
    .Y(_9345_)
);

OAI21X1 _20627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6213_),
    .B(_9343__bF$buf4),
    .C(_9345_),
    .Y(_5216_)
);

NAND2X1 _20628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [2]),
    .B(_9343__bF$buf3),
    .Y(_9346_)
);

OAI21X1 _20629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6283_),
    .B(_9343__bF$buf2),
    .C(_9346_),
    .Y(_5227_)
);

NOR2X1 _20630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [3]),
    .B(_9343__bF$buf1),
    .Y(_9347_)
);

AOI21X1 _20631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf3),
    .B(_9343__bF$buf0),
    .C(_9347_),
    .Y(_5230_)
);

NOR2X1 _20632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [4]),
    .B(_9343__bF$buf7),
    .Y(_9348_)
);

AOI21X1 _20633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf1),
    .B(_9343__bF$buf6),
    .C(_9348_),
    .Y(_5231_)
);

NOR2X1 _20634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [5]),
    .B(_9343__bF$buf5),
    .Y(_9349_)
);

AOI21X1 _20635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf2),
    .B(_9343__bF$buf4),
    .C(_9349_),
    .Y(_5232_)
);

NAND2X1 _20636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [6]),
    .B(_9343__bF$buf3),
    .Y(_9350_)
);

OAI21X1 _20637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7893_),
    .B(_9343__bF$buf2),
    .C(_9350_),
    .Y(_5233_)
);

NAND2X1 _20638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [7]),
    .B(_9343__bF$buf1),
    .Y(_9351_)
);

OAI21X1 _20639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7939_),
    .B(_9343__bF$buf0),
    .C(_9351_),
    .Y(_5234_)
);

NAND2X1 _20640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [8]),
    .B(_9343__bF$buf7),
    .Y(_9352_)
);

OAI21X1 _20641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8009_),
    .B(_9343__bF$buf6),
    .C(_9352_),
    .Y(_5235_)
);

NOR2X1 _20642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [9]),
    .B(_9343__bF$buf5),
    .Y(_9353_)
);

AOI21X1 _20643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf1),
    .B(_9343__bF$buf4),
    .C(_9353_),
    .Y(_5236_)
);

NOR2X1 _20644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [10]),
    .B(_9343__bF$buf3),
    .Y(_9354_)
);

AOI21X1 _20645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf3),
    .B(_9343__bF$buf2),
    .C(_9354_),
    .Y(_5206_)
);

NOR2X1 _20646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [11]),
    .B(_9343__bF$buf1),
    .Y(_9355_)
);

AOI21X1 _20647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf2),
    .B(_9343__bF$buf0),
    .C(_9355_),
    .Y(_5207_)
);

NOR2X1 _20648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [12]),
    .B(_9343__bF$buf7),
    .Y(_9356_)
);

AOI21X1 _20649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf3),
    .B(_9343__bF$buf6),
    .C(_9356_),
    .Y(_5208_)
);

NOR2X1 _20650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [13]),
    .B(_9343__bF$buf5),
    .Y(_9357_)
);

AOI21X1 _20651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf3),
    .B(_9343__bF$buf4),
    .C(_9357_),
    .Y(_5209_)
);

NAND2X1 _20652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [14]),
    .B(_9343__bF$buf3),
    .Y(_9358_)
);

OAI21X1 _20653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8280_),
    .B(_9343__bF$buf2),
    .C(_9358_),
    .Y(_5210_)
);

NOR2X1 _20654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [15]),
    .B(_9343__bF$buf1),
    .Y(_9359_)
);

AOI21X1 _20655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf1),
    .B(_9343__bF$buf0),
    .C(_9359_),
    .Y(_5211_)
);

NOR2X1 _20656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [16]),
    .B(_9343__bF$buf7),
    .Y(_9360_)
);

AOI21X1 _20657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf3),
    .B(_9343__bF$buf6),
    .C(_9360_),
    .Y(_5212_)
);

NOR2X1 _20658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [17]),
    .B(_9343__bF$buf5),
    .Y(_9361_)
);

AOI21X1 _20659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf3),
    .B(_9343__bF$buf4),
    .C(_9361_),
    .Y(_5213_)
);

NOR2X1 _20660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [18]),
    .B(_9343__bF$buf3),
    .Y(_9362_)
);

AOI21X1 _20661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf2),
    .B(_9343__bF$buf2),
    .C(_9362_),
    .Y(_5214_)
);

NAND2X1 _20662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [19]),
    .B(_9343__bF$buf1),
    .Y(_9363_)
);

OAI21X1 _20663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7052_),
    .B(_9343__bF$buf0),
    .C(_9363_),
    .Y(_5215_)
);

NOR2X1 _20664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [20]),
    .B(_9343__bF$buf7),
    .Y(_9364_)
);

AOI21X1 _20665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf2),
    .B(_9343__bF$buf6),
    .C(_9364_),
    .Y(_5217_)
);

NOR2X1 _20666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [21]),
    .B(_9343__bF$buf5),
    .Y(_9365_)
);

AOI21X1 _20667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf3),
    .B(_9343__bF$buf4),
    .C(_9365_),
    .Y(_5218_)
);

NOR2X1 _20668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [22]),
    .B(_9343__bF$buf3),
    .Y(_9366_)
);

AOI21X1 _20669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf2),
    .B(_9343__bF$buf2),
    .C(_9366_),
    .Y(_5219_)
);

NOR2X1 _20670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [23]),
    .B(_9343__bF$buf1),
    .Y(_9367_)
);

AOI21X1 _20671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf1),
    .B(_9343__bF$buf0),
    .C(_9367_),
    .Y(_5220_)
);

NAND2X1 _20672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [24]),
    .B(_9343__bF$buf7),
    .Y(_9368_)
);

OAI21X1 _20673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8721_),
    .B(_9343__bF$buf6),
    .C(_9368_),
    .Y(_5221_)
);

NAND2X1 _20674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [25]),
    .B(_9343__bF$buf5),
    .Y(_9369_)
);

OAI21X1 _20675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7293_),
    .B(_9343__bF$buf4),
    .C(_9369_),
    .Y(_5222_)
);

NOR2X1 _20676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [26]),
    .B(_9343__bF$buf3),
    .Y(_9370_)
);

AOI21X1 _20677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf1),
    .B(_9343__bF$buf2),
    .C(_9370_),
    .Y(_5223_)
);

NAND2X1 _20678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [27]),
    .B(_9343__bF$buf1),
    .Y(_9371_)
);

OAI21X1 _20679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7395_),
    .B(_9343__bF$buf0),
    .C(_9371_),
    .Y(_5224_)
);

NAND2X1 _20680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [28]),
    .B(_9343__bF$buf7),
    .Y(_9372_)
);

OAI21X1 _20681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7465_),
    .B(_9343__bF$buf6),
    .C(_9372_),
    .Y(_5225_)
);

NAND2X1 _20682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [29]),
    .B(_9343__bF$buf5),
    .Y(_9373_)
);

OAI21X1 _20683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8944_),
    .B(_9343__bF$buf4),
    .C(_9373_),
    .Y(_5226_)
);

NAND2X1 _20684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.rd [30]),
    .B(_9343__bF$buf3),
    .Y(_9374_)
);

OAI21X1 _20685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7554_),
    .B(_9343__bF$buf2),
    .C(_9374_),
    .Y(_5228_)
);

NOR2X1 _20686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[3] [31]),
    .B(_9343__bF$buf1),
    .Y(_9375_)
);

AOI21X1 _20687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf2),
    .B(_9343__bF$buf0),
    .C(_9375_),
    .Y(_5229_)
);

INVX1 _20688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5505__bF$buf5),
    .Y(_9376_)
);

NAND2X1 _20689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9376_),
    .B(_5508_),
    .Y(_9377_)
);

OAI21X1 _20690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf15),
    .B(_5505__bF$buf4),
    .C(\datapath.registers.1226[2] [0]),
    .Y(_9378_)
);

OAI21X1 _20691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf2),
    .B(_9377__bF$buf4),
    .C(_9378_),
    .Y(_5109_)
);

OAI21X1 _20692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf14),
    .B(_5505__bF$buf3),
    .C(\datapath.registers.1226[2] [1]),
    .Y(_9379_)
);

OAI21X1 _20693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf2),
    .B(_9377__bF$buf3),
    .C(_9379_),
    .Y(_5120_)
);

OAI21X1 _20694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf13),
    .B(_5505__bF$buf2),
    .C(\datapath.registers.1226[2] [2]),
    .Y(_9380_)
);

OAI21X1 _20695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf1),
    .B(_9377__bF$buf2),
    .C(_9380_),
    .Y(_5131_)
);

OAI21X1 _20696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf12),
    .B(_5505__bF$buf1),
    .C(\datapath.registers.1226[2] [3]),
    .Y(_9381_)
);

OAI21X1 _20697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf2),
    .B(_9377__bF$buf1),
    .C(_9381_),
    .Y(_5134_)
);

OAI21X1 _20698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf11),
    .B(_5505__bF$buf0),
    .C(\datapath.registers.1226[2] [4]),
    .Y(_9382_)
);

OAI21X1 _20699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf0),
    .B(_9377__bF$buf0),
    .C(_9382_),
    .Y(_5135_)
);

OAI21X1 _20700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf10),
    .B(_5505__bF$buf7),
    .C(\datapath.registers.1226[2] [5]),
    .Y(_9383_)
);

OAI21X1 _20701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf1),
    .B(_9377__bF$buf4),
    .C(_9383_),
    .Y(_5136_)
);

OAI21X1 _20702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf9),
    .B(_5505__bF$buf6),
    .C(\datapath.registers.1226[2] [6]),
    .Y(_9384_)
);

OAI21X1 _20703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf2),
    .B(_9377__bF$buf3),
    .C(_9384_),
    .Y(_5137_)
);

OAI21X1 _20704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf8),
    .B(_5505__bF$buf5),
    .C(\datapath.registers.1226[2] [7]),
    .Y(_9385_)
);

OAI21X1 _20705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf2),
    .B(_9377__bF$buf2),
    .C(_9385_),
    .Y(_5138_)
);

OAI21X1 _20706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf7),
    .B(_5505__bF$buf4),
    .C(\datapath.registers.1226[2] [8]),
    .Y(_9386_)
);

OAI21X1 _20707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf2),
    .B(_9377__bF$buf1),
    .C(_9386_),
    .Y(_5139_)
);

OAI21X1 _20708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf6),
    .B(_5505__bF$buf3),
    .C(\datapath.registers.1226[2] [9]),
    .Y(_9387_)
);

OAI21X1 _20709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf0),
    .B(_9377__bF$buf0),
    .C(_9387_),
    .Y(_5140_)
);

OAI21X1 _20710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf5),
    .B(_5505__bF$buf2),
    .C(\datapath.registers.1226[2] [10]),
    .Y(_9388_)
);

OAI21X1 _20711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf2),
    .B(_9377__bF$buf4),
    .C(_9388_),
    .Y(_5110_)
);

OAI21X1 _20712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf4),
    .B(_5505__bF$buf1),
    .C(\datapath.registers.1226[2] [11]),
    .Y(_9389_)
);

OAI21X1 _20713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf1),
    .B(_9377__bF$buf3),
    .C(_9389_),
    .Y(_5111_)
);

OAI21X1 _20714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf3),
    .B(_5505__bF$buf0),
    .C(\datapath.registers.1226[2] [12]),
    .Y(_9390_)
);

OAI21X1 _20715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf2),
    .B(_9377__bF$buf2),
    .C(_9390_),
    .Y(_5112_)
);

OAI21X1 _20716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf2),
    .B(_5505__bF$buf7),
    .C(\datapath.registers.1226[2] [13]),
    .Y(_9391_)
);

OAI21X1 _20717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf2),
    .B(_9377__bF$buf1),
    .C(_9391_),
    .Y(_5113_)
);

OAI21X1 _20718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf1),
    .B(_5505__bF$buf6),
    .C(\datapath.registers.1226[2] [14]),
    .Y(_9392_)
);

OAI21X1 _20719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf1),
    .B(_9377__bF$buf0),
    .C(_9392_),
    .Y(_5114_)
);

OAI21X1 _20720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf0),
    .B(_5505__bF$buf5),
    .C(\datapath.registers.1226[2] [15]),
    .Y(_9393_)
);

OAI21X1 _20721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf0),
    .B(_9377__bF$buf4),
    .C(_9393_),
    .Y(_5115_)
);

OAI21X1 _20722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf15),
    .B(_5505__bF$buf4),
    .C(\datapath.registers.1226[2] [16]),
    .Y(_9394_)
);

OAI21X1 _20723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf2),
    .B(_9377__bF$buf3),
    .C(_9394_),
    .Y(_5116_)
);

OAI21X1 _20724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf14),
    .B(_5505__bF$buf3),
    .C(\datapath.registers.1226[2] [17]),
    .Y(_9395_)
);

OAI21X1 _20725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf2),
    .B(_9377__bF$buf2),
    .C(_9395_),
    .Y(_5117_)
);

OAI21X1 _20726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf13),
    .B(_5505__bF$buf2),
    .C(\datapath.registers.1226[2] [18]),
    .Y(_9396_)
);

OAI21X1 _20727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf1),
    .B(_9377__bF$buf1),
    .C(_9396_),
    .Y(_5118_)
);

OAI21X1 _20728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf12),
    .B(_5505__bF$buf1),
    .C(\datapath.registers.1226[2] [19]),
    .Y(_9397_)
);

OAI21X1 _20729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf1),
    .B(_9377__bF$buf0),
    .C(_9397_),
    .Y(_5119_)
);

OAI21X1 _20730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf11),
    .B(_5505__bF$buf0),
    .C(\datapath.registers.1226[2] [20]),
    .Y(_9398_)
);

OAI21X1 _20731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf1),
    .B(_9377__bF$buf4),
    .C(_9398_),
    .Y(_5121_)
);

OAI21X1 _20732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf10),
    .B(_5505__bF$buf7),
    .C(\datapath.registers.1226[2] [21]),
    .Y(_9399_)
);

OAI21X1 _20733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf2),
    .B(_9377__bF$buf3),
    .C(_9399_),
    .Y(_5122_)
);

OAI21X1 _20734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf9),
    .B(_5505__bF$buf6),
    .C(\datapath.registers.1226[2] [22]),
    .Y(_9400_)
);

OAI21X1 _20735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf1),
    .B(_9377__bF$buf2),
    .C(_9400_),
    .Y(_5123_)
);

OAI21X1 _20736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf8),
    .B(_5505__bF$buf5),
    .C(\datapath.registers.1226[2] [23]),
    .Y(_9401_)
);

OAI21X1 _20737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf0),
    .B(_9377__bF$buf1),
    .C(_9401_),
    .Y(_5124_)
);

OAI21X1 _20738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf7),
    .B(_5505__bF$buf4),
    .C(\datapath.registers.1226[2] [24]),
    .Y(_9402_)
);

OAI21X1 _20739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf1),
    .B(_9377__bF$buf0),
    .C(_9402_),
    .Y(_5125_)
);

OAI21X1 _20740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf6),
    .B(_5505__bF$buf3),
    .C(\datapath.registers.1226[2] [25]),
    .Y(_9403_)
);

OAI21X1 _20741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486__bF$buf3),
    .B(_9377__bF$buf4),
    .C(_9403_),
    .Y(_5126_)
);

OAI21X1 _20742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf5),
    .B(_5505__bF$buf2),
    .C(\datapath.registers.1226[2] [26]),
    .Y(_9404_)
);

OAI21X1 _20743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf0),
    .B(_9377__bF$buf3),
    .C(_9404_),
    .Y(_5127_)
);

OAI21X1 _20744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf4),
    .B(_5505__bF$buf1),
    .C(\datapath.registers.1226[2] [27]),
    .Y(_9405_)
);

OAI21X1 _20745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf2),
    .B(_9377__bF$buf2),
    .C(_9405_),
    .Y(_5128_)
);

OAI21X1 _20746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf3),
    .B(_5505__bF$buf0),
    .C(\datapath.registers.1226[2] [28]),
    .Y(_9406_)
);

OAI21X1 _20747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf2),
    .B(_9377__bF$buf1),
    .C(_9406_),
    .Y(_5129_)
);

OAI21X1 _20748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf2),
    .B(_5505__bF$buf7),
    .C(\datapath.registers.1226[2] [29]),
    .Y(_9407_)
);

OAI21X1 _20749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf1),
    .B(_9377__bF$buf0),
    .C(_9407_),
    .Y(_5130_)
);

OAI21X1 _20750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf1),
    .B(_5505__bF$buf6),
    .C(\datapath.registers.1226[2] [30]),
    .Y(_9408_)
);

OAI21X1 _20751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf1),
    .B(_9377__bF$buf4),
    .C(_9408_),
    .Y(_5132_)
);

OAI21X1 _20752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510__bF$buf0),
    .B(_5505__bF$buf5),
    .C(\datapath.registers.1226[2] [31]),
    .Y(_9409_)
);

OAI21X1 _20753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf1),
    .B(_9377__bF$buf3),
    .C(_9409_),
    .Y(_5133_)
);

NAND2X1 _20754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9376_),
    .B(_5544_),
    .Y(_9410_)
);

OAI21X1 _20755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf15),
    .B(_5505__bF$buf4),
    .C(\datapath.registers.1226[1] [0]),
    .Y(_9411_)
);

OAI21X1 _20756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5429__bF$buf1),
    .B(_9410__bF$buf4),
    .C(_9411_),
    .Y(_4757_)
);

OAI21X1 _20757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf14),
    .B(_5505__bF$buf3),
    .C(\datapath.registers.1226[1] [1]),
    .Y(_9412_)
);

OAI21X1 _20758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438__bF$buf1),
    .B(_9410__bF$buf3),
    .C(_9412_),
    .Y(_4768_)
);

OAI21X1 _20759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf13),
    .B(_5505__bF$buf2),
    .C(\datapath.registers.1226[1] [2]),
    .Y(_9413_)
);

OAI21X1 _20760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440__bF$buf0),
    .B(_9410__bF$buf2),
    .C(_9413_),
    .Y(_4779_)
);

OAI21X1 _20761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf12),
    .B(_5505__bF$buf1),
    .C(\datapath.registers.1226[1] [3]),
    .Y(_9414_)
);

OAI21X1 _20762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442__bF$buf1),
    .B(_9410__bF$buf1),
    .C(_9414_),
    .Y(_4782_)
);

OAI21X1 _20763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf11),
    .B(_5505__bF$buf0),
    .C(\datapath.registers.1226[1] [4]),
    .Y(_9415_)
);

OAI21X1 _20764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444__bF$buf4),
    .B(_9410__bF$buf0),
    .C(_9415_),
    .Y(_4783_)
);

OAI21X1 _20765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf10),
    .B(_5505__bF$buf7),
    .C(\datapath.registers.1226[1] [5]),
    .Y(_9416_)
);

OAI21X1 _20766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446__bF$buf0),
    .B(_9410__bF$buf4),
    .C(_9416_),
    .Y(_4784_)
);

OAI21X1 _20767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf9),
    .B(_5505__bF$buf6),
    .C(\datapath.registers.1226[1] [6]),
    .Y(_9417_)
);

OAI21X1 _20768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448__bF$buf1),
    .B(_9410__bF$buf3),
    .C(_9417_),
    .Y(_4785_)
);

OAI21X1 _20769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf8),
    .B(_5505__bF$buf5),
    .C(\datapath.registers.1226[1] [7]),
    .Y(_9418_)
);

OAI21X1 _20770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5450__bF$buf1),
    .B(_9410__bF$buf2),
    .C(_9418_),
    .Y(_4786_)
);

OAI21X1 _20771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf7),
    .B(_5505__bF$buf4),
    .C(\datapath.registers.1226[1] [8]),
    .Y(_9419_)
);

OAI21X1 _20772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452__bF$buf1),
    .B(_9410__bF$buf1),
    .C(_9419_),
    .Y(_4787_)
);

OAI21X1 _20773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf6),
    .B(_5505__bF$buf3),
    .C(\datapath.registers.1226[1] [9]),
    .Y(_9420_)
);

OAI21X1 _20774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5454__bF$buf4),
    .B(_9410__bF$buf0),
    .C(_9420_),
    .Y(_4788_)
);

OAI21X1 _20775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf5),
    .B(_5505__bF$buf2),
    .C(\datapath.registers.1226[1] [10]),
    .Y(_9421_)
);

OAI21X1 _20776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5456__bF$buf1),
    .B(_9410__bF$buf4),
    .C(_9421_),
    .Y(_4758_)
);

OAI21X1 _20777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf4),
    .B(_5505__bF$buf1),
    .C(\datapath.registers.1226[1] [11]),
    .Y(_9422_)
);

OAI21X1 _20778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5458__bF$buf0),
    .B(_9410__bF$buf3),
    .C(_9422_),
    .Y(_4759_)
);

OAI21X1 _20779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf3),
    .B(_5505__bF$buf0),
    .C(\datapath.registers.1226[1] [12]),
    .Y(_9423_)
);

OAI21X1 _20780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460__bF$buf1),
    .B(_9410__bF$buf2),
    .C(_9423_),
    .Y(_4760_)
);

OAI21X1 _20781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf2),
    .B(_5505__bF$buf7),
    .C(\datapath.registers.1226[1] [13]),
    .Y(_9424_)
);

OAI21X1 _20782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5462__bF$buf1),
    .B(_9410__bF$buf1),
    .C(_9424_),
    .Y(_4761_)
);

OAI21X1 _20783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf1),
    .B(_5505__bF$buf6),
    .C(\datapath.registers.1226[1] [14]),
    .Y(_9425_)
);

OAI21X1 _20784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5464__bF$buf0),
    .B(_9410__bF$buf0),
    .C(_9425_),
    .Y(_4762_)
);

OAI21X1 _20785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf0),
    .B(_5505__bF$buf5),
    .C(\datapath.registers.1226[1] [15]),
    .Y(_9426_)
);

OAI21X1 _20786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466__bF$buf4),
    .B(_9410__bF$buf4),
    .C(_9426_),
    .Y(_4763_)
);

OAI21X1 _20787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf15),
    .B(_5505__bF$buf4),
    .C(\datapath.registers.1226[1] [16]),
    .Y(_9427_)
);

OAI21X1 _20788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468__bF$buf1),
    .B(_9410__bF$buf3),
    .C(_9427_),
    .Y(_4764_)
);

OAI21X1 _20789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf14),
    .B(_5505__bF$buf3),
    .C(\datapath.registers.1226[1] [17]),
    .Y(_9428_)
);

OAI21X1 _20790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470__bF$buf1),
    .B(_9410__bF$buf2),
    .C(_9428_),
    .Y(_4765_)
);

OAI21X1 _20791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf13),
    .B(_5505__bF$buf2),
    .C(\datapath.registers.1226[1] [18]),
    .Y(_9429_)
);

OAI21X1 _20792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5472__bF$buf0),
    .B(_9410__bF$buf1),
    .C(_9429_),
    .Y(_4766_)
);

OAI21X1 _20793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf12),
    .B(_5505__bF$buf1),
    .C(\datapath.registers.1226[1] [19]),
    .Y(_9430_)
);

OAI21X1 _20794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474__bF$buf0),
    .B(_9410__bF$buf0),
    .C(_9430_),
    .Y(_4767_)
);

OAI21X1 _20795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf11),
    .B(_5505__bF$buf0),
    .C(\datapath.registers.1226[1] [20]),
    .Y(_9431_)
);

OAI21X1 _20796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476__bF$buf0),
    .B(_9410__bF$buf4),
    .C(_9431_),
    .Y(_4769_)
);

OAI21X1 _20797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf10),
    .B(_5505__bF$buf7),
    .C(\datapath.registers.1226[1] [21]),
    .Y(_9432_)
);

OAI21X1 _20798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478__bF$buf1),
    .B(_9410__bF$buf3),
    .C(_9432_),
    .Y(_4770_)
);

OAI21X1 _20799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf9),
    .B(_5505__bF$buf6),
    .C(\datapath.registers.1226[1] [22]),
    .Y(_9433_)
);

OAI21X1 _20800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480__bF$buf0),
    .B(_9410__bF$buf2),
    .C(_9433_),
    .Y(_4771_)
);

OAI21X1 _20801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf8),
    .B(_5505__bF$buf5),
    .C(\datapath.registers.1226[1] [23]),
    .Y(_9434_)
);

OAI21X1 _20802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5482__bF$buf4),
    .B(_9410__bF$buf1),
    .C(_9434_),
    .Y(_4772_)
);

OAI21X1 _20803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf7),
    .B(_5505__bF$buf4),
    .C(\datapath.registers.1226[1] [24]),
    .Y(_9435_)
);

OAI21X1 _20804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5484__bF$buf0),
    .B(_9410__bF$buf0),
    .C(_9435_),
    .Y(_4773_)
);

OAI21X1 _20805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf6),
    .B(_5505__bF$buf3),
    .C(\datapath.registers.1226[1] [25]),
    .Y(_9436_)
);

OAI21X1 _20806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5486__bF$buf2),
    .B(_9410__bF$buf4),
    .C(_9436_),
    .Y(_4774_)
);

OAI21X1 _20807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf5),
    .B(_5505__bF$buf2),
    .C(\datapath.registers.1226[1] [26]),
    .Y(_9437_)
);

OAI21X1 _20808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488__bF$buf4),
    .B(_9410__bF$buf3),
    .C(_9437_),
    .Y(_4775_)
);

OAI21X1 _20809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf4),
    .B(_5505__bF$buf1),
    .C(\datapath.registers.1226[1] [27]),
    .Y(_9438_)
);

OAI21X1 _20810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5490__bF$buf1),
    .B(_9410__bF$buf2),
    .C(_9438_),
    .Y(_4776_)
);

OAI21X1 _20811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf3),
    .B(_5505__bF$buf0),
    .C(\datapath.registers.1226[1] [28]),
    .Y(_9439_)
);

OAI21X1 _20812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5492__bF$buf1),
    .B(_9410__bF$buf1),
    .C(_9439_),
    .Y(_4777_)
);

OAI21X1 _20813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf2),
    .B(_5505__bF$buf7),
    .C(\datapath.registers.1226[1] [29]),
    .Y(_9440_)
);

OAI21X1 _20814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494__bF$buf0),
    .B(_9410__bF$buf0),
    .C(_9440_),
    .Y(_4778_)
);

OAI21X1 _20815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf1),
    .B(_5505__bF$buf6),
    .C(\datapath.registers.1226[1] [30]),
    .Y(_9441_)
);

OAI21X1 _20816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496__bF$buf0),
    .B(_9410__bF$buf4),
    .C(_9441_),
    .Y(_4780_)
);

OAI21X1 _20817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5546__bF$buf0),
    .B(_5505__bF$buf5),
    .C(\datapath.registers.1226[1] [31]),
    .Y(_9442_)
);

OAI21X1 _20818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498__bF$buf0),
    .B(_9410__bF$buf3),
    .C(_9442_),
    .Y(_4781_)
);

BUFX2 _20819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [0]),
    .Y(_4405_)
);

BUFX2 _20820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [1]),
    .Y(_4416_)
);

BUFX2 _20821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [2]),
    .Y(_4427_)
);

BUFX2 _20822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [3]),
    .Y(_4430_)
);

BUFX2 _20823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [4]),
    .Y(_4431_)
);

BUFX2 _20824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [5]),
    .Y(_4432_)
);

BUFX2 _20825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [6]),
    .Y(_4433_)
);

BUFX2 _20826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [7]),
    .Y(_4434_)
);

BUFX2 _20827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [8]),
    .Y(_4435_)
);

BUFX2 _20828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [9]),
    .Y(_4436_)
);

BUFX2 _20829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [10]),
    .Y(_4406_)
);

BUFX2 _20830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [11]),
    .Y(_4407_)
);

BUFX2 _20831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [12]),
    .Y(_4408_)
);

BUFX2 _20832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [13]),
    .Y(_4409_)
);

BUFX2 _20833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [14]),
    .Y(_4410_)
);

BUFX2 _20834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [15]),
    .Y(_4411_)
);

BUFX2 _20835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [16]),
    .Y(_4412_)
);

BUFX2 _20836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [17]),
    .Y(_4413_)
);

BUFX2 _20837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [18]),
    .Y(_4414_)
);

BUFX2 _20838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [19]),
    .Y(_4415_)
);

BUFX2 _20839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [20]),
    .Y(_4417_)
);

BUFX2 _20840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [21]),
    .Y(_4418_)
);

BUFX2 _20841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [22]),
    .Y(_4419_)
);

BUFX2 _20842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [23]),
    .Y(_4420_)
);

BUFX2 _20843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [24]),
    .Y(_4421_)
);

BUFX2 _20844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [25]),
    .Y(_4422_)
);

BUFX2 _20845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [26]),
    .Y(_4423_)
);

BUFX2 _20846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [27]),
    .Y(_4424_)
);

BUFX2 _20847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [28]),
    .Y(_4425_)
);

BUFX2 _20848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [29]),
    .Y(_4426_)
);

BUFX2 _20849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [30]),
    .Y(_4428_)
);

BUFX2 _20850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.registers.1226[0] [31]),
    .Y(_4429_)
);

DFFPOSX1 _20851_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf24),
    .D(_4821_),
    .Q(\datapath.registers.1226[21] [0])
);

DFFPOSX1 _20852_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf23),
    .D(_4832_),
    .Q(\datapath.registers.1226[21] [1])
);

DFFPOSX1 _20853_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf22),
    .D(_4843_),
    .Q(\datapath.registers.1226[21] [2])
);

DFFPOSX1 _20854_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf21),
    .D(_4846_),
    .Q(\datapath.registers.1226[21] [3])
);

DFFPOSX1 _20855_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf20),
    .D(_4847_),
    .Q(\datapath.registers.1226[21] [4])
);

DFFPOSX1 _20856_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf19),
    .D(_4848_),
    .Q(\datapath.registers.1226[21] [5])
);

DFFPOSX1 _20857_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf18),
    .D(_4849_),
    .Q(\datapath.registers.1226[21] [6])
);

DFFPOSX1 _20858_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf17),
    .D(_4850_),
    .Q(\datapath.registers.1226[21] [7])
);

DFFPOSX1 _20859_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf16),
    .D(_4851_),
    .Q(\datapath.registers.1226[21] [8])
);

DFFPOSX1 _20860_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf15),
    .D(_4852_),
    .Q(\datapath.registers.1226[21] [9])
);

DFFPOSX1 _20861_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf14),
    .D(_4822_),
    .Q(\datapath.registers.1226[21] [10])
);

DFFPOSX1 _20862_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf13),
    .D(_4823_),
    .Q(\datapath.registers.1226[21] [11])
);

DFFPOSX1 _20863_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf12),
    .D(_4824_),
    .Q(\datapath.registers.1226[21] [12])
);

DFFPOSX1 _20864_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf11),
    .D(_4825_),
    .Q(\datapath.registers.1226[21] [13])
);

DFFPOSX1 _20865_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf10),
    .D(_4826_),
    .Q(\datapath.registers.1226[21] [14])
);

DFFPOSX1 _20866_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf9),
    .D(_4827_),
    .Q(\datapath.registers.1226[21] [15])
);

DFFPOSX1 _20867_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf8),
    .D(_4828_),
    .Q(\datapath.registers.1226[21] [16])
);

DFFPOSX1 _20868_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf7),
    .D(_4829_),
    .Q(\datapath.registers.1226[21] [17])
);

DFFPOSX1 _20869_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf6),
    .D(_4830_),
    .Q(\datapath.registers.1226[21] [18])
);

DFFPOSX1 _20870_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf5),
    .D(_4831_),
    .Q(\datapath.registers.1226[21] [19])
);

DFFPOSX1 _20871_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf4),
    .D(_4833_),
    .Q(\datapath.registers.1226[21] [20])
);

DFFPOSX1 _20872_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf3),
    .D(_4834_),
    .Q(\datapath.registers.1226[21] [21])
);

DFFPOSX1 _20873_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf2),
    .D(_4835_),
    .Q(\datapath.registers.1226[21] [22])
);

DFFPOSX1 _20874_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf1),
    .D(_4836_),
    .Q(\datapath.registers.1226[21] [23])
);

DFFPOSX1 _20875_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf0),
    .D(_4837_),
    .Q(\datapath.registers.1226[21] [24])
);

DFFPOSX1 _20876_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf153),
    .D(_4838_),
    .Q(\datapath.registers.1226[21] [25])
);

DFFPOSX1 _20877_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf152),
    .D(_4839_),
    .Q(\datapath.registers.1226[21] [26])
);

DFFPOSX1 _20878_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf151),
    .D(_4840_),
    .Q(\datapath.registers.1226[21] [27])
);

DFFPOSX1 _20879_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf150),
    .D(_4841_),
    .Q(\datapath.registers.1226[21] [28])
);

DFFPOSX1 _20880_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf149),
    .D(_4842_),
    .Q(\datapath.registers.1226[21] [29])
);

DFFPOSX1 _20881_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf148),
    .D(_4844_),
    .Q(\datapath.registers.1226[21] [30])
);

DFFPOSX1 _20882_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf147),
    .D(_4845_),
    .Q(\datapath.registers.1226[21] [31])
);

DFFPOSX1 _20883_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf146),
    .D(_4789_),
    .Q(\datapath.registers.1226[20] [0])
);

DFFPOSX1 _20884_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf145),
    .D(_4800_),
    .Q(\datapath.registers.1226[20] [1])
);

DFFPOSX1 _20885_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf144),
    .D(_4811_),
    .Q(\datapath.registers.1226[20] [2])
);

DFFPOSX1 _20886_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf143),
    .D(_4814_),
    .Q(\datapath.registers.1226[20] [3])
);

DFFPOSX1 _20887_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf142),
    .D(_4815_),
    .Q(\datapath.registers.1226[20] [4])
);

DFFPOSX1 _20888_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf141),
    .D(_4816_),
    .Q(\datapath.registers.1226[20] [5])
);

DFFPOSX1 _20889_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf140),
    .D(_4817_),
    .Q(\datapath.registers.1226[20] [6])
);

DFFPOSX1 _20890_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf139),
    .D(_4818_),
    .Q(\datapath.registers.1226[20] [7])
);

DFFPOSX1 _20891_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf138),
    .D(_4819_),
    .Q(\datapath.registers.1226[20] [8])
);

DFFPOSX1 _20892_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf137),
    .D(_4820_),
    .Q(\datapath.registers.1226[20] [9])
);

DFFPOSX1 _20893_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf136),
    .D(_4790_),
    .Q(\datapath.registers.1226[20] [10])
);

DFFPOSX1 _20894_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf135),
    .D(_4791_),
    .Q(\datapath.registers.1226[20] [11])
);

DFFPOSX1 _20895_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf134),
    .D(_4792_),
    .Q(\datapath.registers.1226[20] [12])
);

DFFPOSX1 _20896_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf133),
    .D(_4793_),
    .Q(\datapath.registers.1226[20] [13])
);

DFFPOSX1 _20897_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf132),
    .D(_4794_),
    .Q(\datapath.registers.1226[20] [14])
);

DFFPOSX1 _20898_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf131),
    .D(_4795_),
    .Q(\datapath.registers.1226[20] [15])
);

DFFPOSX1 _20899_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf130),
    .D(_4796_),
    .Q(\datapath.registers.1226[20] [16])
);

DFFPOSX1 _20900_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf129),
    .D(_4797_),
    .Q(\datapath.registers.1226[20] [17])
);

DFFPOSX1 _20901_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf128),
    .D(_4798_),
    .Q(\datapath.registers.1226[20] [18])
);

DFFPOSX1 _20902_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf127),
    .D(_4799_),
    .Q(\datapath.registers.1226[20] [19])
);

DFFPOSX1 _20903_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf126),
    .D(_4801_),
    .Q(\datapath.registers.1226[20] [20])
);

DFFPOSX1 _20904_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf125),
    .D(_4802_),
    .Q(\datapath.registers.1226[20] [21])
);

DFFPOSX1 _20905_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf124),
    .D(_4803_),
    .Q(\datapath.registers.1226[20] [22])
);

DFFPOSX1 _20906_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf123),
    .D(_4804_),
    .Q(\datapath.registers.1226[20] [23])
);

DFFPOSX1 _20907_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf122),
    .D(_4805_),
    .Q(\datapath.registers.1226[20] [24])
);

DFFPOSX1 _20908_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf121),
    .D(_4806_),
    .Q(\datapath.registers.1226[20] [25])
);

DFFPOSX1 _20909_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf120),
    .D(_4807_),
    .Q(\datapath.registers.1226[20] [26])
);

DFFPOSX1 _20910_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf119),
    .D(_4808_),
    .Q(\datapath.registers.1226[20] [27])
);

DFFPOSX1 _20911_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf118),
    .D(_4809_),
    .Q(\datapath.registers.1226[20] [28])
);

DFFPOSX1 _20912_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf117),
    .D(_4810_),
    .Q(\datapath.registers.1226[20] [29])
);

DFFPOSX1 _20913_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf116),
    .D(_4812_),
    .Q(\datapath.registers.1226[20] [30])
);

DFFPOSX1 _20914_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf115),
    .D(_4813_),
    .Q(\datapath.registers.1226[20] [31])
);

DFFPOSX1 _20915_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf114),
    .D(_4885_),
    .Q(\datapath.registers.1226[23] [0])
);

DFFPOSX1 _20916_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf113),
    .D(_4896_),
    .Q(\datapath.registers.1226[23] [1])
);

DFFPOSX1 _20917_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf112),
    .D(_4907_),
    .Q(\datapath.registers.1226[23] [2])
);

DFFPOSX1 _20918_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf111),
    .D(_4910_),
    .Q(\datapath.registers.1226[23] [3])
);

DFFPOSX1 _20919_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf110),
    .D(_4911_),
    .Q(\datapath.registers.1226[23] [4])
);

DFFPOSX1 _20920_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf109),
    .D(_4912_),
    .Q(\datapath.registers.1226[23] [5])
);

DFFPOSX1 _20921_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf108),
    .D(_4913_),
    .Q(\datapath.registers.1226[23] [6])
);

DFFPOSX1 _20922_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf107),
    .D(_4914_),
    .Q(\datapath.registers.1226[23] [7])
);

DFFPOSX1 _20923_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf106),
    .D(_4915_),
    .Q(\datapath.registers.1226[23] [8])
);

DFFPOSX1 _20924_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf105),
    .D(_4916_),
    .Q(\datapath.registers.1226[23] [9])
);

DFFPOSX1 _20925_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf104),
    .D(_4886_),
    .Q(\datapath.registers.1226[23] [10])
);

DFFPOSX1 _20926_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf103),
    .D(_4887_),
    .Q(\datapath.registers.1226[23] [11])
);

DFFPOSX1 _20927_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf102),
    .D(_4888_),
    .Q(\datapath.registers.1226[23] [12])
);

DFFPOSX1 _20928_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf101),
    .D(_4889_),
    .Q(\datapath.registers.1226[23] [13])
);

DFFPOSX1 _20929_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf100),
    .D(_4890_),
    .Q(\datapath.registers.1226[23] [14])
);

DFFPOSX1 _20930_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf99),
    .D(_4891_),
    .Q(\datapath.registers.1226[23] [15])
);

DFFPOSX1 _20931_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf98),
    .D(_4892_),
    .Q(\datapath.registers.1226[23] [16])
);

DFFPOSX1 _20932_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf97),
    .D(_4893_),
    .Q(\datapath.registers.1226[23] [17])
);

DFFPOSX1 _20933_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf96),
    .D(_4894_),
    .Q(\datapath.registers.1226[23] [18])
);

DFFPOSX1 _20934_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf95),
    .D(_4895_),
    .Q(\datapath.registers.1226[23] [19])
);

DFFPOSX1 _20935_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf94),
    .D(_4897_),
    .Q(\datapath.registers.1226[23] [20])
);

DFFPOSX1 _20936_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf93),
    .D(_4898_),
    .Q(\datapath.registers.1226[23] [21])
);

DFFPOSX1 _20937_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf92),
    .D(_4899_),
    .Q(\datapath.registers.1226[23] [22])
);

DFFPOSX1 _20938_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf91),
    .D(_4900_),
    .Q(\datapath.registers.1226[23] [23])
);

DFFPOSX1 _20939_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf90),
    .D(_4901_),
    .Q(\datapath.registers.1226[23] [24])
);

DFFPOSX1 _20940_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf89),
    .D(_4902_),
    .Q(\datapath.registers.1226[23] [25])
);

DFFPOSX1 _20941_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf88),
    .D(_4903_),
    .Q(\datapath.registers.1226[23] [26])
);

DFFPOSX1 _20942_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf87),
    .D(_4904_),
    .Q(\datapath.registers.1226[23] [27])
);

DFFPOSX1 _20943_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf86),
    .D(_4905_),
    .Q(\datapath.registers.1226[23] [28])
);

DFFPOSX1 _20944_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf85),
    .D(_4906_),
    .Q(\datapath.registers.1226[23] [29])
);

DFFPOSX1 _20945_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf84),
    .D(_4908_),
    .Q(\datapath.registers.1226[23] [30])
);

DFFPOSX1 _20946_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf83),
    .D(_4909_),
    .Q(\datapath.registers.1226[23] [31])
);

DFFPOSX1 _20947_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf82),
    .D(_4853_),
    .Q(\datapath.registers.1226[22] [0])
);

DFFPOSX1 _20948_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf81),
    .D(_4864_),
    .Q(\datapath.registers.1226[22] [1])
);

DFFPOSX1 _20949_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf80),
    .D(_4875_),
    .Q(\datapath.registers.1226[22] [2])
);

DFFPOSX1 _20950_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf79),
    .D(_4878_),
    .Q(\datapath.registers.1226[22] [3])
);

DFFPOSX1 _20951_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf78),
    .D(_4879_),
    .Q(\datapath.registers.1226[22] [4])
);

DFFPOSX1 _20952_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf77),
    .D(_4880_),
    .Q(\datapath.registers.1226[22] [5])
);

DFFPOSX1 _20953_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf76),
    .D(_4881_),
    .Q(\datapath.registers.1226[22] [6])
);

DFFPOSX1 _20954_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf75),
    .D(_4882_),
    .Q(\datapath.registers.1226[22] [7])
);

DFFPOSX1 _20955_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf74),
    .D(_4883_),
    .Q(\datapath.registers.1226[22] [8])
);

DFFPOSX1 _20956_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf73),
    .D(_4884_),
    .Q(\datapath.registers.1226[22] [9])
);

DFFPOSX1 _20957_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf72),
    .D(_4854_),
    .Q(\datapath.registers.1226[22] [10])
);

DFFPOSX1 _20958_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf71),
    .D(_4855_),
    .Q(\datapath.registers.1226[22] [11])
);

DFFPOSX1 _20959_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf70),
    .D(_4856_),
    .Q(\datapath.registers.1226[22] [12])
);

DFFPOSX1 _20960_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf69),
    .D(_4857_),
    .Q(\datapath.registers.1226[22] [13])
);

DFFPOSX1 _20961_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf68),
    .D(_4858_),
    .Q(\datapath.registers.1226[22] [14])
);

DFFPOSX1 _20962_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf67),
    .D(_4859_),
    .Q(\datapath.registers.1226[22] [15])
);

DFFPOSX1 _20963_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf66),
    .D(_4860_),
    .Q(\datapath.registers.1226[22] [16])
);

DFFPOSX1 _20964_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf65),
    .D(_4861_),
    .Q(\datapath.registers.1226[22] [17])
);

DFFPOSX1 _20965_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf64),
    .D(_4862_),
    .Q(\datapath.registers.1226[22] [18])
);

DFFPOSX1 _20966_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf63),
    .D(_4863_),
    .Q(\datapath.registers.1226[22] [19])
);

DFFPOSX1 _20967_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf62),
    .D(_4865_),
    .Q(\datapath.registers.1226[22] [20])
);

DFFPOSX1 _20968_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf61),
    .D(_4866_),
    .Q(\datapath.registers.1226[22] [21])
);

DFFPOSX1 _20969_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf60),
    .D(_4867_),
    .Q(\datapath.registers.1226[22] [22])
);

DFFPOSX1 _20970_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf59),
    .D(_4868_),
    .Q(\datapath.registers.1226[22] [23])
);

DFFPOSX1 _20971_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf58),
    .D(_4869_),
    .Q(\datapath.registers.1226[22] [24])
);

DFFPOSX1 _20972_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf57),
    .D(_4870_),
    .Q(\datapath.registers.1226[22] [25])
);

DFFPOSX1 _20973_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf56),
    .D(_4871_),
    .Q(\datapath.registers.1226[22] [26])
);

DFFPOSX1 _20974_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf55),
    .D(_4872_),
    .Q(\datapath.registers.1226[22] [27])
);

DFFPOSX1 _20975_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf54),
    .D(_4873_),
    .Q(\datapath.registers.1226[22] [28])
);

DFFPOSX1 _20976_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf53),
    .D(_4874_),
    .Q(\datapath.registers.1226[22] [29])
);

DFFPOSX1 _20977_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf52),
    .D(_4876_),
    .Q(\datapath.registers.1226[22] [30])
);

DFFPOSX1 _20978_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf51),
    .D(_4877_),
    .Q(\datapath.registers.1226[22] [31])
);

DFFPOSX1 _20979_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf50),
    .D(_5397_),
    .Q(\datapath.registers.1226[9] [0])
);

DFFPOSX1 _20980_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf49),
    .D(_5408_),
    .Q(\datapath.registers.1226[9] [1])
);

DFFPOSX1 _20981_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf48),
    .D(_5419_),
    .Q(\datapath.registers.1226[9] [2])
);

DFFPOSX1 _20982_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf47),
    .D(_5422_),
    .Q(\datapath.registers.1226[9] [3])
);

DFFPOSX1 _20983_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf46),
    .D(_5423_),
    .Q(\datapath.registers.1226[9] [4])
);

DFFPOSX1 _20984_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf45),
    .D(_5424_),
    .Q(\datapath.registers.1226[9] [5])
);

DFFPOSX1 _20985_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf44),
    .D(_5425_),
    .Q(\datapath.registers.1226[9] [6])
);

DFFPOSX1 _20986_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf43),
    .D(_5426_),
    .Q(\datapath.registers.1226[9] [7])
);

DFFPOSX1 _20987_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf42),
    .D(_5427_),
    .Q(\datapath.registers.1226[9] [8])
);

DFFPOSX1 _20988_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf41),
    .D(_5428_),
    .Q(\datapath.registers.1226[9] [9])
);

DFFPOSX1 _20989_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf40),
    .D(_5398_),
    .Q(\datapath.registers.1226[9] [10])
);

DFFPOSX1 _20990_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf39),
    .D(_5399_),
    .Q(\datapath.registers.1226[9] [11])
);

DFFPOSX1 _20991_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf38),
    .D(_5400_),
    .Q(\datapath.registers.1226[9] [12])
);

DFFPOSX1 _20992_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf37),
    .D(_5401_),
    .Q(\datapath.registers.1226[9] [13])
);

DFFPOSX1 _20993_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf36),
    .D(_5402_),
    .Q(\datapath.registers.1226[9] [14])
);

DFFPOSX1 _20994_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf35),
    .D(_5403_),
    .Q(\datapath.registers.1226[9] [15])
);

DFFPOSX1 _20995_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf34),
    .D(_5404_),
    .Q(\datapath.registers.1226[9] [16])
);

DFFPOSX1 _20996_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf33),
    .D(_5405_),
    .Q(\datapath.registers.1226[9] [17])
);

DFFPOSX1 _20997_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf32),
    .D(_5406_),
    .Q(\datapath.registers.1226[9] [18])
);

DFFPOSX1 _20998_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf31),
    .D(_5407_),
    .Q(\datapath.registers.1226[9] [19])
);

DFFPOSX1 _20999_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf30),
    .D(_5409_),
    .Q(\datapath.registers.1226[9] [20])
);

DFFPOSX1 _21000_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf29),
    .D(_5410_),
    .Q(\datapath.registers.1226[9] [21])
);

DFFPOSX1 _21001_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf28),
    .D(_5411_),
    .Q(\datapath.registers.1226[9] [22])
);

DFFPOSX1 _21002_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf27),
    .D(_5412_),
    .Q(\datapath.registers.1226[9] [23])
);

DFFPOSX1 _21003_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf26),
    .D(_5413_),
    .Q(\datapath.registers.1226[9] [24])
);

DFFPOSX1 _21004_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf25),
    .D(_5414_),
    .Q(\datapath.registers.1226[9] [25])
);

DFFPOSX1 _21005_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf24),
    .D(_5415_),
    .Q(\datapath.registers.1226[9] [26])
);

DFFPOSX1 _21006_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf23),
    .D(_5416_),
    .Q(\datapath.registers.1226[9] [27])
);

DFFPOSX1 _21007_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf22),
    .D(_5417_),
    .Q(\datapath.registers.1226[9] [28])
);

DFFPOSX1 _21008_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf21),
    .D(_5418_),
    .Q(\datapath.registers.1226[9] [29])
);

DFFPOSX1 _21009_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf20),
    .D(_5420_),
    .Q(\datapath.registers.1226[9] [30])
);

DFFPOSX1 _21010_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf19),
    .D(_5421_),
    .Q(\datapath.registers.1226[9] [31])
);

DFFPOSX1 _21011_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf18),
    .D(_4437_),
    .Q(\datapath.registers.1226[10] [0])
);

DFFPOSX1 _21012_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf17),
    .D(_4448_),
    .Q(\datapath.registers.1226[10] [1])
);

DFFPOSX1 _21013_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf16),
    .D(_4459_),
    .Q(\datapath.registers.1226[10] [2])
);

DFFPOSX1 _21014_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf15),
    .D(_4462_),
    .Q(\datapath.registers.1226[10] [3])
);

DFFPOSX1 _21015_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf14),
    .D(_4463_),
    .Q(\datapath.registers.1226[10] [4])
);

DFFPOSX1 _21016_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf13),
    .D(_4464_),
    .Q(\datapath.registers.1226[10] [5])
);

DFFPOSX1 _21017_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf12),
    .D(_4465_),
    .Q(\datapath.registers.1226[10] [6])
);

DFFPOSX1 _21018_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf11),
    .D(_4466_),
    .Q(\datapath.registers.1226[10] [7])
);

DFFPOSX1 _21019_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf10),
    .D(_4467_),
    .Q(\datapath.registers.1226[10] [8])
);

DFFPOSX1 _21020_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf9),
    .D(_4468_),
    .Q(\datapath.registers.1226[10] [9])
);

DFFPOSX1 _21021_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf8),
    .D(_4438_),
    .Q(\datapath.registers.1226[10] [10])
);

DFFPOSX1 _21022_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf7),
    .D(_4439_),
    .Q(\datapath.registers.1226[10] [11])
);

DFFPOSX1 _21023_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf6),
    .D(_4440_),
    .Q(\datapath.registers.1226[10] [12])
);

DFFPOSX1 _21024_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf5),
    .D(_4441_),
    .Q(\datapath.registers.1226[10] [13])
);

DFFPOSX1 _21025_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf4),
    .D(_4442_),
    .Q(\datapath.registers.1226[10] [14])
);

DFFPOSX1 _21026_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf3),
    .D(_4443_),
    .Q(\datapath.registers.1226[10] [15])
);

DFFPOSX1 _21027_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf2),
    .D(_4444_),
    .Q(\datapath.registers.1226[10] [16])
);

DFFPOSX1 _21028_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf1),
    .D(_4445_),
    .Q(\datapath.registers.1226[10] [17])
);

DFFPOSX1 _21029_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf0),
    .D(_4446_),
    .Q(\datapath.registers.1226[10] [18])
);

DFFPOSX1 _21030_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf153),
    .D(_4447_),
    .Q(\datapath.registers.1226[10] [19])
);

DFFPOSX1 _21031_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf152),
    .D(_4449_),
    .Q(\datapath.registers.1226[10] [20])
);

DFFPOSX1 _21032_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf151),
    .D(_4450_),
    .Q(\datapath.registers.1226[10] [21])
);

DFFPOSX1 _21033_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf150),
    .D(_4451_),
    .Q(\datapath.registers.1226[10] [22])
);

DFFPOSX1 _21034_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf149),
    .D(_4452_),
    .Q(\datapath.registers.1226[10] [23])
);

DFFPOSX1 _21035_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf148),
    .D(_4453_),
    .Q(\datapath.registers.1226[10] [24])
);

DFFPOSX1 _21036_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf147),
    .D(_4454_),
    .Q(\datapath.registers.1226[10] [25])
);

DFFPOSX1 _21037_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf146),
    .D(_4455_),
    .Q(\datapath.registers.1226[10] [26])
);

DFFPOSX1 _21038_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf145),
    .D(_4456_),
    .Q(\datapath.registers.1226[10] [27])
);

DFFPOSX1 _21039_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf144),
    .D(_4457_),
    .Q(\datapath.registers.1226[10] [28])
);

DFFPOSX1 _21040_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf143),
    .D(_4458_),
    .Q(\datapath.registers.1226[10] [29])
);

DFFPOSX1 _21041_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf142),
    .D(_4460_),
    .Q(\datapath.registers.1226[10] [30])
);

DFFPOSX1 _21042_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf141),
    .D(_4461_),
    .Q(\datapath.registers.1226[10] [31])
);

DFFPOSX1 _21043_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf140),
    .D(_5013_),
    .Q(\datapath.registers.1226[27] [0])
);

DFFPOSX1 _21044_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf139),
    .D(_5024_),
    .Q(\datapath.registers.1226[27] [1])
);

DFFPOSX1 _21045_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf138),
    .D(_5035_),
    .Q(\datapath.registers.1226[27] [2])
);

DFFPOSX1 _21046_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf137),
    .D(_5038_),
    .Q(\datapath.registers.1226[27] [3])
);

DFFPOSX1 _21047_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf136),
    .D(_5039_),
    .Q(\datapath.registers.1226[27] [4])
);

DFFPOSX1 _21048_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf135),
    .D(_5040_),
    .Q(\datapath.registers.1226[27] [5])
);

DFFPOSX1 _21049_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf134),
    .D(_5041_),
    .Q(\datapath.registers.1226[27] [6])
);

DFFPOSX1 _21050_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf133),
    .D(_5042_),
    .Q(\datapath.registers.1226[27] [7])
);

DFFPOSX1 _21051_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf132),
    .D(_5043_),
    .Q(\datapath.registers.1226[27] [8])
);

DFFPOSX1 _21052_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf131),
    .D(_5044_),
    .Q(\datapath.registers.1226[27] [9])
);

DFFPOSX1 _21053_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf130),
    .D(_5014_),
    .Q(\datapath.registers.1226[27] [10])
);

DFFPOSX1 _21054_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf129),
    .D(_5015_),
    .Q(\datapath.registers.1226[27] [11])
);

DFFPOSX1 _21055_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf128),
    .D(_5016_),
    .Q(\datapath.registers.1226[27] [12])
);

DFFPOSX1 _21056_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf127),
    .D(_5017_),
    .Q(\datapath.registers.1226[27] [13])
);

DFFPOSX1 _21057_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf126),
    .D(_5018_),
    .Q(\datapath.registers.1226[27] [14])
);

DFFPOSX1 _21058_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf125),
    .D(_5019_),
    .Q(\datapath.registers.1226[27] [15])
);

DFFPOSX1 _21059_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf124),
    .D(_5020_),
    .Q(\datapath.registers.1226[27] [16])
);

DFFPOSX1 _21060_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf123),
    .D(_5021_),
    .Q(\datapath.registers.1226[27] [17])
);

DFFPOSX1 _21061_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf122),
    .D(_5022_),
    .Q(\datapath.registers.1226[27] [18])
);

DFFPOSX1 _21062_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf121),
    .D(_5023_),
    .Q(\datapath.registers.1226[27] [19])
);

DFFPOSX1 _21063_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf120),
    .D(_5025_),
    .Q(\datapath.registers.1226[27] [20])
);

DFFPOSX1 _21064_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf119),
    .D(_5026_),
    .Q(\datapath.registers.1226[27] [21])
);

DFFPOSX1 _21065_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf118),
    .D(_5027_),
    .Q(\datapath.registers.1226[27] [22])
);

DFFPOSX1 _21066_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf117),
    .D(_5028_),
    .Q(\datapath.registers.1226[27] [23])
);

DFFPOSX1 _21067_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf116),
    .D(_5029_),
    .Q(\datapath.registers.1226[27] [24])
);

DFFPOSX1 _21068_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf115),
    .D(_5030_),
    .Q(\datapath.registers.1226[27] [25])
);

DFFPOSX1 _21069_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf114),
    .D(_5031_),
    .Q(\datapath.registers.1226[27] [26])
);

DFFPOSX1 _21070_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf113),
    .D(_5032_),
    .Q(\datapath.registers.1226[27] [27])
);

DFFPOSX1 _21071_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf112),
    .D(_5033_),
    .Q(\datapath.registers.1226[27] [28])
);

DFFPOSX1 _21072_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf111),
    .D(_5034_),
    .Q(\datapath.registers.1226[27] [29])
);

DFFPOSX1 _21073_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf110),
    .D(_5036_),
    .Q(\datapath.registers.1226[27] [30])
);

DFFPOSX1 _21074_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf109),
    .D(_5037_),
    .Q(\datapath.registers.1226[27] [31])
);

DFFPOSX1 _21075_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf108),
    .D(_4597_),
    .Q(\datapath.registers.1226[15] [0])
);

DFFPOSX1 _21076_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf107),
    .D(_4608_),
    .Q(\datapath.registers.1226[15] [1])
);

DFFPOSX1 _21077_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf106),
    .D(_4619_),
    .Q(\datapath.registers.1226[15] [2])
);

DFFPOSX1 _21078_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf105),
    .D(_4622_),
    .Q(\datapath.registers.1226[15] [3])
);

DFFPOSX1 _21079_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf104),
    .D(_4623_),
    .Q(\datapath.registers.1226[15] [4])
);

DFFPOSX1 _21080_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf103),
    .D(_4624_),
    .Q(\datapath.registers.1226[15] [5])
);

DFFPOSX1 _21081_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf102),
    .D(_4625_),
    .Q(\datapath.registers.1226[15] [6])
);

DFFPOSX1 _21082_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf101),
    .D(_4626_),
    .Q(\datapath.registers.1226[15] [7])
);

DFFPOSX1 _21083_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf100),
    .D(_4627_),
    .Q(\datapath.registers.1226[15] [8])
);

DFFPOSX1 _21084_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf99),
    .D(_4628_),
    .Q(\datapath.registers.1226[15] [9])
);

DFFPOSX1 _21085_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf98),
    .D(_4598_),
    .Q(\datapath.registers.1226[15] [10])
);

DFFPOSX1 _21086_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf97),
    .D(_4599_),
    .Q(\datapath.registers.1226[15] [11])
);

DFFPOSX1 _21087_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf96),
    .D(_4600_),
    .Q(\datapath.registers.1226[15] [12])
);

DFFPOSX1 _21088_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf95),
    .D(_4601_),
    .Q(\datapath.registers.1226[15] [13])
);

DFFPOSX1 _21089_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf94),
    .D(_4602_),
    .Q(\datapath.registers.1226[15] [14])
);

DFFPOSX1 _21090_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf93),
    .D(_4603_),
    .Q(\datapath.registers.1226[15] [15])
);

DFFPOSX1 _21091_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf92),
    .D(_4604_),
    .Q(\datapath.registers.1226[15] [16])
);

DFFPOSX1 _21092_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf91),
    .D(_4605_),
    .Q(\datapath.registers.1226[15] [17])
);

DFFPOSX1 _21093_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf90),
    .D(_4606_),
    .Q(\datapath.registers.1226[15] [18])
);

DFFPOSX1 _21094_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf89),
    .D(_4607_),
    .Q(\datapath.registers.1226[15] [19])
);

DFFPOSX1 _21095_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf88),
    .D(_4609_),
    .Q(\datapath.registers.1226[15] [20])
);

DFFPOSX1 _21096_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf87),
    .D(_4610_),
    .Q(\datapath.registers.1226[15] [21])
);

DFFPOSX1 _21097_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf86),
    .D(_4611_),
    .Q(\datapath.registers.1226[15] [22])
);

DFFPOSX1 _21098_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf85),
    .D(_4612_),
    .Q(\datapath.registers.1226[15] [23])
);

DFFPOSX1 _21099_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf84),
    .D(_4613_),
    .Q(\datapath.registers.1226[15] [24])
);

DFFPOSX1 _21100_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf83),
    .D(_4614_),
    .Q(\datapath.registers.1226[15] [25])
);

DFFPOSX1 _21101_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf82),
    .D(_4615_),
    .Q(\datapath.registers.1226[15] [26])
);

DFFPOSX1 _21102_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf81),
    .D(_4616_),
    .Q(\datapath.registers.1226[15] [27])
);

DFFPOSX1 _21103_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf80),
    .D(_4617_),
    .Q(\datapath.registers.1226[15] [28])
);

DFFPOSX1 _21104_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf79),
    .D(_4618_),
    .Q(\datapath.registers.1226[15] [29])
);

DFFPOSX1 _21105_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf78),
    .D(_4620_),
    .Q(\datapath.registers.1226[15] [30])
);

DFFPOSX1 _21106_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf77),
    .D(_4621_),
    .Q(\datapath.registers.1226[15] [31])
);

DFFPOSX1 _21107_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf76),
    .D(_5173_),
    .Q(\datapath.registers.1226[31] [0])
);

DFFPOSX1 _21108_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf75),
    .D(_5184_),
    .Q(\datapath.registers.1226[31] [1])
);

DFFPOSX1 _21109_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf74),
    .D(_5195_),
    .Q(\datapath.registers.1226[31] [2])
);

DFFPOSX1 _21110_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf73),
    .D(_5198_),
    .Q(\datapath.registers.1226[31] [3])
);

DFFPOSX1 _21111_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf72),
    .D(_5199_),
    .Q(\datapath.registers.1226[31] [4])
);

DFFPOSX1 _21112_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf71),
    .D(_5200_),
    .Q(\datapath.registers.1226[31] [5])
);

DFFPOSX1 _21113_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf70),
    .D(_5201_),
    .Q(\datapath.registers.1226[31] [6])
);

DFFPOSX1 _21114_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf69),
    .D(_5202_),
    .Q(\datapath.registers.1226[31] [7])
);

DFFPOSX1 _21115_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf68),
    .D(_5203_),
    .Q(\datapath.registers.1226[31] [8])
);

DFFPOSX1 _21116_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf67),
    .D(_5204_),
    .Q(\datapath.registers.1226[31] [9])
);

DFFPOSX1 _21117_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf66),
    .D(_5174_),
    .Q(\datapath.registers.1226[31] [10])
);

DFFPOSX1 _21118_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf65),
    .D(_5175_),
    .Q(\datapath.registers.1226[31] [11])
);

DFFPOSX1 _21119_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf64),
    .D(_5176_),
    .Q(\datapath.registers.1226[31] [12])
);

DFFPOSX1 _21120_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf63),
    .D(_5177_),
    .Q(\datapath.registers.1226[31] [13])
);

DFFPOSX1 _21121_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf62),
    .D(_5178_),
    .Q(\datapath.registers.1226[31] [14])
);

DFFPOSX1 _21122_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf61),
    .D(_5179_),
    .Q(\datapath.registers.1226[31] [15])
);

DFFPOSX1 _21123_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf60),
    .D(_5180_),
    .Q(\datapath.registers.1226[31] [16])
);

DFFPOSX1 _21124_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf59),
    .D(_5181_),
    .Q(\datapath.registers.1226[31] [17])
);

DFFPOSX1 _21125_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf58),
    .D(_5182_),
    .Q(\datapath.registers.1226[31] [18])
);

DFFPOSX1 _21126_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf57),
    .D(_5183_),
    .Q(\datapath.registers.1226[31] [19])
);

DFFPOSX1 _21127_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf56),
    .D(_5185_),
    .Q(\datapath.registers.1226[31] [20])
);

DFFPOSX1 _21128_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf55),
    .D(_5186_),
    .Q(\datapath.registers.1226[31] [21])
);

DFFPOSX1 _21129_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf54),
    .D(_5187_),
    .Q(\datapath.registers.1226[31] [22])
);

DFFPOSX1 _21130_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf53),
    .D(_5188_),
    .Q(\datapath.registers.1226[31] [23])
);

DFFPOSX1 _21131_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf52),
    .D(_5189_),
    .Q(\datapath.registers.1226[31] [24])
);

DFFPOSX1 _21132_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf51),
    .D(_5190_),
    .Q(\datapath.registers.1226[31] [25])
);

DFFPOSX1 _21133_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf50),
    .D(_5191_),
    .Q(\datapath.registers.1226[31] [26])
);

DFFPOSX1 _21134_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf49),
    .D(_5192_),
    .Q(\datapath.registers.1226[31] [27])
);

DFFPOSX1 _21135_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf48),
    .D(_5193_),
    .Q(\datapath.registers.1226[31] [28])
);

DFFPOSX1 _21136_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf47),
    .D(_5194_),
    .Q(\datapath.registers.1226[31] [29])
);

DFFPOSX1 _21137_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf46),
    .D(_5196_),
    .Q(\datapath.registers.1226[31] [30])
);

DFFPOSX1 _21138_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf45),
    .D(_5197_),
    .Q(\datapath.registers.1226[31] [31])
);

DFFPOSX1 _21139_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf44),
    .D(_5109_),
    .Q(\datapath.registers.1226[2] [0])
);

DFFPOSX1 _21140_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf43),
    .D(_5120_),
    .Q(\datapath.registers.1226[2] [1])
);

DFFPOSX1 _21141_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf42),
    .D(_5131_),
    .Q(\datapath.registers.1226[2] [2])
);

DFFPOSX1 _21142_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf41),
    .D(_5134_),
    .Q(\datapath.registers.1226[2] [3])
);

DFFPOSX1 _21143_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf40),
    .D(_5135_),
    .Q(\datapath.registers.1226[2] [4])
);

DFFPOSX1 _21144_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf39),
    .D(_5136_),
    .Q(\datapath.registers.1226[2] [5])
);

DFFPOSX1 _21145_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf38),
    .D(_5137_),
    .Q(\datapath.registers.1226[2] [6])
);

DFFPOSX1 _21146_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf37),
    .D(_5138_),
    .Q(\datapath.registers.1226[2] [7])
);

DFFPOSX1 _21147_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf36),
    .D(_5139_),
    .Q(\datapath.registers.1226[2] [8])
);

DFFPOSX1 _21148_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf35),
    .D(_5140_),
    .Q(\datapath.registers.1226[2] [9])
);

DFFPOSX1 _21149_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf34),
    .D(_5110_),
    .Q(\datapath.registers.1226[2] [10])
);

DFFPOSX1 _21150_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf33),
    .D(_5111_),
    .Q(\datapath.registers.1226[2] [11])
);

DFFPOSX1 _21151_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf32),
    .D(_5112_),
    .Q(\datapath.registers.1226[2] [12])
);

DFFPOSX1 _21152_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf31),
    .D(_5113_),
    .Q(\datapath.registers.1226[2] [13])
);

DFFPOSX1 _21153_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf30),
    .D(_5114_),
    .Q(\datapath.registers.1226[2] [14])
);

DFFPOSX1 _21154_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf29),
    .D(_5115_),
    .Q(\datapath.registers.1226[2] [15])
);

DFFPOSX1 _21155_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf28),
    .D(_5116_),
    .Q(\datapath.registers.1226[2] [16])
);

DFFPOSX1 _21156_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf27),
    .D(_5117_),
    .Q(\datapath.registers.1226[2] [17])
);

DFFPOSX1 _21157_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf26),
    .D(_5118_),
    .Q(\datapath.registers.1226[2] [18])
);

DFFPOSX1 _21158_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf25),
    .D(_5119_),
    .Q(\datapath.registers.1226[2] [19])
);

DFFPOSX1 _21159_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf24),
    .D(_5121_),
    .Q(\datapath.registers.1226[2] [20])
);

DFFPOSX1 _21160_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf23),
    .D(_5122_),
    .Q(\datapath.registers.1226[2] [21])
);

DFFPOSX1 _21161_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf22),
    .D(_5123_),
    .Q(\datapath.registers.1226[2] [22])
);

DFFPOSX1 _21162_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf21),
    .D(_5124_),
    .Q(\datapath.registers.1226[2] [23])
);

DFFPOSX1 _21163_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf20),
    .D(_5125_),
    .Q(\datapath.registers.1226[2] [24])
);

DFFPOSX1 _21164_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf19),
    .D(_5126_),
    .Q(\datapath.registers.1226[2] [25])
);

DFFPOSX1 _21165_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf18),
    .D(_5127_),
    .Q(\datapath.registers.1226[2] [26])
);

DFFPOSX1 _21166_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf17),
    .D(_5128_),
    .Q(\datapath.registers.1226[2] [27])
);

DFFPOSX1 _21167_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf16),
    .D(_5129_),
    .Q(\datapath.registers.1226[2] [28])
);

DFFPOSX1 _21168_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf15),
    .D(_5130_),
    .Q(\datapath.registers.1226[2] [29])
);

DFFPOSX1 _21169_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf14),
    .D(_5132_),
    .Q(\datapath.registers.1226[2] [30])
);

DFFPOSX1 _21170_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf13),
    .D(_5133_),
    .Q(\datapath.registers.1226[2] [31])
);

DFFPOSX1 _21171_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf12),
    .D(_5205_),
    .Q(\datapath.registers.1226[3] [0])
);

DFFPOSX1 _21172_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf11),
    .D(_5216_),
    .Q(\datapath.registers.1226[3] [1])
);

DFFPOSX1 _21173_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf10),
    .D(_5227_),
    .Q(\datapath.registers.1226[3] [2])
);

DFFPOSX1 _21174_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf9),
    .D(_5230_),
    .Q(\datapath.registers.1226[3] [3])
);

DFFPOSX1 _21175_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf8),
    .D(_5231_),
    .Q(\datapath.registers.1226[3] [4])
);

DFFPOSX1 _21176_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf7),
    .D(_5232_),
    .Q(\datapath.registers.1226[3] [5])
);

DFFPOSX1 _21177_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf6),
    .D(_5233_),
    .Q(\datapath.registers.1226[3] [6])
);

DFFPOSX1 _21178_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf5),
    .D(_5234_),
    .Q(\datapath.registers.1226[3] [7])
);

DFFPOSX1 _21179_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf4),
    .D(_5235_),
    .Q(\datapath.registers.1226[3] [8])
);

DFFPOSX1 _21180_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf3),
    .D(_5236_),
    .Q(\datapath.registers.1226[3] [9])
);

DFFPOSX1 _21181_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf2),
    .D(_5206_),
    .Q(\datapath.registers.1226[3] [10])
);

DFFPOSX1 _21182_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf1),
    .D(_5207_),
    .Q(\datapath.registers.1226[3] [11])
);

DFFPOSX1 _21183_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf0),
    .D(_5208_),
    .Q(\datapath.registers.1226[3] [12])
);

DFFPOSX1 _21184_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf153),
    .D(_5209_),
    .Q(\datapath.registers.1226[3] [13])
);

DFFPOSX1 _21185_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf152),
    .D(_5210_),
    .Q(\datapath.registers.1226[3] [14])
);

DFFPOSX1 _21186_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf151),
    .D(_5211_),
    .Q(\datapath.registers.1226[3] [15])
);

DFFPOSX1 _21187_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf150),
    .D(_5212_),
    .Q(\datapath.registers.1226[3] [16])
);

DFFPOSX1 _21188_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf149),
    .D(_5213_),
    .Q(\datapath.registers.1226[3] [17])
);

DFFPOSX1 _21189_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf148),
    .D(_5214_),
    .Q(\datapath.registers.1226[3] [18])
);

DFFPOSX1 _21190_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf147),
    .D(_5215_),
    .Q(\datapath.registers.1226[3] [19])
);

DFFPOSX1 _21191_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf146),
    .D(_5217_),
    .Q(\datapath.registers.1226[3] [20])
);

DFFPOSX1 _21192_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf145),
    .D(_5218_),
    .Q(\datapath.registers.1226[3] [21])
);

DFFPOSX1 _21193_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf144),
    .D(_5219_),
    .Q(\datapath.registers.1226[3] [22])
);

DFFPOSX1 _21194_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf143),
    .D(_5220_),
    .Q(\datapath.registers.1226[3] [23])
);

DFFPOSX1 _21195_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf142),
    .D(_5221_),
    .Q(\datapath.registers.1226[3] [24])
);

DFFPOSX1 _21196_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf141),
    .D(_5222_),
    .Q(\datapath.registers.1226[3] [25])
);

DFFPOSX1 _21197_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf140),
    .D(_5223_),
    .Q(\datapath.registers.1226[3] [26])
);

DFFPOSX1 _21198_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf139),
    .D(_5224_),
    .Q(\datapath.registers.1226[3] [27])
);

DFFPOSX1 _21199_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf138),
    .D(_5225_),
    .Q(\datapath.registers.1226[3] [28])
);

DFFPOSX1 _21200_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf137),
    .D(_5226_),
    .Q(\datapath.registers.1226[3] [29])
);

DFFPOSX1 _21201_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf136),
    .D(_5228_),
    .Q(\datapath.registers.1226[3] [30])
);

DFFPOSX1 _21202_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf135),
    .D(_5229_),
    .Q(\datapath.registers.1226[3] [31])
);

DFFPOSX1 _21203_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf134),
    .D(_4629_),
    .Q(\datapath.registers.1226[16] [0])
);

DFFPOSX1 _21204_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf133),
    .D(_4640_),
    .Q(\datapath.registers.1226[16] [1])
);

DFFPOSX1 _21205_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf132),
    .D(_4651_),
    .Q(\datapath.registers.1226[16] [2])
);

DFFPOSX1 _21206_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf131),
    .D(_4654_),
    .Q(\datapath.registers.1226[16] [3])
);

DFFPOSX1 _21207_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf130),
    .D(_4655_),
    .Q(\datapath.registers.1226[16] [4])
);

DFFPOSX1 _21208_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf129),
    .D(_4656_),
    .Q(\datapath.registers.1226[16] [5])
);

DFFPOSX1 _21209_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf128),
    .D(_4657_),
    .Q(\datapath.registers.1226[16] [6])
);

DFFPOSX1 _21210_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf127),
    .D(_4658_),
    .Q(\datapath.registers.1226[16] [7])
);

DFFPOSX1 _21211_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf126),
    .D(_4659_),
    .Q(\datapath.registers.1226[16] [8])
);

DFFPOSX1 _21212_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf125),
    .D(_4660_),
    .Q(\datapath.registers.1226[16] [9])
);

DFFPOSX1 _21213_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf124),
    .D(_4630_),
    .Q(\datapath.registers.1226[16] [10])
);

DFFPOSX1 _21214_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf123),
    .D(_4631_),
    .Q(\datapath.registers.1226[16] [11])
);

DFFPOSX1 _21215_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf122),
    .D(_4632_),
    .Q(\datapath.registers.1226[16] [12])
);

DFFPOSX1 _21216_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf121),
    .D(_4633_),
    .Q(\datapath.registers.1226[16] [13])
);

DFFPOSX1 _21217_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf120),
    .D(_4634_),
    .Q(\datapath.registers.1226[16] [14])
);

DFFPOSX1 _21218_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf119),
    .D(_4635_),
    .Q(\datapath.registers.1226[16] [15])
);

DFFPOSX1 _21219_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf118),
    .D(_4636_),
    .Q(\datapath.registers.1226[16] [16])
);

DFFPOSX1 _21220_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf117),
    .D(_4637_),
    .Q(\datapath.registers.1226[16] [17])
);

DFFPOSX1 _21221_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf116),
    .D(_4638_),
    .Q(\datapath.registers.1226[16] [18])
);

DFFPOSX1 _21222_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf115),
    .D(_4639_),
    .Q(\datapath.registers.1226[16] [19])
);

DFFPOSX1 _21223_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf114),
    .D(_4641_),
    .Q(\datapath.registers.1226[16] [20])
);

DFFPOSX1 _21224_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf113),
    .D(_4642_),
    .Q(\datapath.registers.1226[16] [21])
);

DFFPOSX1 _21225_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf112),
    .D(_4643_),
    .Q(\datapath.registers.1226[16] [22])
);

DFFPOSX1 _21226_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf111),
    .D(_4644_),
    .Q(\datapath.registers.1226[16] [23])
);

DFFPOSX1 _21227_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf110),
    .D(_4645_),
    .Q(\datapath.registers.1226[16] [24])
);

DFFPOSX1 _21228_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf109),
    .D(_4646_),
    .Q(\datapath.registers.1226[16] [25])
);

DFFPOSX1 _21229_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf108),
    .D(_4647_),
    .Q(\datapath.registers.1226[16] [26])
);

DFFPOSX1 _21230_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf107),
    .D(_4648_),
    .Q(\datapath.registers.1226[16] [27])
);

DFFPOSX1 _21231_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf106),
    .D(_4649_),
    .Q(\datapath.registers.1226[16] [28])
);

DFFPOSX1 _21232_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf105),
    .D(_4650_),
    .Q(\datapath.registers.1226[16] [29])
);

DFFPOSX1 _21233_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf104),
    .D(_4652_),
    .Q(\datapath.registers.1226[16] [30])
);

DFFPOSX1 _21234_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf103),
    .D(_4653_),
    .Q(\datapath.registers.1226[16] [31])
);

DFFPOSX1 _21235_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf102),
    .D(_5237_),
    .Q(\datapath.registers.1226[4] [0])
);

DFFPOSX1 _21236_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf101),
    .D(_5248_),
    .Q(\datapath.registers.1226[4] [1])
);

DFFPOSX1 _21237_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf100),
    .D(_5259_),
    .Q(\datapath.registers.1226[4] [2])
);

DFFPOSX1 _21238_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf99),
    .D(_5262_),
    .Q(\datapath.registers.1226[4] [3])
);

DFFPOSX1 _21239_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf98),
    .D(_5263_),
    .Q(\datapath.registers.1226[4] [4])
);

DFFPOSX1 _21240_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf97),
    .D(_5264_),
    .Q(\datapath.registers.1226[4] [5])
);

DFFPOSX1 _21241_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf96),
    .D(_5265_),
    .Q(\datapath.registers.1226[4] [6])
);

DFFPOSX1 _21242_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf95),
    .D(_5266_),
    .Q(\datapath.registers.1226[4] [7])
);

DFFPOSX1 _21243_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf94),
    .D(_5267_),
    .Q(\datapath.registers.1226[4] [8])
);

DFFPOSX1 _21244_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf93),
    .D(_5268_),
    .Q(\datapath.registers.1226[4] [9])
);

DFFPOSX1 _21245_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf92),
    .D(_5238_),
    .Q(\datapath.registers.1226[4] [10])
);

DFFPOSX1 _21246_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf91),
    .D(_5239_),
    .Q(\datapath.registers.1226[4] [11])
);

DFFPOSX1 _21247_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf90),
    .D(_5240_),
    .Q(\datapath.registers.1226[4] [12])
);

DFFPOSX1 _21248_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf89),
    .D(_5241_),
    .Q(\datapath.registers.1226[4] [13])
);

DFFPOSX1 _21249_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf88),
    .D(_5242_),
    .Q(\datapath.registers.1226[4] [14])
);

DFFPOSX1 _21250_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf87),
    .D(_5243_),
    .Q(\datapath.registers.1226[4] [15])
);

DFFPOSX1 _21251_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf86),
    .D(_5244_),
    .Q(\datapath.registers.1226[4] [16])
);

DFFPOSX1 _21252_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf85),
    .D(_5245_),
    .Q(\datapath.registers.1226[4] [17])
);

DFFPOSX1 _21253_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf84),
    .D(_5246_),
    .Q(\datapath.registers.1226[4] [18])
);

DFFPOSX1 _21254_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf83),
    .D(_5247_),
    .Q(\datapath.registers.1226[4] [19])
);

DFFPOSX1 _21255_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf82),
    .D(_5249_),
    .Q(\datapath.registers.1226[4] [20])
);

DFFPOSX1 _21256_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf81),
    .D(_5250_),
    .Q(\datapath.registers.1226[4] [21])
);

DFFPOSX1 _21257_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf80),
    .D(_5251_),
    .Q(\datapath.registers.1226[4] [22])
);

DFFPOSX1 _21258_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf79),
    .D(_5252_),
    .Q(\datapath.registers.1226[4] [23])
);

DFFPOSX1 _21259_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf78),
    .D(_5253_),
    .Q(\datapath.registers.1226[4] [24])
);

DFFPOSX1 _21260_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf77),
    .D(_5254_),
    .Q(\datapath.registers.1226[4] [25])
);

DFFPOSX1 _21261_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf76),
    .D(_5255_),
    .Q(\datapath.registers.1226[4] [26])
);

DFFPOSX1 _21262_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf75),
    .D(_5256_),
    .Q(\datapath.registers.1226[4] [27])
);

DFFPOSX1 _21263_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf74),
    .D(_5257_),
    .Q(\datapath.registers.1226[4] [28])
);

DFFPOSX1 _21264_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf73),
    .D(_5258_),
    .Q(\datapath.registers.1226[4] [29])
);

DFFPOSX1 _21265_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf72),
    .D(_5260_),
    .Q(\datapath.registers.1226[4] [30])
);

DFFPOSX1 _21266_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf71),
    .D(_5261_),
    .Q(\datapath.registers.1226[4] [31])
);

DFFPOSX1 _21267_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf70),
    .D(_5365_),
    .Q(\datapath.registers.1226[8] [0])
);

DFFPOSX1 _21268_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf69),
    .D(_5376_),
    .Q(\datapath.registers.1226[8] [1])
);

DFFPOSX1 _21269_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf68),
    .D(_5387_),
    .Q(\datapath.registers.1226[8] [2])
);

DFFPOSX1 _21270_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf67),
    .D(_5390_),
    .Q(\datapath.registers.1226[8] [3])
);

DFFPOSX1 _21271_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf66),
    .D(_5391_),
    .Q(\datapath.registers.1226[8] [4])
);

DFFPOSX1 _21272_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf65),
    .D(_5392_),
    .Q(\datapath.registers.1226[8] [5])
);

DFFPOSX1 _21273_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf64),
    .D(_5393_),
    .Q(\datapath.registers.1226[8] [6])
);

DFFPOSX1 _21274_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf63),
    .D(_5394_),
    .Q(\datapath.registers.1226[8] [7])
);

DFFPOSX1 _21275_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf62),
    .D(_5395_),
    .Q(\datapath.registers.1226[8] [8])
);

DFFPOSX1 _21276_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf61),
    .D(_5396_),
    .Q(\datapath.registers.1226[8] [9])
);

DFFPOSX1 _21277_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf60),
    .D(_5366_),
    .Q(\datapath.registers.1226[8] [10])
);

DFFPOSX1 _21278_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf59),
    .D(_5367_),
    .Q(\datapath.registers.1226[8] [11])
);

DFFPOSX1 _21279_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf58),
    .D(_5368_),
    .Q(\datapath.registers.1226[8] [12])
);

DFFPOSX1 _21280_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf57),
    .D(_5369_),
    .Q(\datapath.registers.1226[8] [13])
);

DFFPOSX1 _21281_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf56),
    .D(_5370_),
    .Q(\datapath.registers.1226[8] [14])
);

DFFPOSX1 _21282_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf55),
    .D(_5371_),
    .Q(\datapath.registers.1226[8] [15])
);

DFFPOSX1 _21283_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf54),
    .D(_5372_),
    .Q(\datapath.registers.1226[8] [16])
);

DFFPOSX1 _21284_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf53),
    .D(_5373_),
    .Q(\datapath.registers.1226[8] [17])
);

DFFPOSX1 _21285_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf52),
    .D(_5374_),
    .Q(\datapath.registers.1226[8] [18])
);

DFFPOSX1 _21286_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf51),
    .D(_5375_),
    .Q(\datapath.registers.1226[8] [19])
);

DFFPOSX1 _21287_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf50),
    .D(_5377_),
    .Q(\datapath.registers.1226[8] [20])
);

DFFPOSX1 _21288_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf49),
    .D(_5378_),
    .Q(\datapath.registers.1226[8] [21])
);

DFFPOSX1 _21289_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf48),
    .D(_5379_),
    .Q(\datapath.registers.1226[8] [22])
);

DFFPOSX1 _21290_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf47),
    .D(_5380_),
    .Q(\datapath.registers.1226[8] [23])
);

DFFPOSX1 _21291_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf46),
    .D(_5381_),
    .Q(\datapath.registers.1226[8] [24])
);

DFFPOSX1 _21292_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf45),
    .D(_5382_),
    .Q(\datapath.registers.1226[8] [25])
);

DFFPOSX1 _21293_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf44),
    .D(_5383_),
    .Q(\datapath.registers.1226[8] [26])
);

DFFPOSX1 _21294_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf43),
    .D(_5384_),
    .Q(\datapath.registers.1226[8] [27])
);

DFFPOSX1 _21295_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf42),
    .D(_5385_),
    .Q(\datapath.registers.1226[8] [28])
);

DFFPOSX1 _21296_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf41),
    .D(_5386_),
    .Q(\datapath.registers.1226[8] [29])
);

DFFPOSX1 _21297_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf40),
    .D(_5388_),
    .Q(\datapath.registers.1226[8] [30])
);

DFFPOSX1 _21298_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf39),
    .D(_5389_),
    .Q(\datapath.registers.1226[8] [31])
);

DFFPOSX1 _21299_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf38),
    .D(_4533_),
    .Q(\datapath.registers.1226[13] [0])
);

DFFPOSX1 _21300_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf37),
    .D(_4544_),
    .Q(\datapath.registers.1226[13] [1])
);

DFFPOSX1 _21301_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf36),
    .D(_4555_),
    .Q(\datapath.registers.1226[13] [2])
);

DFFPOSX1 _21302_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf35),
    .D(_4558_),
    .Q(\datapath.registers.1226[13] [3])
);

DFFPOSX1 _21303_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf34),
    .D(_4559_),
    .Q(\datapath.registers.1226[13] [4])
);

DFFPOSX1 _21304_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf33),
    .D(_4560_),
    .Q(\datapath.registers.1226[13] [5])
);

DFFPOSX1 _21305_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf32),
    .D(_4561_),
    .Q(\datapath.registers.1226[13] [6])
);

DFFPOSX1 _21306_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf31),
    .D(_4562_),
    .Q(\datapath.registers.1226[13] [7])
);

DFFPOSX1 _21307_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf30),
    .D(_4563_),
    .Q(\datapath.registers.1226[13] [8])
);

DFFPOSX1 _21308_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf29),
    .D(_4564_),
    .Q(\datapath.registers.1226[13] [9])
);

DFFPOSX1 _21309_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf28),
    .D(_4534_),
    .Q(\datapath.registers.1226[13] [10])
);

DFFPOSX1 _21310_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf27),
    .D(_4535_),
    .Q(\datapath.registers.1226[13] [11])
);

DFFPOSX1 _21311_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf26),
    .D(_4536_),
    .Q(\datapath.registers.1226[13] [12])
);

DFFPOSX1 _21312_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf25),
    .D(_4537_),
    .Q(\datapath.registers.1226[13] [13])
);

DFFPOSX1 _21313_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf24),
    .D(_4538_),
    .Q(\datapath.registers.1226[13] [14])
);

DFFPOSX1 _21314_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf23),
    .D(_4539_),
    .Q(\datapath.registers.1226[13] [15])
);

DFFPOSX1 _21315_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf22),
    .D(_4540_),
    .Q(\datapath.registers.1226[13] [16])
);

DFFPOSX1 _21316_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf21),
    .D(_4541_),
    .Q(\datapath.registers.1226[13] [17])
);

DFFPOSX1 _21317_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf20),
    .D(_4542_),
    .Q(\datapath.registers.1226[13] [18])
);

DFFPOSX1 _21318_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf19),
    .D(_4543_),
    .Q(\datapath.registers.1226[13] [19])
);

DFFPOSX1 _21319_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf18),
    .D(_4545_),
    .Q(\datapath.registers.1226[13] [20])
);

DFFPOSX1 _21320_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf17),
    .D(_4546_),
    .Q(\datapath.registers.1226[13] [21])
);

DFFPOSX1 _21321_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf16),
    .D(_4547_),
    .Q(\datapath.registers.1226[13] [22])
);

DFFPOSX1 _21322_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf15),
    .D(_4548_),
    .Q(\datapath.registers.1226[13] [23])
);

DFFPOSX1 _21323_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf14),
    .D(_4549_),
    .Q(\datapath.registers.1226[13] [24])
);

DFFPOSX1 _21324_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf13),
    .D(_4550_),
    .Q(\datapath.registers.1226[13] [25])
);

DFFPOSX1 _21325_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf12),
    .D(_4551_),
    .Q(\datapath.registers.1226[13] [26])
);

DFFPOSX1 _21326_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf11),
    .D(_4552_),
    .Q(\datapath.registers.1226[13] [27])
);

DFFPOSX1 _21327_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf10),
    .D(_4553_),
    .Q(\datapath.registers.1226[13] [28])
);

DFFPOSX1 _21328_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf9),
    .D(_4554_),
    .Q(\datapath.registers.1226[13] [29])
);

DFFPOSX1 _21329_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf8),
    .D(_4556_),
    .Q(\datapath.registers.1226[13] [30])
);

DFFPOSX1 _21330_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf7),
    .D(_4557_),
    .Q(\datapath.registers.1226[13] [31])
);

DFFPOSX1 _21331_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf6),
    .D(_4757_),
    .Q(\datapath.registers.1226[1] [0])
);

DFFPOSX1 _21332_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf5),
    .D(_4768_),
    .Q(\datapath.registers.1226[1] [1])
);

DFFPOSX1 _21333_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf4),
    .D(_4779_),
    .Q(\datapath.registers.1226[1] [2])
);

DFFPOSX1 _21334_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf3),
    .D(_4782_),
    .Q(\datapath.registers.1226[1] [3])
);

DFFPOSX1 _21335_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf2),
    .D(_4783_),
    .Q(\datapath.registers.1226[1] [4])
);

DFFPOSX1 _21336_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf1),
    .D(_4784_),
    .Q(\datapath.registers.1226[1] [5])
);

DFFPOSX1 _21337_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf0),
    .D(_4785_),
    .Q(\datapath.registers.1226[1] [6])
);

DFFPOSX1 _21338_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf153),
    .D(_4786_),
    .Q(\datapath.registers.1226[1] [7])
);

DFFPOSX1 _21339_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf152),
    .D(_4787_),
    .Q(\datapath.registers.1226[1] [8])
);

DFFPOSX1 _21340_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf151),
    .D(_4788_),
    .Q(\datapath.registers.1226[1] [9])
);

DFFPOSX1 _21341_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf150),
    .D(_4758_),
    .Q(\datapath.registers.1226[1] [10])
);

DFFPOSX1 _21342_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf149),
    .D(_4759_),
    .Q(\datapath.registers.1226[1] [11])
);

DFFPOSX1 _21343_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf148),
    .D(_4760_),
    .Q(\datapath.registers.1226[1] [12])
);

DFFPOSX1 _21344_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf147),
    .D(_4761_),
    .Q(\datapath.registers.1226[1] [13])
);

DFFPOSX1 _21345_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf146),
    .D(_4762_),
    .Q(\datapath.registers.1226[1] [14])
);

DFFPOSX1 _21346_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf145),
    .D(_4763_),
    .Q(\datapath.registers.1226[1] [15])
);

DFFPOSX1 _21347_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf144),
    .D(_4764_),
    .Q(\datapath.registers.1226[1] [16])
);

DFFPOSX1 _21348_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf143),
    .D(_4765_),
    .Q(\datapath.registers.1226[1] [17])
);

DFFPOSX1 _21349_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf142),
    .D(_4766_),
    .Q(\datapath.registers.1226[1] [18])
);

DFFPOSX1 _21350_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf141),
    .D(_4767_),
    .Q(\datapath.registers.1226[1] [19])
);

DFFPOSX1 _21351_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf140),
    .D(_4769_),
    .Q(\datapath.registers.1226[1] [20])
);

DFFPOSX1 _21352_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf139),
    .D(_4770_),
    .Q(\datapath.registers.1226[1] [21])
);

DFFPOSX1 _21353_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf138),
    .D(_4771_),
    .Q(\datapath.registers.1226[1] [22])
);

DFFPOSX1 _21354_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf137),
    .D(_4772_),
    .Q(\datapath.registers.1226[1] [23])
);

DFFPOSX1 _21355_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf136),
    .D(_4773_),
    .Q(\datapath.registers.1226[1] [24])
);

DFFPOSX1 _21356_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf135),
    .D(_4774_),
    .Q(\datapath.registers.1226[1] [25])
);

DFFPOSX1 _21357_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf134),
    .D(_4775_),
    .Q(\datapath.registers.1226[1] [26])
);

DFFPOSX1 _21358_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf133),
    .D(_4776_),
    .Q(\datapath.registers.1226[1] [27])
);

DFFPOSX1 _21359_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf132),
    .D(_4777_),
    .Q(\datapath.registers.1226[1] [28])
);

DFFPOSX1 _21360_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf131),
    .D(_4778_),
    .Q(\datapath.registers.1226[1] [29])
);

DFFPOSX1 _21361_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf130),
    .D(_4780_),
    .Q(\datapath.registers.1226[1] [30])
);

DFFPOSX1 _21362_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf129),
    .D(_4781_),
    .Q(\datapath.registers.1226[1] [31])
);

DFFPOSX1 _21363_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf128),
    .D(_4917_),
    .Q(\datapath.registers.1226[24] [0])
);

DFFPOSX1 _21364_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf127),
    .D(_4928_),
    .Q(\datapath.registers.1226[24] [1])
);

DFFPOSX1 _21365_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf126),
    .D(_4939_),
    .Q(\datapath.registers.1226[24] [2])
);

DFFPOSX1 _21366_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf125),
    .D(_4942_),
    .Q(\datapath.registers.1226[24] [3])
);

DFFPOSX1 _21367_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf124),
    .D(_4943_),
    .Q(\datapath.registers.1226[24] [4])
);

DFFPOSX1 _21368_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf123),
    .D(_4944_),
    .Q(\datapath.registers.1226[24] [5])
);

DFFPOSX1 _21369_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf122),
    .D(_4945_),
    .Q(\datapath.registers.1226[24] [6])
);

DFFPOSX1 _21370_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf121),
    .D(_4946_),
    .Q(\datapath.registers.1226[24] [7])
);

DFFPOSX1 _21371_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf120),
    .D(_4947_),
    .Q(\datapath.registers.1226[24] [8])
);

DFFPOSX1 _21372_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf119),
    .D(_4948_),
    .Q(\datapath.registers.1226[24] [9])
);

DFFPOSX1 _21373_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf118),
    .D(_4918_),
    .Q(\datapath.registers.1226[24] [10])
);

DFFPOSX1 _21374_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf117),
    .D(_4919_),
    .Q(\datapath.registers.1226[24] [11])
);

DFFPOSX1 _21375_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf116),
    .D(_4920_),
    .Q(\datapath.registers.1226[24] [12])
);

DFFPOSX1 _21376_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf115),
    .D(_4921_),
    .Q(\datapath.registers.1226[24] [13])
);

DFFPOSX1 _21377_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf114),
    .D(_4922_),
    .Q(\datapath.registers.1226[24] [14])
);

DFFPOSX1 _21378_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf113),
    .D(_4923_),
    .Q(\datapath.registers.1226[24] [15])
);

DFFPOSX1 _21379_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf112),
    .D(_4924_),
    .Q(\datapath.registers.1226[24] [16])
);

DFFPOSX1 _21380_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf111),
    .D(_4925_),
    .Q(\datapath.registers.1226[24] [17])
);

DFFPOSX1 _21381_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf110),
    .D(_4926_),
    .Q(\datapath.registers.1226[24] [18])
);

DFFPOSX1 _21382_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf109),
    .D(_4927_),
    .Q(\datapath.registers.1226[24] [19])
);

DFFPOSX1 _21383_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf108),
    .D(_4929_),
    .Q(\datapath.registers.1226[24] [20])
);

DFFPOSX1 _21384_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf107),
    .D(_4930_),
    .Q(\datapath.registers.1226[24] [21])
);

DFFPOSX1 _21385_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf106),
    .D(_4931_),
    .Q(\datapath.registers.1226[24] [22])
);

DFFPOSX1 _21386_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf105),
    .D(_4932_),
    .Q(\datapath.registers.1226[24] [23])
);

DFFPOSX1 _21387_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf104),
    .D(_4933_),
    .Q(\datapath.registers.1226[24] [24])
);

DFFPOSX1 _21388_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf103),
    .D(_4934_),
    .Q(\datapath.registers.1226[24] [25])
);

DFFPOSX1 _21389_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf102),
    .D(_4935_),
    .Q(\datapath.registers.1226[24] [26])
);

DFFPOSX1 _21390_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf101),
    .D(_4936_),
    .Q(\datapath.registers.1226[24] [27])
);

DFFPOSX1 _21391_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf100),
    .D(_4937_),
    .Q(\datapath.registers.1226[24] [28])
);

DFFPOSX1 _21392_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf99),
    .D(_4938_),
    .Q(\datapath.registers.1226[24] [29])
);

DFFPOSX1 _21393_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf98),
    .D(_4940_),
    .Q(\datapath.registers.1226[24] [30])
);

DFFPOSX1 _21394_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf97),
    .D(_4941_),
    .Q(\datapath.registers.1226[24] [31])
);

DFFPOSX1 _21395_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf96),
    .D(_4501_),
    .Q(\datapath.registers.1226[12] [0])
);

DFFPOSX1 _21396_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf95),
    .D(_4512_),
    .Q(\datapath.registers.1226[12] [1])
);

DFFPOSX1 _21397_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf94),
    .D(_4523_),
    .Q(\datapath.registers.1226[12] [2])
);

DFFPOSX1 _21398_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf93),
    .D(_4526_),
    .Q(\datapath.registers.1226[12] [3])
);

DFFPOSX1 _21399_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf92),
    .D(_4527_),
    .Q(\datapath.registers.1226[12] [4])
);

DFFPOSX1 _21400_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf91),
    .D(_4528_),
    .Q(\datapath.registers.1226[12] [5])
);

DFFPOSX1 _21401_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf90),
    .D(_4529_),
    .Q(\datapath.registers.1226[12] [6])
);

DFFPOSX1 _21402_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf89),
    .D(_4530_),
    .Q(\datapath.registers.1226[12] [7])
);

DFFPOSX1 _21403_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf88),
    .D(_4531_),
    .Q(\datapath.registers.1226[12] [8])
);

DFFPOSX1 _21404_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf87),
    .D(_4532_),
    .Q(\datapath.registers.1226[12] [9])
);

DFFPOSX1 _21405_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf86),
    .D(_4502_),
    .Q(\datapath.registers.1226[12] [10])
);

DFFPOSX1 _21406_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf85),
    .D(_4503_),
    .Q(\datapath.registers.1226[12] [11])
);

DFFPOSX1 _21407_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf84),
    .D(_4504_),
    .Q(\datapath.registers.1226[12] [12])
);

DFFPOSX1 _21408_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf83),
    .D(_4505_),
    .Q(\datapath.registers.1226[12] [13])
);

DFFPOSX1 _21409_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf82),
    .D(_4506_),
    .Q(\datapath.registers.1226[12] [14])
);

DFFPOSX1 _21410_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf81),
    .D(_4507_),
    .Q(\datapath.registers.1226[12] [15])
);

DFFPOSX1 _21411_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf80),
    .D(_4508_),
    .Q(\datapath.registers.1226[12] [16])
);

DFFPOSX1 _21412_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf79),
    .D(_4509_),
    .Q(\datapath.registers.1226[12] [17])
);

DFFPOSX1 _21413_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf78),
    .D(_4510_),
    .Q(\datapath.registers.1226[12] [18])
);

DFFPOSX1 _21414_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf77),
    .D(_4511_),
    .Q(\datapath.registers.1226[12] [19])
);

DFFPOSX1 _21415_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf76),
    .D(_4513_),
    .Q(\datapath.registers.1226[12] [20])
);

DFFPOSX1 _21416_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf75),
    .D(_4514_),
    .Q(\datapath.registers.1226[12] [21])
);

DFFPOSX1 _21417_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf74),
    .D(_4515_),
    .Q(\datapath.registers.1226[12] [22])
);

DFFPOSX1 _21418_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf73),
    .D(_4516_),
    .Q(\datapath.registers.1226[12] [23])
);

DFFPOSX1 _21419_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf72),
    .D(_4517_),
    .Q(\datapath.registers.1226[12] [24])
);

DFFPOSX1 _21420_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf71),
    .D(_4518_),
    .Q(\datapath.registers.1226[12] [25])
);

DFFPOSX1 _21421_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf70),
    .D(_4519_),
    .Q(\datapath.registers.1226[12] [26])
);

DFFPOSX1 _21422_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf69),
    .D(_4520_),
    .Q(\datapath.registers.1226[12] [27])
);

DFFPOSX1 _21423_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf68),
    .D(_4521_),
    .Q(\datapath.registers.1226[12] [28])
);

DFFPOSX1 _21424_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf67),
    .D(_4522_),
    .Q(\datapath.registers.1226[12] [29])
);

DFFPOSX1 _21425_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf66),
    .D(_4524_),
    .Q(\datapath.registers.1226[12] [30])
);

DFFPOSX1 _21426_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf65),
    .D(_4525_),
    .Q(\datapath.registers.1226[12] [31])
);

DFFPOSX1 _21427_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf64),
    .D(_5269_),
    .Q(\datapath.registers.1226[5] [0])
);

DFFPOSX1 _21428_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf63),
    .D(_5280_),
    .Q(\datapath.registers.1226[5] [1])
);

DFFPOSX1 _21429_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf62),
    .D(_5291_),
    .Q(\datapath.registers.1226[5] [2])
);

DFFPOSX1 _21430_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf61),
    .D(_5294_),
    .Q(\datapath.registers.1226[5] [3])
);

DFFPOSX1 _21431_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf60),
    .D(_5295_),
    .Q(\datapath.registers.1226[5] [4])
);

DFFPOSX1 _21432_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf59),
    .D(_5296_),
    .Q(\datapath.registers.1226[5] [5])
);

DFFPOSX1 _21433_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf58),
    .D(_5297_),
    .Q(\datapath.registers.1226[5] [6])
);

DFFPOSX1 _21434_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf57),
    .D(_5298_),
    .Q(\datapath.registers.1226[5] [7])
);

DFFPOSX1 _21435_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf56),
    .D(_5299_),
    .Q(\datapath.registers.1226[5] [8])
);

DFFPOSX1 _21436_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf55),
    .D(_5300_),
    .Q(\datapath.registers.1226[5] [9])
);

DFFPOSX1 _21437_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf54),
    .D(_5270_),
    .Q(\datapath.registers.1226[5] [10])
);

DFFPOSX1 _21438_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf53),
    .D(_5271_),
    .Q(\datapath.registers.1226[5] [11])
);

DFFPOSX1 _21439_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf52),
    .D(_5272_),
    .Q(\datapath.registers.1226[5] [12])
);

DFFPOSX1 _21440_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf51),
    .D(_5273_),
    .Q(\datapath.registers.1226[5] [13])
);

DFFPOSX1 _21441_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf50),
    .D(_5274_),
    .Q(\datapath.registers.1226[5] [14])
);

DFFPOSX1 _21442_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf49),
    .D(_5275_),
    .Q(\datapath.registers.1226[5] [15])
);

DFFPOSX1 _21443_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf48),
    .D(_5276_),
    .Q(\datapath.registers.1226[5] [16])
);

DFFPOSX1 _21444_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf47),
    .D(_5277_),
    .Q(\datapath.registers.1226[5] [17])
);

DFFPOSX1 _21445_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf46),
    .D(_5278_),
    .Q(\datapath.registers.1226[5] [18])
);

DFFPOSX1 _21446_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf45),
    .D(_5279_),
    .Q(\datapath.registers.1226[5] [19])
);

DFFPOSX1 _21447_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf44),
    .D(_5281_),
    .Q(\datapath.registers.1226[5] [20])
);

DFFPOSX1 _21448_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf43),
    .D(_5282_),
    .Q(\datapath.registers.1226[5] [21])
);

DFFPOSX1 _21449_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf42),
    .D(_5283_),
    .Q(\datapath.registers.1226[5] [22])
);

DFFPOSX1 _21450_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf41),
    .D(_5284_),
    .Q(\datapath.registers.1226[5] [23])
);

DFFPOSX1 _21451_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf40),
    .D(_5285_),
    .Q(\datapath.registers.1226[5] [24])
);

DFFPOSX1 _21452_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf39),
    .D(_5286_),
    .Q(\datapath.registers.1226[5] [25])
);

DFFPOSX1 _21453_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf38),
    .D(_5287_),
    .Q(\datapath.registers.1226[5] [26])
);

DFFPOSX1 _21454_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf37),
    .D(_5288_),
    .Q(\datapath.registers.1226[5] [27])
);

DFFPOSX1 _21455_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf36),
    .D(_5289_),
    .Q(\datapath.registers.1226[5] [28])
);

DFFPOSX1 _21456_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf35),
    .D(_5290_),
    .Q(\datapath.registers.1226[5] [29])
);

DFFPOSX1 _21457_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf34),
    .D(_5292_),
    .Q(\datapath.registers.1226[5] [30])
);

DFFPOSX1 _21458_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf33),
    .D(_5293_),
    .Q(\datapath.registers.1226[5] [31])
);

DFFPOSX1 _21459_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf32),
    .D(_4981_),
    .Q(\datapath.registers.1226[26] [0])
);

DFFPOSX1 _21460_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf31),
    .D(_4992_),
    .Q(\datapath.registers.1226[26] [1])
);

DFFPOSX1 _21461_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf30),
    .D(_5003_),
    .Q(\datapath.registers.1226[26] [2])
);

DFFPOSX1 _21462_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf29),
    .D(_5006_),
    .Q(\datapath.registers.1226[26] [3])
);

DFFPOSX1 _21463_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf28),
    .D(_5007_),
    .Q(\datapath.registers.1226[26] [4])
);

DFFPOSX1 _21464_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf27),
    .D(_5008_),
    .Q(\datapath.registers.1226[26] [5])
);

DFFPOSX1 _21465_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf26),
    .D(_5009_),
    .Q(\datapath.registers.1226[26] [6])
);

DFFPOSX1 _21466_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf25),
    .D(_5010_),
    .Q(\datapath.registers.1226[26] [7])
);

DFFPOSX1 _21467_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf24),
    .D(_5011_),
    .Q(\datapath.registers.1226[26] [8])
);

DFFPOSX1 _21468_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf23),
    .D(_5012_),
    .Q(\datapath.registers.1226[26] [9])
);

DFFPOSX1 _21469_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf22),
    .D(_4982_),
    .Q(\datapath.registers.1226[26] [10])
);

DFFPOSX1 _21470_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf21),
    .D(_4983_),
    .Q(\datapath.registers.1226[26] [11])
);

DFFPOSX1 _21471_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf20),
    .D(_4984_),
    .Q(\datapath.registers.1226[26] [12])
);

DFFPOSX1 _21472_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf19),
    .D(_4985_),
    .Q(\datapath.registers.1226[26] [13])
);

DFFPOSX1 _21473_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf18),
    .D(_4986_),
    .Q(\datapath.registers.1226[26] [14])
);

DFFPOSX1 _21474_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf17),
    .D(_4987_),
    .Q(\datapath.registers.1226[26] [15])
);

DFFPOSX1 _21475_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf16),
    .D(_4988_),
    .Q(\datapath.registers.1226[26] [16])
);

DFFPOSX1 _21476_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf15),
    .D(_4989_),
    .Q(\datapath.registers.1226[26] [17])
);

DFFPOSX1 _21477_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf14),
    .D(_4990_),
    .Q(\datapath.registers.1226[26] [18])
);

DFFPOSX1 _21478_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf13),
    .D(_4991_),
    .Q(\datapath.registers.1226[26] [19])
);

DFFPOSX1 _21479_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf12),
    .D(_4993_),
    .Q(\datapath.registers.1226[26] [20])
);

DFFPOSX1 _21480_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf11),
    .D(_4994_),
    .Q(\datapath.registers.1226[26] [21])
);

DFFPOSX1 _21481_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf10),
    .D(_4995_),
    .Q(\datapath.registers.1226[26] [22])
);

DFFPOSX1 _21482_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf9),
    .D(_4996_),
    .Q(\datapath.registers.1226[26] [23])
);

DFFPOSX1 _21483_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf8),
    .D(_4997_),
    .Q(\datapath.registers.1226[26] [24])
);

DFFPOSX1 _21484_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf7),
    .D(_4998_),
    .Q(\datapath.registers.1226[26] [25])
);

DFFPOSX1 _21485_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf6),
    .D(_4999_),
    .Q(\datapath.registers.1226[26] [26])
);

DFFPOSX1 _21486_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf5),
    .D(_5000_),
    .Q(\datapath.registers.1226[26] [27])
);

DFFPOSX1 _21487_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf4),
    .D(_5001_),
    .Q(\datapath.registers.1226[26] [28])
);

DFFPOSX1 _21488_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf3),
    .D(_5002_),
    .Q(\datapath.registers.1226[26] [29])
);

DFFPOSX1 _21489_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf2),
    .D(_5004_),
    .Q(\datapath.registers.1226[26] [30])
);

DFFPOSX1 _21490_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf1),
    .D(_5005_),
    .Q(\datapath.registers.1226[26] [31])
);

DFFPOSX1 _21491_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf0),
    .D(_4725_),
    .Q(\datapath.registers.1226[19] [0])
);

DFFPOSX1 _21492_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf153),
    .D(_4736_),
    .Q(\datapath.registers.1226[19] [1])
);

DFFPOSX1 _21493_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf152),
    .D(_4747_),
    .Q(\datapath.registers.1226[19] [2])
);

DFFPOSX1 _21494_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf151),
    .D(_4750_),
    .Q(\datapath.registers.1226[19] [3])
);

DFFPOSX1 _21495_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf150),
    .D(_4751_),
    .Q(\datapath.registers.1226[19] [4])
);

DFFPOSX1 _21496_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf149),
    .D(_4752_),
    .Q(\datapath.registers.1226[19] [5])
);

DFFPOSX1 _21497_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf148),
    .D(_4753_),
    .Q(\datapath.registers.1226[19] [6])
);

DFFPOSX1 _21498_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf147),
    .D(_4754_),
    .Q(\datapath.registers.1226[19] [7])
);

DFFPOSX1 _21499_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf146),
    .D(_4755_),
    .Q(\datapath.registers.1226[19] [8])
);

DFFPOSX1 _21500_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf145),
    .D(_4756_),
    .Q(\datapath.registers.1226[19] [9])
);

DFFPOSX1 _21501_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf144),
    .D(_4726_),
    .Q(\datapath.registers.1226[19] [10])
);

DFFPOSX1 _21502_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf143),
    .D(_4727_),
    .Q(\datapath.registers.1226[19] [11])
);

DFFPOSX1 _21503_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf142),
    .D(_4728_),
    .Q(\datapath.registers.1226[19] [12])
);

DFFPOSX1 _21504_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf141),
    .D(_4729_),
    .Q(\datapath.registers.1226[19] [13])
);

DFFPOSX1 _21505_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf140),
    .D(_4730_),
    .Q(\datapath.registers.1226[19] [14])
);

DFFPOSX1 _21506_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf139),
    .D(_4731_),
    .Q(\datapath.registers.1226[19] [15])
);

DFFPOSX1 _21507_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf138),
    .D(_4732_),
    .Q(\datapath.registers.1226[19] [16])
);

DFFPOSX1 _21508_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf137),
    .D(_4733_),
    .Q(\datapath.registers.1226[19] [17])
);

DFFPOSX1 _21509_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf136),
    .D(_4734_),
    .Q(\datapath.registers.1226[19] [18])
);

DFFPOSX1 _21510_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf135),
    .D(_4735_),
    .Q(\datapath.registers.1226[19] [19])
);

DFFPOSX1 _21511_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf134),
    .D(_4737_),
    .Q(\datapath.registers.1226[19] [20])
);

DFFPOSX1 _21512_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf133),
    .D(_4738_),
    .Q(\datapath.registers.1226[19] [21])
);

DFFPOSX1 _21513_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf132),
    .D(_4739_),
    .Q(\datapath.registers.1226[19] [22])
);

DFFPOSX1 _21514_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf131),
    .D(_4740_),
    .Q(\datapath.registers.1226[19] [23])
);

DFFPOSX1 _21515_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf130),
    .D(_4741_),
    .Q(\datapath.registers.1226[19] [24])
);

DFFPOSX1 _21516_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf129),
    .D(_4742_),
    .Q(\datapath.registers.1226[19] [25])
);

DFFPOSX1 _21517_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf128),
    .D(_4743_),
    .Q(\datapath.registers.1226[19] [26])
);

DFFPOSX1 _21518_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf127),
    .D(_4744_),
    .Q(\datapath.registers.1226[19] [27])
);

DFFPOSX1 _21519_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf126),
    .D(_4745_),
    .Q(\datapath.registers.1226[19] [28])
);

DFFPOSX1 _21520_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf125),
    .D(_4746_),
    .Q(\datapath.registers.1226[19] [29])
);

DFFPOSX1 _21521_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf124),
    .D(_4748_),
    .Q(\datapath.registers.1226[19] [30])
);

DFFPOSX1 _21522_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf123),
    .D(_4749_),
    .Q(\datapath.registers.1226[19] [31])
);

DFFPOSX1 _21523_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf122),
    .D(_4405_),
    .Q(\datapath.registers.1226[0] [0])
);

DFFPOSX1 _21524_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf121),
    .D(_4416_),
    .Q(\datapath.registers.1226[0] [1])
);

DFFPOSX1 _21525_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf120),
    .D(_4427_),
    .Q(\datapath.registers.1226[0] [2])
);

DFFPOSX1 _21526_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf119),
    .D(_4430_),
    .Q(\datapath.registers.1226[0] [3])
);

DFFPOSX1 _21527_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf118),
    .D(_4431_),
    .Q(\datapath.registers.1226[0] [4])
);

DFFPOSX1 _21528_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf117),
    .D(_4432_),
    .Q(\datapath.registers.1226[0] [5])
);

DFFPOSX1 _21529_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf116),
    .D(_4433_),
    .Q(\datapath.registers.1226[0] [6])
);

DFFPOSX1 _21530_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf115),
    .D(_4434_),
    .Q(\datapath.registers.1226[0] [7])
);

DFFPOSX1 _21531_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf114),
    .D(_4435_),
    .Q(\datapath.registers.1226[0] [8])
);

DFFPOSX1 _21532_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf113),
    .D(_4436_),
    .Q(\datapath.registers.1226[0] [9])
);

DFFPOSX1 _21533_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf112),
    .D(_4406_),
    .Q(\datapath.registers.1226[0] [10])
);

DFFPOSX1 _21534_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf111),
    .D(_4407_),
    .Q(\datapath.registers.1226[0] [11])
);

DFFPOSX1 _21535_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf110),
    .D(_4408_),
    .Q(\datapath.registers.1226[0] [12])
);

DFFPOSX1 _21536_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf109),
    .D(_4409_),
    .Q(\datapath.registers.1226[0] [13])
);

DFFPOSX1 _21537_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf108),
    .D(_4410_),
    .Q(\datapath.registers.1226[0] [14])
);

DFFPOSX1 _21538_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf107),
    .D(_4411_),
    .Q(\datapath.registers.1226[0] [15])
);

DFFPOSX1 _21539_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf106),
    .D(_4412_),
    .Q(\datapath.registers.1226[0] [16])
);

DFFPOSX1 _21540_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf105),
    .D(_4413_),
    .Q(\datapath.registers.1226[0] [17])
);

DFFPOSX1 _21541_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf104),
    .D(_4414_),
    .Q(\datapath.registers.1226[0] [18])
);

DFFPOSX1 _21542_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf103),
    .D(_4415_),
    .Q(\datapath.registers.1226[0] [19])
);

DFFPOSX1 _21543_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf102),
    .D(_4417_),
    .Q(\datapath.registers.1226[0] [20])
);

DFFPOSX1 _21544_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf101),
    .D(_4418_),
    .Q(\datapath.registers.1226[0] [21])
);

DFFPOSX1 _21545_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf100),
    .D(_4419_),
    .Q(\datapath.registers.1226[0] [22])
);

DFFPOSX1 _21546_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf99),
    .D(_4420_),
    .Q(\datapath.registers.1226[0] [23])
);

DFFPOSX1 _21547_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf98),
    .D(_4421_),
    .Q(\datapath.registers.1226[0] [24])
);

DFFPOSX1 _21548_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf97),
    .D(_4422_),
    .Q(\datapath.registers.1226[0] [25])
);

DFFPOSX1 _21549_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf96),
    .D(_4423_),
    .Q(\datapath.registers.1226[0] [26])
);

DFFPOSX1 _21550_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf95),
    .D(_4424_),
    .Q(\datapath.registers.1226[0] [27])
);

DFFPOSX1 _21551_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf94),
    .D(_4425_),
    .Q(\datapath.registers.1226[0] [28])
);

DFFPOSX1 _21552_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf93),
    .D(_4426_),
    .Q(\datapath.registers.1226[0] [29])
);

DFFPOSX1 _21553_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf92),
    .D(_4428_),
    .Q(\datapath.registers.1226[0] [30])
);

DFFPOSX1 _21554_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf91),
    .D(_4429_),
    .Q(\datapath.registers.1226[0] [31])
);

DFFPOSX1 _21555_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf90),
    .D(_4693_),
    .Q(\datapath.registers.1226[18] [0])
);

DFFPOSX1 _21556_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf89),
    .D(_4704_),
    .Q(\datapath.registers.1226[18] [1])
);

DFFPOSX1 _21557_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf88),
    .D(_4715_),
    .Q(\datapath.registers.1226[18] [2])
);

DFFPOSX1 _21558_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf87),
    .D(_4718_),
    .Q(\datapath.registers.1226[18] [3])
);

DFFPOSX1 _21559_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf86),
    .D(_4719_),
    .Q(\datapath.registers.1226[18] [4])
);

DFFPOSX1 _21560_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf85),
    .D(_4720_),
    .Q(\datapath.registers.1226[18] [5])
);

DFFPOSX1 _21561_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf84),
    .D(_4721_),
    .Q(\datapath.registers.1226[18] [6])
);

DFFPOSX1 _21562_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf83),
    .D(_4722_),
    .Q(\datapath.registers.1226[18] [7])
);

DFFPOSX1 _21563_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf82),
    .D(_4723_),
    .Q(\datapath.registers.1226[18] [8])
);

DFFPOSX1 _21564_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf81),
    .D(_4724_),
    .Q(\datapath.registers.1226[18] [9])
);

DFFPOSX1 _21565_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf80),
    .D(_4694_),
    .Q(\datapath.registers.1226[18] [10])
);

DFFPOSX1 _21566_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf79),
    .D(_4695_),
    .Q(\datapath.registers.1226[18] [11])
);

DFFPOSX1 _21567_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf78),
    .D(_4696_),
    .Q(\datapath.registers.1226[18] [12])
);

DFFPOSX1 _21568_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf77),
    .D(_4697_),
    .Q(\datapath.registers.1226[18] [13])
);

DFFPOSX1 _21569_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf76),
    .D(_4698_),
    .Q(\datapath.registers.1226[18] [14])
);

DFFPOSX1 _21570_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf75),
    .D(_4699_),
    .Q(\datapath.registers.1226[18] [15])
);

DFFPOSX1 _21571_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf74),
    .D(_4700_),
    .Q(\datapath.registers.1226[18] [16])
);

DFFPOSX1 _21572_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf73),
    .D(_4701_),
    .Q(\datapath.registers.1226[18] [17])
);

DFFPOSX1 _21573_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf72),
    .D(_4702_),
    .Q(\datapath.registers.1226[18] [18])
);

DFFPOSX1 _21574_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf71),
    .D(_4703_),
    .Q(\datapath.registers.1226[18] [19])
);

DFFPOSX1 _21575_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf70),
    .D(_4705_),
    .Q(\datapath.registers.1226[18] [20])
);

DFFPOSX1 _21576_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf69),
    .D(_4706_),
    .Q(\datapath.registers.1226[18] [21])
);

DFFPOSX1 _21577_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf68),
    .D(_4707_),
    .Q(\datapath.registers.1226[18] [22])
);

DFFPOSX1 _21578_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf67),
    .D(_4708_),
    .Q(\datapath.registers.1226[18] [23])
);

DFFPOSX1 _21579_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf66),
    .D(_4709_),
    .Q(\datapath.registers.1226[18] [24])
);

DFFPOSX1 _21580_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf65),
    .D(_4710_),
    .Q(\datapath.registers.1226[18] [25])
);

DFFPOSX1 _21581_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf64),
    .D(_4711_),
    .Q(\datapath.registers.1226[18] [26])
);

DFFPOSX1 _21582_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf63),
    .D(_4712_),
    .Q(\datapath.registers.1226[18] [27])
);

DFFPOSX1 _21583_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf62),
    .D(_4713_),
    .Q(\datapath.registers.1226[18] [28])
);

DFFPOSX1 _21584_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf61),
    .D(_4714_),
    .Q(\datapath.registers.1226[18] [29])
);

DFFPOSX1 _21585_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf60),
    .D(_4716_),
    .Q(\datapath.registers.1226[18] [30])
);

DFFPOSX1 _21586_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf59),
    .D(_4717_),
    .Q(\datapath.registers.1226[18] [31])
);

DFFPOSX1 _21587_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf58),
    .D(_4661_),
    .Q(\datapath.registers.1226[17] [0])
);

DFFPOSX1 _21588_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf57),
    .D(_4672_),
    .Q(\datapath.registers.1226[17] [1])
);

DFFPOSX1 _21589_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf56),
    .D(_4683_),
    .Q(\datapath.registers.1226[17] [2])
);

DFFPOSX1 _21590_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf55),
    .D(_4686_),
    .Q(\datapath.registers.1226[17] [3])
);

DFFPOSX1 _21591_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf54),
    .D(_4687_),
    .Q(\datapath.registers.1226[17] [4])
);

DFFPOSX1 _21592_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf53),
    .D(_4688_),
    .Q(\datapath.registers.1226[17] [5])
);

DFFPOSX1 _21593_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf52),
    .D(_4689_),
    .Q(\datapath.registers.1226[17] [6])
);

DFFPOSX1 _21594_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf51),
    .D(_4690_),
    .Q(\datapath.registers.1226[17] [7])
);

DFFPOSX1 _21595_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf50),
    .D(_4691_),
    .Q(\datapath.registers.1226[17] [8])
);

DFFPOSX1 _21596_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf49),
    .D(_4692_),
    .Q(\datapath.registers.1226[17] [9])
);

DFFPOSX1 _21597_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf48),
    .D(_4662_),
    .Q(\datapath.registers.1226[17] [10])
);

DFFPOSX1 _21598_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf47),
    .D(_4663_),
    .Q(\datapath.registers.1226[17] [11])
);

DFFPOSX1 _21599_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf46),
    .D(_4664_),
    .Q(\datapath.registers.1226[17] [12])
);

DFFPOSX1 _21600_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf45),
    .D(_4665_),
    .Q(\datapath.registers.1226[17] [13])
);

DFFPOSX1 _21601_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf44),
    .D(_4666_),
    .Q(\datapath.registers.1226[17] [14])
);

DFFPOSX1 _21602_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf43),
    .D(_4667_),
    .Q(\datapath.registers.1226[17] [15])
);

DFFPOSX1 _21603_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf42),
    .D(_4668_),
    .Q(\datapath.registers.1226[17] [16])
);

DFFPOSX1 _21604_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf41),
    .D(_4669_),
    .Q(\datapath.registers.1226[17] [17])
);

DFFPOSX1 _21605_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf40),
    .D(_4670_),
    .Q(\datapath.registers.1226[17] [18])
);

DFFPOSX1 _21606_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf39),
    .D(_4671_),
    .Q(\datapath.registers.1226[17] [19])
);

DFFPOSX1 _21607_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf38),
    .D(_4673_),
    .Q(\datapath.registers.1226[17] [20])
);

DFFPOSX1 _21608_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf37),
    .D(_4674_),
    .Q(\datapath.registers.1226[17] [21])
);

DFFPOSX1 _21609_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf36),
    .D(_4675_),
    .Q(\datapath.registers.1226[17] [22])
);

DFFPOSX1 _21610_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf35),
    .D(_4676_),
    .Q(\datapath.registers.1226[17] [23])
);

DFFPOSX1 _21611_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf34),
    .D(_4677_),
    .Q(\datapath.registers.1226[17] [24])
);

DFFPOSX1 _21612_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf33),
    .D(_4678_),
    .Q(\datapath.registers.1226[17] [25])
);

DFFPOSX1 _21613_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf32),
    .D(_4679_),
    .Q(\datapath.registers.1226[17] [26])
);

DFFPOSX1 _21614_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf31),
    .D(_4680_),
    .Q(\datapath.registers.1226[17] [27])
);

DFFPOSX1 _21615_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf30),
    .D(_4681_),
    .Q(\datapath.registers.1226[17] [28])
);

DFFPOSX1 _21616_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf29),
    .D(_4682_),
    .Q(\datapath.registers.1226[17] [29])
);

DFFPOSX1 _21617_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf28),
    .D(_4684_),
    .Q(\datapath.registers.1226[17] [30])
);

DFFPOSX1 _21618_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf27),
    .D(_4685_),
    .Q(\datapath.registers.1226[17] [31])
);

DFFPOSX1 _21619_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf26),
    .D(_4469_),
    .Q(\datapath.registers.1226[11] [0])
);

DFFPOSX1 _21620_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf25),
    .D(_4480_),
    .Q(\datapath.registers.1226[11] [1])
);

DFFPOSX1 _21621_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf24),
    .D(_4491_),
    .Q(\datapath.registers.1226[11] [2])
);

DFFPOSX1 _21622_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf23),
    .D(_4494_),
    .Q(\datapath.registers.1226[11] [3])
);

DFFPOSX1 _21623_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf22),
    .D(_4495_),
    .Q(\datapath.registers.1226[11] [4])
);

DFFPOSX1 _21624_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf21),
    .D(_4496_),
    .Q(\datapath.registers.1226[11] [5])
);

DFFPOSX1 _21625_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf20),
    .D(_4497_),
    .Q(\datapath.registers.1226[11] [6])
);

DFFPOSX1 _21626_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf19),
    .D(_4498_),
    .Q(\datapath.registers.1226[11] [7])
);

DFFPOSX1 _21627_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf18),
    .D(_4499_),
    .Q(\datapath.registers.1226[11] [8])
);

DFFPOSX1 _21628_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf17),
    .D(_4500_),
    .Q(\datapath.registers.1226[11] [9])
);

DFFPOSX1 _21629_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf16),
    .D(_4470_),
    .Q(\datapath.registers.1226[11] [10])
);

DFFPOSX1 _21630_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf15),
    .D(_4471_),
    .Q(\datapath.registers.1226[11] [11])
);

DFFPOSX1 _21631_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf14),
    .D(_4472_),
    .Q(\datapath.registers.1226[11] [12])
);

DFFPOSX1 _21632_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf13),
    .D(_4473_),
    .Q(\datapath.registers.1226[11] [13])
);

DFFPOSX1 _21633_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf12),
    .D(_4474_),
    .Q(\datapath.registers.1226[11] [14])
);

DFFPOSX1 _21634_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf11),
    .D(_4475_),
    .Q(\datapath.registers.1226[11] [15])
);

DFFPOSX1 _21635_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf10),
    .D(_4476_),
    .Q(\datapath.registers.1226[11] [16])
);

DFFPOSX1 _21636_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf9),
    .D(_4477_),
    .Q(\datapath.registers.1226[11] [17])
);

DFFPOSX1 _21637_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf8),
    .D(_4478_),
    .Q(\datapath.registers.1226[11] [18])
);

DFFPOSX1 _21638_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf7),
    .D(_4479_),
    .Q(\datapath.registers.1226[11] [19])
);

DFFPOSX1 _21639_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf6),
    .D(_4481_),
    .Q(\datapath.registers.1226[11] [20])
);

DFFPOSX1 _21640_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf5),
    .D(_4482_),
    .Q(\datapath.registers.1226[11] [21])
);

DFFPOSX1 _21641_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf4),
    .D(_4483_),
    .Q(\datapath.registers.1226[11] [22])
);

DFFPOSX1 _21642_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf3),
    .D(_4484_),
    .Q(\datapath.registers.1226[11] [23])
);

DFFPOSX1 _21643_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf2),
    .D(_4485_),
    .Q(\datapath.registers.1226[11] [24])
);

DFFPOSX1 _21644_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf1),
    .D(_4486_),
    .Q(\datapath.registers.1226[11] [25])
);

DFFPOSX1 _21645_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf0),
    .D(_4487_),
    .Q(\datapath.registers.1226[11] [26])
);

DFFPOSX1 _21646_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf153),
    .D(_4488_),
    .Q(\datapath.registers.1226[11] [27])
);

DFFPOSX1 _21647_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf152),
    .D(_4489_),
    .Q(\datapath.registers.1226[11] [28])
);

DFFPOSX1 _21648_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf151),
    .D(_4490_),
    .Q(\datapath.registers.1226[11] [29])
);

DFFPOSX1 _21649_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf150),
    .D(_4492_),
    .Q(\datapath.registers.1226[11] [30])
);

DFFPOSX1 _21650_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf149),
    .D(_4493_),
    .Q(\datapath.registers.1226[11] [31])
);

DFFPOSX1 _21651_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf148),
    .D(_4565_),
    .Q(\datapath.registers.1226[14] [0])
);

DFFPOSX1 _21652_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf147),
    .D(_4576_),
    .Q(\datapath.registers.1226[14] [1])
);

DFFPOSX1 _21653_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf146),
    .D(_4587_),
    .Q(\datapath.registers.1226[14] [2])
);

DFFPOSX1 _21654_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf145),
    .D(_4590_),
    .Q(\datapath.registers.1226[14] [3])
);

DFFPOSX1 _21655_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf144),
    .D(_4591_),
    .Q(\datapath.registers.1226[14] [4])
);

DFFPOSX1 _21656_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf143),
    .D(_4592_),
    .Q(\datapath.registers.1226[14] [5])
);

DFFPOSX1 _21657_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf142),
    .D(_4593_),
    .Q(\datapath.registers.1226[14] [6])
);

DFFPOSX1 _21658_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf141),
    .D(_4594_),
    .Q(\datapath.registers.1226[14] [7])
);

DFFPOSX1 _21659_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf140),
    .D(_4595_),
    .Q(\datapath.registers.1226[14] [8])
);

DFFPOSX1 _21660_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf139),
    .D(_4596_),
    .Q(\datapath.registers.1226[14] [9])
);

DFFPOSX1 _21661_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf138),
    .D(_4566_),
    .Q(\datapath.registers.1226[14] [10])
);

DFFPOSX1 _21662_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf137),
    .D(_4567_),
    .Q(\datapath.registers.1226[14] [11])
);

DFFPOSX1 _21663_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf136),
    .D(_4568_),
    .Q(\datapath.registers.1226[14] [12])
);

DFFPOSX1 _21664_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf135),
    .D(_4569_),
    .Q(\datapath.registers.1226[14] [13])
);

DFFPOSX1 _21665_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf134),
    .D(_4570_),
    .Q(\datapath.registers.1226[14] [14])
);

DFFPOSX1 _21666_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf133),
    .D(_4571_),
    .Q(\datapath.registers.1226[14] [15])
);

DFFPOSX1 _21667_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf132),
    .D(_4572_),
    .Q(\datapath.registers.1226[14] [16])
);

DFFPOSX1 _21668_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf131),
    .D(_4573_),
    .Q(\datapath.registers.1226[14] [17])
);

DFFPOSX1 _21669_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf130),
    .D(_4574_),
    .Q(\datapath.registers.1226[14] [18])
);

DFFPOSX1 _21670_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf129),
    .D(_4575_),
    .Q(\datapath.registers.1226[14] [19])
);

DFFPOSX1 _21671_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf128),
    .D(_4577_),
    .Q(\datapath.registers.1226[14] [20])
);

DFFPOSX1 _21672_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf127),
    .D(_4578_),
    .Q(\datapath.registers.1226[14] [21])
);

DFFPOSX1 _21673_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf126),
    .D(_4579_),
    .Q(\datapath.registers.1226[14] [22])
);

DFFPOSX1 _21674_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf125),
    .D(_4580_),
    .Q(\datapath.registers.1226[14] [23])
);

DFFPOSX1 _21675_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf124),
    .D(_4581_),
    .Q(\datapath.registers.1226[14] [24])
);

DFFPOSX1 _21676_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf123),
    .D(_4582_),
    .Q(\datapath.registers.1226[14] [25])
);

DFFPOSX1 _21677_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf122),
    .D(_4583_),
    .Q(\datapath.registers.1226[14] [26])
);

DFFPOSX1 _21678_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf121),
    .D(_4584_),
    .Q(\datapath.registers.1226[14] [27])
);

DFFPOSX1 _21679_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf120),
    .D(_4585_),
    .Q(\datapath.registers.1226[14] [28])
);

DFFPOSX1 _21680_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf119),
    .D(_4586_),
    .Q(\datapath.registers.1226[14] [29])
);

DFFPOSX1 _21681_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf118),
    .D(_4588_),
    .Q(\datapath.registers.1226[14] [30])
);

DFFPOSX1 _21682_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf117),
    .D(_4589_),
    .Q(\datapath.registers.1226[14] [31])
);

DFFPOSX1 _21683_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf116),
    .D(_5333_),
    .Q(\datapath.registers.1226[7] [0])
);

DFFPOSX1 _21684_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf115),
    .D(_5344_),
    .Q(\datapath.registers.1226[7] [1])
);

DFFPOSX1 _21685_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf114),
    .D(_5355_),
    .Q(\datapath.registers.1226[7] [2])
);

DFFPOSX1 _21686_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf113),
    .D(_5358_),
    .Q(\datapath.registers.1226[7] [3])
);

DFFPOSX1 _21687_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf112),
    .D(_5359_),
    .Q(\datapath.registers.1226[7] [4])
);

DFFPOSX1 _21688_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf111),
    .D(_5360_),
    .Q(\datapath.registers.1226[7] [5])
);

DFFPOSX1 _21689_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf110),
    .D(_5361_),
    .Q(\datapath.registers.1226[7] [6])
);

DFFPOSX1 _21690_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf109),
    .D(_5362_),
    .Q(\datapath.registers.1226[7] [7])
);

DFFPOSX1 _21691_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf108),
    .D(_5363_),
    .Q(\datapath.registers.1226[7] [8])
);

DFFPOSX1 _21692_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf107),
    .D(_5364_),
    .Q(\datapath.registers.1226[7] [9])
);

DFFPOSX1 _21693_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf106),
    .D(_5334_),
    .Q(\datapath.registers.1226[7] [10])
);

DFFPOSX1 _21694_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf105),
    .D(_5335_),
    .Q(\datapath.registers.1226[7] [11])
);

DFFPOSX1 _21695_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf104),
    .D(_5336_),
    .Q(\datapath.registers.1226[7] [12])
);

DFFPOSX1 _21696_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf103),
    .D(_5337_),
    .Q(\datapath.registers.1226[7] [13])
);

DFFPOSX1 _21697_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf102),
    .D(_5338_),
    .Q(\datapath.registers.1226[7] [14])
);

DFFPOSX1 _21698_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf101),
    .D(_5339_),
    .Q(\datapath.registers.1226[7] [15])
);

DFFPOSX1 _21699_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf100),
    .D(_5340_),
    .Q(\datapath.registers.1226[7] [16])
);

DFFPOSX1 _21700_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf99),
    .D(_5341_),
    .Q(\datapath.registers.1226[7] [17])
);

DFFPOSX1 _21701_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf98),
    .D(_5342_),
    .Q(\datapath.registers.1226[7] [18])
);

DFFPOSX1 _21702_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf97),
    .D(_5343_),
    .Q(\datapath.registers.1226[7] [19])
);

DFFPOSX1 _21703_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf96),
    .D(_5345_),
    .Q(\datapath.registers.1226[7] [20])
);

DFFPOSX1 _21704_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf95),
    .D(_5346_),
    .Q(\datapath.registers.1226[7] [21])
);

DFFPOSX1 _21705_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf94),
    .D(_5347_),
    .Q(\datapath.registers.1226[7] [22])
);

DFFPOSX1 _21706_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf93),
    .D(_5348_),
    .Q(\datapath.registers.1226[7] [23])
);

DFFPOSX1 _21707_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf92),
    .D(_5349_),
    .Q(\datapath.registers.1226[7] [24])
);

DFFPOSX1 _21708_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf91),
    .D(_5350_),
    .Q(\datapath.registers.1226[7] [25])
);

DFFPOSX1 _21709_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf90),
    .D(_5351_),
    .Q(\datapath.registers.1226[7] [26])
);

DFFPOSX1 _21710_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf89),
    .D(_5352_),
    .Q(\datapath.registers.1226[7] [27])
);

DFFPOSX1 _21711_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf88),
    .D(_5353_),
    .Q(\datapath.registers.1226[7] [28])
);

DFFPOSX1 _21712_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf87),
    .D(_5354_),
    .Q(\datapath.registers.1226[7] [29])
);

DFFPOSX1 _21713_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf86),
    .D(_5356_),
    .Q(\datapath.registers.1226[7] [30])
);

DFFPOSX1 _21714_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf85),
    .D(_5357_),
    .Q(\datapath.registers.1226[7] [31])
);

DFFPOSX1 _21715_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf84),
    .D(_5141_),
    .Q(\datapath.registers.1226[30] [0])
);

DFFPOSX1 _21716_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf83),
    .D(_5152_),
    .Q(\datapath.registers.1226[30] [1])
);

DFFPOSX1 _21717_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf82),
    .D(_5163_),
    .Q(\datapath.registers.1226[30] [2])
);

DFFPOSX1 _21718_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf81),
    .D(_5166_),
    .Q(\datapath.registers.1226[30] [3])
);

DFFPOSX1 _21719_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf80),
    .D(_5167_),
    .Q(\datapath.registers.1226[30] [4])
);

DFFPOSX1 _21720_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf79),
    .D(_5168_),
    .Q(\datapath.registers.1226[30] [5])
);

DFFPOSX1 _21721_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf78),
    .D(_5169_),
    .Q(\datapath.registers.1226[30] [6])
);

DFFPOSX1 _21722_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf77),
    .D(_5170_),
    .Q(\datapath.registers.1226[30] [7])
);

DFFPOSX1 _21723_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf76),
    .D(_5171_),
    .Q(\datapath.registers.1226[30] [8])
);

DFFPOSX1 _21724_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf75),
    .D(_5172_),
    .Q(\datapath.registers.1226[30] [9])
);

DFFPOSX1 _21725_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf74),
    .D(_5142_),
    .Q(\datapath.registers.1226[30] [10])
);

DFFPOSX1 _21726_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf73),
    .D(_5143_),
    .Q(\datapath.registers.1226[30] [11])
);

DFFPOSX1 _21727_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf72),
    .D(_5144_),
    .Q(\datapath.registers.1226[30] [12])
);

DFFPOSX1 _21728_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf71),
    .D(_5145_),
    .Q(\datapath.registers.1226[30] [13])
);

DFFPOSX1 _21729_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf70),
    .D(_5146_),
    .Q(\datapath.registers.1226[30] [14])
);

DFFPOSX1 _21730_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf69),
    .D(_5147_),
    .Q(\datapath.registers.1226[30] [15])
);

DFFPOSX1 _21731_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf68),
    .D(_5148_),
    .Q(\datapath.registers.1226[30] [16])
);

DFFPOSX1 _21732_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf67),
    .D(_5149_),
    .Q(\datapath.registers.1226[30] [17])
);

DFFPOSX1 _21733_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf66),
    .D(_5150_),
    .Q(\datapath.registers.1226[30] [18])
);

DFFPOSX1 _21734_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf65),
    .D(_5151_),
    .Q(\datapath.registers.1226[30] [19])
);

DFFPOSX1 _21735_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf64),
    .D(_5153_),
    .Q(\datapath.registers.1226[30] [20])
);

DFFPOSX1 _21736_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf63),
    .D(_5154_),
    .Q(\datapath.registers.1226[30] [21])
);

DFFPOSX1 _21737_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf62),
    .D(_5155_),
    .Q(\datapath.registers.1226[30] [22])
);

DFFPOSX1 _21738_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf61),
    .D(_5156_),
    .Q(\datapath.registers.1226[30] [23])
);

DFFPOSX1 _21739_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf60),
    .D(_5157_),
    .Q(\datapath.registers.1226[30] [24])
);

DFFPOSX1 _21740_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf59),
    .D(_5158_),
    .Q(\datapath.registers.1226[30] [25])
);

DFFPOSX1 _21741_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf58),
    .D(_5159_),
    .Q(\datapath.registers.1226[30] [26])
);

DFFPOSX1 _21742_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf57),
    .D(_5160_),
    .Q(\datapath.registers.1226[30] [27])
);

DFFPOSX1 _21743_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf56),
    .D(_5161_),
    .Q(\datapath.registers.1226[30] [28])
);

DFFPOSX1 _21744_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf55),
    .D(_5162_),
    .Q(\datapath.registers.1226[30] [29])
);

DFFPOSX1 _21745_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf54),
    .D(_5164_),
    .Q(\datapath.registers.1226[30] [30])
);

DFFPOSX1 _21746_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf53),
    .D(_5165_),
    .Q(\datapath.registers.1226[30] [31])
);

DFFPOSX1 _21747_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf52),
    .D(_5077_),
    .Q(\datapath.registers.1226[29] [0])
);

DFFPOSX1 _21748_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf51),
    .D(_5088_),
    .Q(\datapath.registers.1226[29] [1])
);

DFFPOSX1 _21749_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf50),
    .D(_5099_),
    .Q(\datapath.registers.1226[29] [2])
);

DFFPOSX1 _21750_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf49),
    .D(_5102_),
    .Q(\datapath.registers.1226[29] [3])
);

DFFPOSX1 _21751_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf48),
    .D(_5103_),
    .Q(\datapath.registers.1226[29] [4])
);

DFFPOSX1 _21752_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf47),
    .D(_5104_),
    .Q(\datapath.registers.1226[29] [5])
);

DFFPOSX1 _21753_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf46),
    .D(_5105_),
    .Q(\datapath.registers.1226[29] [6])
);

DFFPOSX1 _21754_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf45),
    .D(_5106_),
    .Q(\datapath.registers.1226[29] [7])
);

DFFPOSX1 _21755_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf44),
    .D(_5107_),
    .Q(\datapath.registers.1226[29] [8])
);

DFFPOSX1 _21756_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf43),
    .D(_5108_),
    .Q(\datapath.registers.1226[29] [9])
);

DFFPOSX1 _21757_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf42),
    .D(_5078_),
    .Q(\datapath.registers.1226[29] [10])
);

DFFPOSX1 _21758_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf41),
    .D(_5079_),
    .Q(\datapath.registers.1226[29] [11])
);

DFFPOSX1 _21759_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf40),
    .D(_5080_),
    .Q(\datapath.registers.1226[29] [12])
);

DFFPOSX1 _21760_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf39),
    .D(_5081_),
    .Q(\datapath.registers.1226[29] [13])
);

DFFPOSX1 _21761_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf38),
    .D(_5082_),
    .Q(\datapath.registers.1226[29] [14])
);

DFFPOSX1 _21762_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf37),
    .D(_5083_),
    .Q(\datapath.registers.1226[29] [15])
);

DFFPOSX1 _21763_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf36),
    .D(_5084_),
    .Q(\datapath.registers.1226[29] [16])
);

DFFPOSX1 _21764_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf35),
    .D(_5085_),
    .Q(\datapath.registers.1226[29] [17])
);

DFFPOSX1 _21765_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf34),
    .D(_5086_),
    .Q(\datapath.registers.1226[29] [18])
);

DFFPOSX1 _21766_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf33),
    .D(_5087_),
    .Q(\datapath.registers.1226[29] [19])
);

DFFPOSX1 _21767_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf32),
    .D(_5089_),
    .Q(\datapath.registers.1226[29] [20])
);

DFFPOSX1 _21768_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf31),
    .D(_5090_),
    .Q(\datapath.registers.1226[29] [21])
);

DFFPOSX1 _21769_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf30),
    .D(_5091_),
    .Q(\datapath.registers.1226[29] [22])
);

DFFPOSX1 _21770_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf29),
    .D(_5092_),
    .Q(\datapath.registers.1226[29] [23])
);

DFFPOSX1 _21771_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf28),
    .D(_5093_),
    .Q(\datapath.registers.1226[29] [24])
);

DFFPOSX1 _21772_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf27),
    .D(_5094_),
    .Q(\datapath.registers.1226[29] [25])
);

DFFPOSX1 _21773_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf26),
    .D(_5095_),
    .Q(\datapath.registers.1226[29] [26])
);

DFFPOSX1 _21774_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf25),
    .D(_5096_),
    .Q(\datapath.registers.1226[29] [27])
);

DFFPOSX1 _21775_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf24),
    .D(_5097_),
    .Q(\datapath.registers.1226[29] [28])
);

DFFPOSX1 _21776_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf23),
    .D(_5098_),
    .Q(\datapath.registers.1226[29] [29])
);

DFFPOSX1 _21777_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf22),
    .D(_5100_),
    .Q(\datapath.registers.1226[29] [30])
);

DFFPOSX1 _21778_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf21),
    .D(_5101_),
    .Q(\datapath.registers.1226[29] [31])
);

DFFPOSX1 _21779_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf20),
    .D(_5301_),
    .Q(\datapath.registers.1226[6] [0])
);

DFFPOSX1 _21780_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf19),
    .D(_5312_),
    .Q(\datapath.registers.1226[6] [1])
);

DFFPOSX1 _21781_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf18),
    .D(_5323_),
    .Q(\datapath.registers.1226[6] [2])
);

DFFPOSX1 _21782_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf17),
    .D(_5326_),
    .Q(\datapath.registers.1226[6] [3])
);

DFFPOSX1 _21783_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf16),
    .D(_5327_),
    .Q(\datapath.registers.1226[6] [4])
);

DFFPOSX1 _21784_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf15),
    .D(_5328_),
    .Q(\datapath.registers.1226[6] [5])
);

DFFPOSX1 _21785_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf14),
    .D(_5329_),
    .Q(\datapath.registers.1226[6] [6])
);

DFFPOSX1 _21786_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf13),
    .D(_5330_),
    .Q(\datapath.registers.1226[6] [7])
);

DFFPOSX1 _21787_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf12),
    .D(_5331_),
    .Q(\datapath.registers.1226[6] [8])
);

DFFPOSX1 _21788_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf11),
    .D(_5332_),
    .Q(\datapath.registers.1226[6] [9])
);

DFFPOSX1 _21789_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf10),
    .D(_5302_),
    .Q(\datapath.registers.1226[6] [10])
);

DFFPOSX1 _21790_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf9),
    .D(_5303_),
    .Q(\datapath.registers.1226[6] [11])
);

DFFPOSX1 _21791_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf8),
    .D(_5304_),
    .Q(\datapath.registers.1226[6] [12])
);

DFFPOSX1 _21792_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf7),
    .D(_5305_),
    .Q(\datapath.registers.1226[6] [13])
);

DFFPOSX1 _21793_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf6),
    .D(_5306_),
    .Q(\datapath.registers.1226[6] [14])
);

DFFPOSX1 _21794_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf5),
    .D(_5307_),
    .Q(\datapath.registers.1226[6] [15])
);

DFFPOSX1 _21795_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf4),
    .D(_5308_),
    .Q(\datapath.registers.1226[6] [16])
);

DFFPOSX1 _21796_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf3),
    .D(_5309_),
    .Q(\datapath.registers.1226[6] [17])
);

DFFPOSX1 _21797_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf2),
    .D(_5310_),
    .Q(\datapath.registers.1226[6] [18])
);

DFFPOSX1 _21798_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf1),
    .D(_5311_),
    .Q(\datapath.registers.1226[6] [19])
);

DFFPOSX1 _21799_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf0),
    .D(_5313_),
    .Q(\datapath.registers.1226[6] [20])
);

DFFPOSX1 _21800_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf153),
    .D(_5314_),
    .Q(\datapath.registers.1226[6] [21])
);

DFFPOSX1 _21801_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf152),
    .D(_5315_),
    .Q(\datapath.registers.1226[6] [22])
);

DFFPOSX1 _21802_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf151),
    .D(_5316_),
    .Q(\datapath.registers.1226[6] [23])
);

DFFPOSX1 _21803_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf150),
    .D(_5317_),
    .Q(\datapath.registers.1226[6] [24])
);

DFFPOSX1 _21804_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf149),
    .D(_5318_),
    .Q(\datapath.registers.1226[6] [25])
);

DFFPOSX1 _21805_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf148),
    .D(_5319_),
    .Q(\datapath.registers.1226[6] [26])
);

DFFPOSX1 _21806_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf147),
    .D(_5320_),
    .Q(\datapath.registers.1226[6] [27])
);

DFFPOSX1 _21807_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf146),
    .D(_5321_),
    .Q(\datapath.registers.1226[6] [28])
);

DFFPOSX1 _21808_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf145),
    .D(_5322_),
    .Q(\datapath.registers.1226[6] [29])
);

DFFPOSX1 _21809_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf144),
    .D(_5324_),
    .Q(\datapath.registers.1226[6] [30])
);

DFFPOSX1 _21810_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf143),
    .D(_5325_),
    .Q(\datapath.registers.1226[6] [31])
);

DFFPOSX1 _21811_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf142),
    .D(_4949_),
    .Q(\datapath.registers.1226[25] [0])
);

DFFPOSX1 _21812_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf141),
    .D(_4960_),
    .Q(\datapath.registers.1226[25] [1])
);

DFFPOSX1 _21813_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf140),
    .D(_4971_),
    .Q(\datapath.registers.1226[25] [2])
);

DFFPOSX1 _21814_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf139),
    .D(_4974_),
    .Q(\datapath.registers.1226[25] [3])
);

DFFPOSX1 _21815_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf138),
    .D(_4975_),
    .Q(\datapath.registers.1226[25] [4])
);

DFFPOSX1 _21816_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf137),
    .D(_4976_),
    .Q(\datapath.registers.1226[25] [5])
);

DFFPOSX1 _21817_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf136),
    .D(_4977_),
    .Q(\datapath.registers.1226[25] [6])
);

DFFPOSX1 _21818_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf135),
    .D(_4978_),
    .Q(\datapath.registers.1226[25] [7])
);

DFFPOSX1 _21819_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf134),
    .D(_4979_),
    .Q(\datapath.registers.1226[25] [8])
);

DFFPOSX1 _21820_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf133),
    .D(_4980_),
    .Q(\datapath.registers.1226[25] [9])
);

DFFPOSX1 _21821_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf132),
    .D(_4950_),
    .Q(\datapath.registers.1226[25] [10])
);

DFFPOSX1 _21822_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf131),
    .D(_4951_),
    .Q(\datapath.registers.1226[25] [11])
);

DFFPOSX1 _21823_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf130),
    .D(_4952_),
    .Q(\datapath.registers.1226[25] [12])
);

DFFPOSX1 _21824_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf129),
    .D(_4953_),
    .Q(\datapath.registers.1226[25] [13])
);

DFFPOSX1 _21825_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf128),
    .D(_4954_),
    .Q(\datapath.registers.1226[25] [14])
);

DFFPOSX1 _21826_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf127),
    .D(_4955_),
    .Q(\datapath.registers.1226[25] [15])
);

DFFPOSX1 _21827_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf126),
    .D(_4956_),
    .Q(\datapath.registers.1226[25] [16])
);

DFFPOSX1 _21828_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf125),
    .D(_4957_),
    .Q(\datapath.registers.1226[25] [17])
);

DFFPOSX1 _21829_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf124),
    .D(_4958_),
    .Q(\datapath.registers.1226[25] [18])
);

DFFPOSX1 _21830_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf123),
    .D(_4959_),
    .Q(\datapath.registers.1226[25] [19])
);

DFFPOSX1 _21831_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf122),
    .D(_4961_),
    .Q(\datapath.registers.1226[25] [20])
);

DFFPOSX1 _21832_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf121),
    .D(_4962_),
    .Q(\datapath.registers.1226[25] [21])
);

DFFPOSX1 _21833_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf120),
    .D(_4963_),
    .Q(\datapath.registers.1226[25] [22])
);

DFFPOSX1 _21834_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf119),
    .D(_4964_),
    .Q(\datapath.registers.1226[25] [23])
);

DFFPOSX1 _21835_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf118),
    .D(_4965_),
    .Q(\datapath.registers.1226[25] [24])
);

DFFPOSX1 _21836_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf117),
    .D(_4966_),
    .Q(\datapath.registers.1226[25] [25])
);

DFFPOSX1 _21837_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf116),
    .D(_4967_),
    .Q(\datapath.registers.1226[25] [26])
);

DFFPOSX1 _21838_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf115),
    .D(_4968_),
    .Q(\datapath.registers.1226[25] [27])
);

DFFPOSX1 _21839_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf114),
    .D(_4969_),
    .Q(\datapath.registers.1226[25] [28])
);

DFFPOSX1 _21840_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf113),
    .D(_4970_),
    .Q(\datapath.registers.1226[25] [29])
);

DFFPOSX1 _21841_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf112),
    .D(_4972_),
    .Q(\datapath.registers.1226[25] [30])
);

DFFPOSX1 _21842_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf111),
    .D(_4973_),
    .Q(\datapath.registers.1226[25] [31])
);

DFFPOSX1 _21843_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf110),
    .D(_5045_),
    .Q(\datapath.registers.1226[28] [0])
);

DFFPOSX1 _21844_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf109),
    .D(_5056_),
    .Q(\datapath.registers.1226[28] [1])
);

DFFPOSX1 _21845_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf108),
    .D(_5067_),
    .Q(\datapath.registers.1226[28] [2])
);

DFFPOSX1 _21846_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf107),
    .D(_5070_),
    .Q(\datapath.registers.1226[28] [3])
);

DFFPOSX1 _21847_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf106),
    .D(_5071_),
    .Q(\datapath.registers.1226[28] [4])
);

DFFPOSX1 _21848_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf105),
    .D(_5072_),
    .Q(\datapath.registers.1226[28] [5])
);

DFFPOSX1 _21849_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf104),
    .D(_5073_),
    .Q(\datapath.registers.1226[28] [6])
);

DFFPOSX1 _21850_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf103),
    .D(_5074_),
    .Q(\datapath.registers.1226[28] [7])
);

DFFPOSX1 _21851_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf102),
    .D(_5075_),
    .Q(\datapath.registers.1226[28] [8])
);

DFFPOSX1 _21852_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf101),
    .D(_5076_),
    .Q(\datapath.registers.1226[28] [9])
);

DFFPOSX1 _21853_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf100),
    .D(_5046_),
    .Q(\datapath.registers.1226[28] [10])
);

DFFPOSX1 _21854_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf99),
    .D(_5047_),
    .Q(\datapath.registers.1226[28] [11])
);

DFFPOSX1 _21855_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf98),
    .D(_5048_),
    .Q(\datapath.registers.1226[28] [12])
);

DFFPOSX1 _21856_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf97),
    .D(_5049_),
    .Q(\datapath.registers.1226[28] [13])
);

DFFPOSX1 _21857_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf96),
    .D(_5050_),
    .Q(\datapath.registers.1226[28] [14])
);

DFFPOSX1 _21858_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf95),
    .D(_5051_),
    .Q(\datapath.registers.1226[28] [15])
);

DFFPOSX1 _21859_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf94),
    .D(_5052_),
    .Q(\datapath.registers.1226[28] [16])
);

DFFPOSX1 _21860_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf93),
    .D(_5053_),
    .Q(\datapath.registers.1226[28] [17])
);

DFFPOSX1 _21861_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf92),
    .D(_5054_),
    .Q(\datapath.registers.1226[28] [18])
);

DFFPOSX1 _21862_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf91),
    .D(_5055_),
    .Q(\datapath.registers.1226[28] [19])
);

DFFPOSX1 _21863_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf90),
    .D(_5057_),
    .Q(\datapath.registers.1226[28] [20])
);

DFFPOSX1 _21864_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf89),
    .D(_5058_),
    .Q(\datapath.registers.1226[28] [21])
);

DFFPOSX1 _21865_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf88),
    .D(_5059_),
    .Q(\datapath.registers.1226[28] [22])
);

DFFPOSX1 _21866_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf87),
    .D(_5060_),
    .Q(\datapath.registers.1226[28] [23])
);

DFFPOSX1 _21867_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf86),
    .D(_5061_),
    .Q(\datapath.registers.1226[28] [24])
);

DFFPOSX1 _21868_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf85),
    .D(_5062_),
    .Q(\datapath.registers.1226[28] [25])
);

DFFPOSX1 _21869_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf84),
    .D(_5063_),
    .Q(\datapath.registers.1226[28] [26])
);

DFFPOSX1 _21870_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf83),
    .D(_5064_),
    .Q(\datapath.registers.1226[28] [27])
);

DFFPOSX1 _21871_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf82),
    .D(_5065_),
    .Q(\datapath.registers.1226[28] [28])
);

DFFPOSX1 _21872_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf81),
    .D(_5066_),
    .Q(\datapath.registers.1226[28] [29])
);

DFFPOSX1 _21873_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf80),
    .D(_5068_),
    .Q(\datapath.registers.1226[28] [30])
);

DFFPOSX1 _21874_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(CLK_bF$buf79),
    .D(_5069_),
    .Q(\datapath.registers.1226[28] [31])
);

BUFX2 _9443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__0_bF$buf4),
    .Y(DMEM_ADDR[0])
);

BUFX2 _9444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf5),
    .Y(DMEM_ADDR[1])
);

BUFX2 _9445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[2]),
    .Y(DMEM_ADDR[2])
);

BUFX2 _9446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[3]),
    .Y(DMEM_ADDR[3])
);

BUFX2 _9447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[4]),
    .Y(DMEM_ADDR[4])
);

BUFX2 _9448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[5]),
    .Y(DMEM_ADDR[5])
);

BUFX2 _9449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[6]),
    .Y(DMEM_ADDR[6])
);

BUFX2 _9450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[7]),
    .Y(DMEM_ADDR[7])
);

BUFX2 _9451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[8]),
    .Y(DMEM_ADDR[8])
);

BUFX2 _9452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[9]),
    .Y(DMEM_ADDR[9])
);

BUFX2 _9453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[10]),
    .Y(DMEM_ADDR[10])
);

BUFX2 _9454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[11]),
    .Y(DMEM_ADDR[11])
);

BUFX2 _9455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[12]),
    .Y(DMEM_ADDR[12])
);

BUFX2 _9456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[13]),
    .Y(DMEM_ADDR[13])
);

BUFX2 _9457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[14]),
    .Y(DMEM_ADDR[14])
);

BUFX2 _9458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[15]),
    .Y(DMEM_ADDR[15])
);

BUFX2 _9459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[16]),
    .Y(DMEM_ADDR[16])
);

BUFX2 _9460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[17]),
    .Y(DMEM_ADDR[17])
);

BUFX2 _9461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[18]),
    .Y(DMEM_ADDR[18])
);

BUFX2 _9462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[19]),
    .Y(DMEM_ADDR[19])
);

BUFX2 _9463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[20]),
    .Y(DMEM_ADDR[20])
);

BUFX2 _9464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[21]),
    .Y(DMEM_ADDR[21])
);

BUFX2 _9465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[22]),
    .Y(DMEM_ADDR[22])
);

BUFX2 _9466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[23]),
    .Y(DMEM_ADDR[23])
);

BUFX2 _9467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[24]),
    .Y(DMEM_ADDR[24])
);

BUFX2 _9468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[25]),
    .Y(DMEM_ADDR[25])
);

BUFX2 _9469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[26]),
    .Y(DMEM_ADDR[26])
);

BUFX2 _9470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[27]),
    .Y(DMEM_ADDR[27])
);

BUFX2 _9471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[28]),
    .Y(DMEM_ADDR[28])
);

BUFX2 _9472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[29]),
    .Y(DMEM_ADDR[29])
);

BUFX2 _9473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[30]),
    .Y(DMEM_ADDR[30])
);

BUFX2 _9474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[31]),
    .Y(DMEM_ADDR[31])
);

BUFX2 _9475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[0]),
    .Y(DMEM_DATA_S[0])
);

BUFX2 _9476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[1]),
    .Y(DMEM_DATA_S[1])
);

BUFX2 _9477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[2]),
    .Y(DMEM_DATA_S[2])
);

BUFX2 _9478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[3]),
    .Y(DMEM_DATA_S[3])
);

BUFX2 _9479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[4]),
    .Y(DMEM_DATA_S[4])
);

BUFX2 _9480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[5]),
    .Y(DMEM_DATA_S[5])
);

BUFX2 _9481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[6]),
    .Y(DMEM_DATA_S[6])
);

BUFX2 _9482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[7]),
    .Y(DMEM_DATA_S[7])
);

BUFX2 _9483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[8]),
    .Y(DMEM_DATA_S[8])
);

BUFX2 _9484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[9]),
    .Y(DMEM_DATA_S[9])
);

BUFX2 _9485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[10]),
    .Y(DMEM_DATA_S[10])
);

BUFX2 _9486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[11]),
    .Y(DMEM_DATA_S[11])
);

BUFX2 _9487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[12]),
    .Y(DMEM_DATA_S[12])
);

BUFX2 _9488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[13]),
    .Y(DMEM_DATA_S[13])
);

BUFX2 _9489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[14]),
    .Y(DMEM_DATA_S[14])
);

BUFX2 _9490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[15]),
    .Y(DMEM_DATA_S[15])
);

BUFX2 _9491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[16]),
    .Y(DMEM_DATA_S[16])
);

BUFX2 _9492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[17]),
    .Y(DMEM_DATA_S[17])
);

BUFX2 _9493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[18]),
    .Y(DMEM_DATA_S[18])
);

BUFX2 _9494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[19]),
    .Y(DMEM_DATA_S[19])
);

BUFX2 _9495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[20]),
    .Y(DMEM_DATA_S[20])
);

BUFX2 _9496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[21]),
    .Y(DMEM_DATA_S[21])
);

BUFX2 _9497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[22]),
    .Y(DMEM_DATA_S[22])
);

BUFX2 _9498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[23]),
    .Y(DMEM_DATA_S[23])
);

BUFX2 _9499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[24]),
    .Y(DMEM_DATA_S[24])
);

BUFX2 _9500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[25]),
    .Y(DMEM_DATA_S[25])
);

BUFX2 _9501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[26]),
    .Y(DMEM_DATA_S[26])
);

BUFX2 _9502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[27]),
    .Y(DMEM_DATA_S[27])
);

BUFX2 _9503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[28]),
    .Y(DMEM_DATA_S[28])
);

BUFX2 _9504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[29]),
    .Y(DMEM_DATA_S[29])
);

BUFX2 _9505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[30]),
    .Y(DMEM_DATA_S[30])
);

BUFX2 _9506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1_[31]),
    .Y(DMEM_DATA_S[31])
);

BUFX2 _9507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_),
    .Y(DMEM_WEN)
);

BUFX2 _9508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [0]),
    .Y(IMEM_ADDR[0])
);

BUFX2 _9509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [1]),
    .Y(IMEM_ADDR[1])
);

BUFX2 _9510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [2]),
    .Y(IMEM_ADDR[2])
);

BUFX2 _9511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [3]),
    .Y(IMEM_ADDR[3])
);

BUFX2 _9512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [4]),
    .Y(IMEM_ADDR[4])
);

BUFX2 _9513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [5]),
    .Y(IMEM_ADDR[5])
);

BUFX2 _9514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [6]),
    .Y(IMEM_ADDR[6])
);

BUFX2 _9515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [7]),
    .Y(IMEM_ADDR[7])
);

BUFX2 _9516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [8]),
    .Y(IMEM_ADDR[8])
);

BUFX2 _9517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [9]),
    .Y(IMEM_ADDR[9])
);

BUFX2 _9518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [10]),
    .Y(IMEM_ADDR[10])
);

BUFX2 _9519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [11]),
    .Y(IMEM_ADDR[11])
);

BUFX2 _9520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [12]),
    .Y(IMEM_ADDR[12])
);

BUFX2 _9521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [13]),
    .Y(IMEM_ADDR[13])
);

BUFX2 _9522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [14]),
    .Y(IMEM_ADDR[14])
);

BUFX2 _9523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [15]),
    .Y(IMEM_ADDR[15])
);

BUFX2 _9524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [16]),
    .Y(IMEM_ADDR[16])
);

BUFX2 _9525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [17]),
    .Y(IMEM_ADDR[17])
);

BUFX2 _9526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [18]),
    .Y(IMEM_ADDR[18])
);

BUFX2 _9527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [19]),
    .Y(IMEM_ADDR[19])
);

BUFX2 _9528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [20]),
    .Y(IMEM_ADDR[20])
);

BUFX2 _9529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [21]),
    .Y(IMEM_ADDR[21])
);

BUFX2 _9530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [22]),
    .Y(IMEM_ADDR[22])
);

BUFX2 _9531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [23]),
    .Y(IMEM_ADDR[23])
);

BUFX2 _9532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [24]),
    .Y(IMEM_ADDR[24])
);

BUFX2 _9533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [25]),
    .Y(IMEM_ADDR[25])
);

BUFX2 _9534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [26]),
    .Y(IMEM_ADDR[26])
);

BUFX2 _9535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [27]),
    .Y(IMEM_ADDR[27])
);

BUFX2 _9536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [28]),
    .Y(IMEM_ADDR[28])
);

BUFX2 _9537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [29]),
    .Y(IMEM_ADDR[29])
);

BUFX2 _9538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [30]),
    .Y(IMEM_ADDR[30])
);

BUFX2 _9539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [31]),
    .Y(IMEM_ADDR[31])
);

NOR2X1 _9540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [4]),
    .B(\datapath.meminstr [6]),
    .Y(_104_)
);

NOR2X1 _9541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [3]),
    .B(\datapath.meminstr [2]),
    .Y(_105_)
);

INVX2 _9542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_105_),
    .Y(_106_)
);

NOR2X1 _9543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [5]),
    .B(_106_),
    .Y(_107_)
);

AND2X2 _9544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_107_),
    .B(_104_),
    .Y(_108_)
);

XOR2X1 _9545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_19_bF$buf5 ),
    .B(\datapath.meminstr [11]),
    .Y(_109_)
);

INVX2 _9546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [8]),
    .Y(_110_)
);

INVX2 _9547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [10]),
    .Y(_111_)
);

OAI22X1 _9548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_110_),
    .B(\datapath.idinstr_16_bF$buf13 ),
    .C(\datapath.idinstr_18_bF$buf3 ),
    .D(_111_),
    .Y(_112_)
);

NOR2X1 _9549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112_),
    .B(_109_),
    .Y(_113_)
);

INVX1 _9550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [9]),
    .Y(_114_)
);

AOI22X1 _9551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114_),
    .B(\datapath.idinstr_17_bF$buf23 ),
    .C(\datapath.idinstr_18_bF$buf2 ),
    .D(_111_),
    .Y(_115_)
);

INVX1 _9552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf22 ),
    .Y(_116_)
);

AOI22X1 _9553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_116_),
    .B(\datapath.meminstr [9]),
    .C(\datapath.idinstr_16_bF$buf12 ),
    .D(_110_),
    .Y(_117_)
);

AND2X2 _9554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_115_),
    .B(_117_),
    .Y(_118_)
);

INVX1 _9555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [4]),
    .Y(_119_)
);

NAND2X1 _9556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [5]),
    .B(_119_),
    .Y(_120_)
);

NOR2X1 _9557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_120_),
    .B(_106_),
    .Y(_121_)
);

XOR2X1 _9558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf29 ),
    .B(\datapath.meminstr [7]),
    .Y(_122_)
);

NOR2X1 _9559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_122_),
    .B(_121_),
    .Y(_123_)
);

NAND3X1 _9560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_113_),
    .B(_118_),
    .C(_123_),
    .Y(_124_)
);

OR2X2 _9561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_124_),
    .B(_108_),
    .Y(_125_)
);

XNOR2X1 _9562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [10]),
    .B(\datapath.idinstr_18_bF$buf1 ),
    .Y(_126_)
);

XNOR2X1 _9563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [11]),
    .B(\datapath.idinstr_19_bF$buf4 ),
    .Y(_127_)
);

XNOR2X1 _9564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [7]),
    .B(\datapath.idinstr_15_bF$buf28 ),
    .Y(_128_)
);

NAND3X1 _9565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_126_),
    .B(_127_),
    .C(_128_),
    .Y(_129_)
);

INVX1 _9566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [4]),
    .Y(_130_)
);

NOR2X1 _9567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [3]),
    .B(\datapath.wbinstr [2]),
    .Y(_131_)
);

NAND3X1 _9568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_130_),
    .B(\datapath.wbinstr [5]),
    .C(_131_),
    .Y(_132_)
);

XNOR2X1 _9569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [9]),
    .B(\datapath.idinstr_17_bF$buf21 ),
    .Y(_133_)
);

XNOR2X1 _9570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [8]),
    .B(\datapath.idinstr_16_bF$buf11 ),
    .Y(_134_)
);

NAND3X1 _9571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_133_),
    .B(_134_),
    .C(_132_),
    .Y(_135_)
);

NOR2X1 _9572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_135_),
    .Y(_136_)
);

NAND2X1 _9573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_136_),
    .B(_124_),
    .Y(_137_)
);

INVX2 _9574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [6]),
    .Y(_138_)
);

INVX2 _9575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [3]),
    .Y(_3_)
);

NOR2X1 _9576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [4]),
    .B(_3_),
    .Y(_4_)
);

AOI21X1 _9577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [5]),
    .B(_4_),
    .C(_138_),
    .Y(_5_)
);

INVX1 _9578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [2]),
    .Y(_6_)
);

AOI21X1 _9579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [4]),
    .B(_3_),
    .C(\datapath.idinstr [6]),
    .Y(_7_)
);

OR2X2 _9580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7_),
    .B(_6_),
    .Y(_8_)
);

NOR2X1 _9581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf27 ),
    .B(\datapath.idinstr_16_bF$buf10 ),
    .Y(_9_)
);

OR2X2 _9582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf20 ),
    .B(\datapath.idinstr_18_bF$buf0 ),
    .Y(_10_)
);

NOR2X1 _9583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_19_bF$buf3 ),
    .B(_10_),
    .Y(_11_)
);

NAND2X1 _9584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9_),
    .B(_11_),
    .Y(_12_)
);

OAI21X1 _9585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8_),
    .B(_5_),
    .C(_12_),
    .Y(_13_)
);

XOR2X1 _9586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_16_bF$buf9 ),
    .B(\datapath.aluinstr [8]),
    .Y(_14_)
);

XOR2X1 _9587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_15_bF$buf26 ),
    .B(\datapath.aluinstr [7]),
    .Y(_15_)
);

XOR2X1 _9588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_17_bF$buf19 ),
    .B(\datapath.aluinstr [9]),
    .Y(_16_)
);

NOR3X1 _9589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_14_),
    .B(_15_),
    .C(_16_),
    .Y(_17_)
);

NOR2X1 _9590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.aluinstr [3]),
    .B(\datapath.aluinstr [2]),
    .Y(_18_)
);

INVX1 _9591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.aluinstr [5]),
    .Y(_19_)
);

NOR2X1 _9592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.aluinstr [4]),
    .B(_19_),
    .Y(_20_)
);

AND2X2 _9593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_19_bF$buf2 ),
    .B(\datapath.aluinstr [11]),
    .Y(_21_)
);

NOR2X1 _9594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_19_bF$buf1 ),
    .B(\datapath.aluinstr [11]),
    .Y(_22_)
);

AND2X2 _9595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_18_bF$buf7 ),
    .B(\datapath.aluinstr [10]),
    .Y(_23_)
);

NOR2X1 _9596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_18_bF$buf6 ),
    .B(\datapath.aluinstr [10]),
    .Y(_24_)
);

OAI22X1 _9597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_21_),
    .B(_22_),
    .C(_23_),
    .D(_24_),
    .Y(_25_)
);

AOI21X1 _9598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_18_),
    .B(_20_),
    .C(_25_),
    .Y(_26_)
);

NAND2X1 _9599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_26_),
    .B(_17_),
    .Y(_27_)
);

INVX1 _9600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_27_),
    .Y(_28_)
);

OR2X2 _9601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_28_),
    .B(_13_),
    .Y(_29_)
);

AOI21X1 _9602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_125_),
    .B(_137_),
    .C(_29_),
    .Y(abpsel[0])
);

AOI21X1 _9603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_27_),
    .B(_125_),
    .C(_13_),
    .Y(abpsel[1])
);

NAND2X1 _9604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_108_),
    .B(_27_),
    .Y(_30_)
);

OR2X2 _9605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_124_),
    .B(_13_),
    .Y(_31_)
);

NOR2X1 _9606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_30_),
    .B(_31_),
    .Y(abpsel[2])
);

INVX1 _9607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_23_bF$buf1 ),
    .Y(_32_)
);

NOR2X1 _9608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf33 ),
    .B(\datapath.idinstr_21_bF$buf13 ),
    .Y(_33_)
);

NOR2X1 _9609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf20 ),
    .B(\datapath.idinstr_24_bF$buf4 ),
    .Y(_34_)
);

NAND3X1 _9610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_32_),
    .B(_33_),
    .C(_34_),
    .Y(_35_)
);

INVX1 _9611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [4]),
    .Y(_36_)
);

AOI21X1 _9612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3_),
    .B(_36_),
    .C(_138_),
    .Y(_37_)
);

NAND2X1 _9613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [5]),
    .B(_6_),
    .Y(_38_)
);

NOR3X1 _9614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7_),
    .B(_38_),
    .C(_37_),
    .Y(_39_)
);

NAND2X1 _9615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_35_),
    .B(_39_),
    .Y(_40_)
);

XOR2X1 _9616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [11]),
    .B(\datapath.idinstr_24_bF$buf3 ),
    .Y(_41_)
);

INVX1 _9617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf12 ),
    .Y(_42_)
);

OAI22X1 _9618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_42_),
    .B(\datapath.meminstr [8]),
    .C(\datapath.meminstr [10]),
    .D(_32_),
    .Y(_43_)
);

NOR2X1 _9619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_43_),
    .B(_41_),
    .Y(_44_)
);

OAI22X1 _9620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114_),
    .B(\datapath.idinstr_22_bF$buf19 ),
    .C(_111_),
    .D(\datapath.idinstr_23_bF$buf0 ),
    .Y(_45_)
);

INVX1 _9621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_22_bF$buf18 ),
    .Y(_46_)
);

OAI22X1 _9622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_110_),
    .B(\datapath.idinstr_21_bF$buf11 ),
    .C(\datapath.meminstr [9]),
    .D(_46_),
    .Y(_47_)
);

NOR2X1 _9623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_45_),
    .B(_47_),
    .Y(_48_)
);

XOR2X1 _9624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [7]),
    .B(\datapath.idinstr_20_bF$buf32 ),
    .Y(_49_)
);

NOR2X1 _9625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_49_),
    .B(_121_),
    .Y(_50_)
);

AND2X2 _9626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_50_),
    .B(_48_),
    .Y(_51_)
);

XNOR2X1 _9627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [11]),
    .B(\datapath.idinstr_24_bF$buf2 ),
    .Y(_52_)
);

XNOR2X1 _9628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [10]),
    .B(\datapath.idinstr_23_bF$buf7 ),
    .Y(_53_)
);

INVX1 _9629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [9]),
    .Y(_54_)
);

AOI22X1 _9630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_54_),
    .B(\datapath.idinstr_22_bF$buf17 ),
    .C(\datapath.wbinstr [8]),
    .D(_42_),
    .Y(_55_)
);

NAND3X1 _9631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_55_),
    .B(_52_),
    .C(_53_),
    .Y(_56_)
);

INVX1 _9632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [8]),
    .Y(_57_)
);

INVX1 _9633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf31 ),
    .Y(_58_)
);

AOI22X1 _9634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_57_),
    .B(\datapath.idinstr_21_bF$buf10 ),
    .C(\datapath.wbinstr [7]),
    .D(_58_),
    .Y(_59_)
);

INVX1 _9635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [7]),
    .Y(_60_)
);

AOI22X1 _9636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_60_),
    .B(\datapath.idinstr_20_bF$buf30 ),
    .C(\datapath.wbinstr [9]),
    .D(_46_),
    .Y(_61_)
);

NAND3X1 _9637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_59_),
    .B(_61_),
    .C(_132_),
    .Y(_62_)
);

NOR2X1 _9638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_56_),
    .B(_62_),
    .Y(_63_)
);

AOI21X1 _9639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_44_),
    .B(_51_),
    .C(_63_),
    .Y(_64_)
);

NAND2X1 _9640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_104_),
    .B(_107_),
    .Y(_65_)
);

NAND3X1 _9641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_44_),
    .B(_48_),
    .C(_50_),
    .Y(_66_)
);

XOR2X1 _9642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.aluinstr [11]),
    .B(\datapath.idinstr_24_bF$buf1 ),
    .Y(_67_)
);

XOR2X1 _9643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.aluinstr [9]),
    .B(\datapath.idinstr_22_bF$buf16 ),
    .Y(_68_)
);

XOR2X1 _9644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.aluinstr [7]),
    .B(\datapath.idinstr_20_bF$buf29 ),
    .Y(_69_)
);

NOR3X1 _9645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_67_),
    .B(_68_),
    .C(_69_),
    .Y(_70_)
);

AND2X2 _9646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.aluinstr [10]),
    .B(\datapath.idinstr_23_bF$buf6 ),
    .Y(_71_)
);

NOR2X1 _9647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.aluinstr [10]),
    .B(\datapath.idinstr_23_bF$buf5 ),
    .Y(_72_)
);

AND2X2 _9648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.aluinstr [8]),
    .B(\datapath.idinstr_21_bF$buf9 ),
    .Y(_73_)
);

NOR2X1 _9649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.aluinstr [8]),
    .B(\datapath.idinstr_21_bF$buf8 ),
    .Y(_74_)
);

OAI22X1 _9650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_71_),
    .B(_72_),
    .C(_73_),
    .D(_74_),
    .Y(_75_)
);

AOI21X1 _9651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_18_),
    .B(_20_),
    .C(_75_),
    .Y(_76_)
);

NAND2X1 _9652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_76_),
    .B(_70_),
    .Y(_77_)
);

OAI21X1 _9653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_66_),
    .B(_65_),
    .C(_77_),
    .Y(_78_)
);

NOR3X1 _9654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_78_),
    .B(_40_),
    .C(_64_),
    .Y(bbpsel[0])
);

OR2X2 _9655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_66_),
    .B(_108_),
    .Y(_79_)
);

AOI21X1 _9656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_77_),
    .B(_79_),
    .C(_40_),
    .Y(bbpsel[1])
);

INVX1 _9657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_77_),
    .Y(_80_)
);

OR2X2 _9658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_66_),
    .B(_65_),
    .Y(_81_)
);

NOR3X1 _9659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_40_),
    .B(_80_),
    .C(_81_),
    .Y(bbpsel[2])
);

NAND3X1 _9660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_138_),
    .B(_3_),
    .C(_36_),
    .Y(_82_)
);

NOR2X1 _9661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_38_),
    .B(_82_),
    .Y(_83_)
);

NAND2X1 _9662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_35_),
    .B(_83_),
    .Y(_84_)
);

NOR3X1 _9663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_78_),
    .B(_84_),
    .C(_64_),
    .Y(\bypassandflushunit.rs2_bypass_sel [0])
);

AOI21X1 _9664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_77_),
    .B(_79_),
    .C(_84_),
    .Y(\bypassandflushunit.rs2_bypass_sel [1])
);

NOR3X1 _9665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_80_),
    .B(_84_),
    .C(_81_),
    .Y(\bypassandflushunit.rs2_bypass_sel [2])
);

NOR2X1 _9666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.regwbtrap ),
    .B(\datapath.regmret_bF$buf2 ),
    .Y(_85_)
);

INVX4 _9667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .Y(\bypassandflushunit.flushsystem )
);

NAND2X1 _9668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [4]),
    .B(\datapath.meminstr [5]),
    .Y(_86_)
);

NOR2X1 _9669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_86_),
    .B(_106_),
    .Y(_87_)
);

NAND2X1 _9670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [5]),
    .B(_131_),
    .Y(_88_)
);

NAND2X1 _9671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.aluinstr [5]),
    .B(_18_),
    .Y(_89_)
);

NAND2X1 _9672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [6]),
    .B(\datapath.wbinstr [4]),
    .Y(_90_)
);

NAND2X1 _9673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.aluinstr [4]),
    .B(\datapath.aluinstr [6]),
    .Y(_91_)
);

OAI22X1 _9674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_88_),
    .B(_90_),
    .C(_89_),
    .D(_91_),
    .Y(_92_)
);

AOI21X1 _9675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [6]),
    .B(_87_),
    .C(_92_),
    .Y(_93_)
);

NOR2X1 _9676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.aluinstr [4]),
    .B(\datapath.aluinstr [6]),
    .Y(_94_)
);

NAND2X1 _9677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_18_),
    .B(_94_),
    .Y(_95_)
);

NOR2X1 _9678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.aluinstr [5]),
    .B(_95_),
    .Y(_96_)
);

OAI21X1 _9679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_39_),
    .B(_83_),
    .C(_35_),
    .Y(_97_)
);

OAI22X1 _9680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_27_),
    .B(_13_),
    .C(_97_),
    .D(_77_),
    .Y(_98_)
);

NAND2X1 _9681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96_),
    .B(_98_),
    .Y(_99_)
);

NAND2X1 _9682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_99_),
    .Y(\bypassandflushunit.stall )
);

NAND2X1 _9683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [2]),
    .B(\datapath.meminstr [6]),
    .Y(_100_)
);

NOR2X1 _9684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_100_),
    .B(_120_),
    .Y(_101_)
);

OR2X2 _9685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.flushsystem ),
    .B(branch),
    .Y(_102_)
);

NOR2X1 _9686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_101_),
    .B(_102_),
    .Y(_103_)
);

INVX4 _9687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_103_),
    .Y(\bypassandflushunit.flushid )
);

NAND3X1 _9688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_103_),
    .C(_99_),
    .Y(\bypassandflushunit.flushalu )
);

NOR2X1 _9689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [3]),
    .B(\datapath.meminstr [2]),
    .Y(_220_)
);

NAND3X1 _9690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [1]),
    .B(\datapath.meminstr [0]),
    .C(_220_),
    .Y(_221_)
);

INVX1 _9691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [6]),
    .Y(_222_)
);

NOR2X1 _9692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.csrfile_trap_wen ),
    .B(\datapath.meminstr [4]),
    .Y(_223_)
);

NAND3X1 _9693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [5]),
    .B(_222_),
    .C(_223_),
    .Y(_224_)
);

NOR2X1 _9694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_221_),
    .B(_224_),
    .Y(_2_)
);

OR2X2 _9695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [13]),
    .B(\datapath.meminstr [14]),
    .Y(_225_)
);

NOR2X1 _9696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [12]),
    .B(_225_),
    .Y(_226_)
);

INVX1 _9697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\controlunit.csrfile_trap_wen ),
    .Y(_227_)
);

AND2X2 _9698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [5]),
    .B(\datapath.meminstr [6]),
    .Y(_228_)
);

NAND3X1 _9699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_227_),
    .B(\datapath.meminstr [4]),
    .C(_228_),
    .Y(_229_)
);

OR2X2 _9700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_229_),
    .B(_221_),
    .Y(_230_)
);

NOR2X1 _9701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_226_),
    .B(_230_),
    .Y(\controlunit.csrfile_wen )
);

INVX1 _9702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [21]),
    .Y(_231_)
);

NOR2X1 _9703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [20]),
    .B(_231_),
    .Y(_232_)
);

NAND3X1 _9704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [29]),
    .B(_232_),
    .C(_226_),
    .Y(_233_)
);

NOR2X1 _9705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_233_),
    .B(_230_),
    .Y(\controlunit.mret )
);

INVX1 _9706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [3]),
    .Y(_234_)
);

NAND3X1 _9707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [1]),
    .B(\datapath.wbinstr [0]),
    .C(_234_),
    .Y(_235_)
);

NOR2X1 _9708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [2]),
    .B(_235_),
    .Y(_236_)
);

INVX2 _9709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [4]),
    .Y(_237_)
);

NAND2X1 _9710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [6]),
    .B(\datapath.wbinstr [5]),
    .Y(_238_)
);

OR2X2 _9711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_238_),
    .B(_237_),
    .Y(_239_)
);

INVX1 _9712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_239_),
    .Y(_240_)
);

INVX1 _9713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [12]),
    .Y(_241_)
);

NOR2X1 _9714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [13]),
    .B(\datapath.wbinstr [14]),
    .Y(_242_)
);

NAND2X1 _9715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_241_),
    .B(_242_),
    .Y(_243_)
);

NAND3X1 _9716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_243_),
    .B(_236_),
    .C(_240_),
    .Y(_244_)
);

NAND3X1 _9717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [1]),
    .B(\datapath.wbinstr [0]),
    .C(\datapath.wbinstr [2]),
    .Y(_245_)
);

NOR2X1 _9718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_238_),
    .B(_245_),
    .Y(_246_)
);

OR2X2 _9719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237_),
    .B(\datapath.wbinstr [6]),
    .Y(_247_)
);

NOR2X1 _9720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [5]),
    .B(\datapath.wbinstr [4]),
    .Y(_139_)
);

NOR2X1 _9721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.wbinstr [2]),
    .B(\datapath.wbinstr [6]),
    .Y(_140_)
);

NAND2X1 _9722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_139_),
    .B(_140_),
    .Y(_141_)
);

AOI21X1 _9723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_141_),
    .B(_247_),
    .C(_235_),
    .Y(_142_)
);

AOI21X1 _9724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237_),
    .B(_246_),
    .C(_142_),
    .Y(_143_)
);

AOI21X1 _9725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_244_),
    .B(_143_),
    .C(\datapath.regwbtrap ),
    .Y(\controlunit.regfile_wen )
);

INVX2 _9726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [13]),
    .Y(_144_)
);

INVX1 _9727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [12]),
    .Y(_145_)
);

NOR2X1 _9728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [2]),
    .B(\datapath.idinstr [3]),
    .Y(_146_)
);

NAND3X1 _9729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [1]),
    .B(\datapath.idinstr [0]),
    .C(_146_),
    .Y(_147_)
);

INVX2 _9730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [4]),
    .Y(_148_)
);

NAND3X1 _9731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [6]),
    .B(\datapath.idinstr [5]),
    .C(_148_),
    .Y(_149_)
);

NOR2X1 _9732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_149_),
    .B(_147_),
    .Y(_150_)
);

INVX1 _9733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_150_),
    .Y(_151_)
);

NAND3X1 _9734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [6]),
    .B(\datapath.idinstr [4]),
    .C(\datapath.idinstr [5]),
    .Y(_152_)
);

NOR2X1 _9735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_152_),
    .B(_147_),
    .Y(_153_)
);

INVX2 _9736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [6]),
    .Y(_154_)
);

NAND2X1 _9737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [4]),
    .B(_154_),
    .Y(_155_)
);

NOR2X1 _9738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_155_),
    .B(_147_),
    .Y(_156_)
);

AOI21X1 _9739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [13]),
    .B(_153_),
    .C(_156_),
    .Y(_157_)
);

OAI22X1 _9740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_144_),
    .B(_151_),
    .C(_157_),
    .D(_145_),
    .Y(alusel[0])
);

NOR3X1 _9741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [6]),
    .B(\datapath.idinstr [5]),
    .C(_148_),
    .Y(_158_)
);

NAND3X1 _9742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [1]),
    .B(\datapath.idinstr [0]),
    .C(\datapath.idinstr [2]),
    .Y(_159_)
);

NOR2X1 _9743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [3]),
    .B(_159_),
    .Y(_160_)
);

NAND2X1 _9744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_158_),
    .B(_160_),
    .Y(_161_)
);

NAND2X1 _9745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [1]),
    .B(\datapath.idinstr [0]),
    .Y(_162_)
);

NOR3X1 _9746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [2]),
    .B(\datapath.idinstr [3]),
    .C(_162_),
    .Y(_163_)
);

INVX2 _9747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [5]),
    .Y(_164_)
);

NOR3X1 _9748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_154_),
    .B(\datapath.idinstr [4]),
    .C(_164_),
    .Y(_165_)
);

INVX2 _9749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_152_),
    .Y(_166_)
);

OAI21X1 _9750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_165_),
    .B(_166_),
    .C(_163_),
    .Y(_167_)
);

AOI22X1 _9751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_160_),
    .B(_165_),
    .C(_154_),
    .D(_163_),
    .Y(_168_)
);

NAND3X1 _9752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_161_),
    .B(_167_),
    .C(_168_),
    .Y(_169_)
);

OAI21X1 _9753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_150_),
    .B(_153_),
    .C(\datapath.idinstr [14]),
    .Y(_170_)
);

OAI21X1 _9754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_153_),
    .B(_156_),
    .C(\datapath.idinstr [13]),
    .Y(_171_)
);

NAND3X1 _9755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .B(_171_),
    .C(_169_),
    .Y(alusel[1])
);

AOI21X1 _9756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [14]),
    .B(_156_),
    .C(_153_),
    .Y(_172_)
);

NAND2X1 _9757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172_),
    .B(_169_),
    .Y(alusel[2])
);

NAND2X1 _9758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [13]),
    .B(_145_),
    .Y(_173_)
);

AOI21X1 _9759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_173_),
    .B(_153_),
    .C(_150_),
    .Y(_174_)
);

INVX1 _9760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [30]),
    .Y(_175_)
);

NAND3X1 _9761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [4]),
    .B(\datapath.idinstr [5]),
    .C(_154_),
    .Y(_176_)
);

NOR3X1 _9762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_175_),
    .B(_176_),
    .C(_147_),
    .Y(_177_)
);

AND2X2 _9763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [12]),
    .B(\datapath.idinstr [30]),
    .Y(_178_)
);

NAND3X1 _9764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_144_),
    .B(\datapath.idinstr [14]),
    .C(_178_),
    .Y(_179_)
);

NOR2X1 _9765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_147_),
    .B(_179_),
    .Y(_180_)
);

AOI21X1 _9766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_158_),
    .B(_180_),
    .C(_177_),
    .Y(_181_)
);

NAND3X1 _9767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_174_),
    .B(_181_),
    .C(_169_),
    .Y(alusel[3])
);

INVX1 _9768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.aluinstr [4]),
    .Y(_182_)
);

NAND3X1 _9769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.aluinstr [5]),
    .B(\datapath.aluinstr [6]),
    .C(_182_),
    .Y(_183_)
);

NAND3X1 _9770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.aluinstr [1]),
    .B(\datapath.aluinstr [0]),
    .C(\datapath.aluinstr [2]),
    .Y(_184_)
);

INVX1 _9771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_184_),
    .Y(_185_)
);

NAND2X1 _9772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.aluinstr [3]),
    .B(_185_),
    .Y(_186_)
);

NOR2X1 _9773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_183_),
    .B(_186_),
    .Y(\controlunit.pc_sel [0])
);

OR2X2 _9774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_184_),
    .B(\datapath.aluinstr [3]),
    .Y(_187_)
);

NOR2X1 _9775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_183_),
    .B(_187_),
    .Y(\controlunit.pc_sel [1])
);

NAND2X1 _9776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_166_),
    .B(_163_),
    .Y(_188_)
);

NOR3X1 _9777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [6]),
    .B(\datapath.idinstr [4]),
    .C(_164_),
    .Y(_189_)
);

NAND2X1 _9778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_189_),
    .B(_163_),
    .Y(_190_)
);

INVX1 _9779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_155_),
    .Y(_191_)
);

NAND2X1 _9780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_160_),
    .B(_191_),
    .Y(_192_)
);

NAND3X1 _9781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(_192_),
    .C(_167_),
    .Y(_193_)
);

NOR2X1 _9782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [6]),
    .B(\datapath.idinstr [5]),
    .Y(_194_)
);

AND2X2 _9783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_194_),
    .B(_148_),
    .Y(_195_)
);

INVX1 _9784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [3]),
    .Y(_196_)
);

NOR2X1 _9785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_196_),
    .B(_159_),
    .Y(_197_)
);

OAI21X1 _9786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_163_),
    .B(_197_),
    .C(_195_),
    .Y(_198_)
);

INVX1 _9787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_159_),
    .Y(_199_)
);

AOI22X1 _9788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_165_),
    .B(_199_),
    .C(_191_),
    .D(_163_),
    .Y(_200_)
);

NAND2X1 _9789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_198_),
    .B(_200_),
    .Y(_201_)
);

INVX1 _9790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf28 ),
    .Y(_202_)
);

NAND3X1 _9791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf7 ),
    .B(\datapath.idinstr [29]),
    .C(_202_),
    .Y(_203_)
);

OR2X2 _9792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_21_bF$buf6 ),
    .B(\datapath.idinstr [29]),
    .Y(_204_)
);

INVX2 _9793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [14]),
    .Y(_205_)
);

NAND2X1 _9794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_144_),
    .B(_205_),
    .Y(_206_)
);

NOR2X1 _9795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [12]),
    .B(_206_),
    .Y(_207_)
);

NAND3X1 _9796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_204_),
    .B(_203_),
    .C(_207_),
    .Y(_208_)
);

OAI22X1 _9797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_188_),
    .B(_208_),
    .C(_193_),
    .D(_201_),
    .Y(\controlunit.ill_op )
);

NAND2X1 _9798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_236_),
    .B(_240_),
    .Y(_209_)
);

OAI21X1 _9799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_235_),
    .B(_141_),
    .C(_209_),
    .Y(\controlunit.wb_sel [0])
);

INVX1 _9800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_142_),
    .Y(\controlunit.wb_sel [1])
);

NAND2X1 _9801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_165_),
    .B(_197_),
    .Y(_210_)
);

OAI21X1 _9802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_147_),
    .B(_152_),
    .C(_210_),
    .Y(\controlunit.imm_sel [2])
);

NAND2X1 _9803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_165_),
    .B(_160_),
    .Y(_211_)
);

NAND2X1 _9804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_194_),
    .B(_163_),
    .Y(_212_)
);

OAI21X1 _9805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_165_),
    .B(_189_),
    .C(_163_),
    .Y(_213_)
);

NAND3X1 _9806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_211_),
    .B(_212_),
    .C(_213_),
    .Y(_214_)
);

OAI21X1 _9807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_189_),
    .B(_166_),
    .C(_163_),
    .Y(_215_)
);

OAI21X1 _9808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_214_),
    .B(\controlunit.imm_sel [2]),
    .C(_215_),
    .Y(\controlunit.imm_sel [0])
);

OAI21X1 _9809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_214_),
    .B(\controlunit.imm_sel [2]),
    .C(_151_),
    .Y(\controlunit.imm_sel [1])
);

OAI21X1 _9810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_147_),
    .B(_176_),
    .C(_167_),
    .Y(_216_)
);

OAI21X1 _9811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_205_),
    .B(_188_),
    .C(_216_),
    .Y(bsel[0])
);

NOR2X1 _9812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [14]),
    .B(_188_),
    .Y(bsel[1])
);

AND2X2 _9813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_168_),
    .B(_167_),
    .Y(asel[0])
);

NOR2X1 _9814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_205_),
    .B(_188_),
    .Y(asel[1])
);

OR2X2 _9815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_188_),
    .B(_204_),
    .Y(_217_)
);

NAND2X1 _9816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr_20_bF$buf27 ),
    .B(_207_),
    .Y(_218_)
);

NOR2X1 _9817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_218_),
    .B(_217_),
    .Y(\controlunit.ebreak )
);

NAND2X1 _9818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_202_),
    .B(_207_),
    .Y(_219_)
);

NOR2X1 _9819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_219_),
    .B(_217_),
    .Y(\controlunit.ecall )
);

INVX8 _9820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.flushid ),
    .Y(_254_)
);

AND2X2 _9821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf2),
    .B(\controlunit.pc_sel [0]),
    .Y(\datapath._32_ [0])
);

AND2X2 _9822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254__bF$buf1),
    .B(\controlunit.pc_sel [1]),
    .Y(\datapath._32_ [1])
);

INVX4 _9823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.flushsystem ),
    .Y(_255_)
);

INVX1 _9824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [0]),
    .Y(_256_)
);

NAND2X1 _9825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(_256_),
    .Y(\datapath._49_ [0])
);

INVX1 _9826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [1]),
    .Y(_257_)
);

NAND2X1 _9827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(_257_),
    .Y(\datapath._49_ [1])
);

INVX1 _9828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [2]),
    .Y(_258_)
);

NOR2X1 _9829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.flushsystem ),
    .B(_258_),
    .Y(\datapath._49_ [2])
);

INVX1 _9830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [3]),
    .Y(_259_)
);

NOR2X1 _9831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.flushsystem ),
    .B(_259_),
    .Y(\datapath._49_ [3])
);

OR2X2 _9832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.flushsystem ),
    .B(\datapath.meminstr [4]),
    .Y(\datapath._49_ [4])
);

INVX2 _9833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [5]),
    .Y(_260_)
);

NOR2X1 _9834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.flushsystem ),
    .B(_260_),
    .Y(\datapath._49_ [5])
);

AND2X2 _9835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(\datapath.meminstr [6]),
    .Y(\datapath._49_ [6])
);

AND2X2 _9836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(\datapath.meminstr [7]),
    .Y(\datapath._49_ [7])
);

AND2X2 _9837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(\datapath.meminstr [8]),
    .Y(\datapath._49_ [8])
);

AND2X2 _9838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(\datapath.meminstr [9]),
    .Y(\datapath._49_ [9])
);

AND2X2 _9839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(\datapath.meminstr [10]),
    .Y(\datapath._49_ [10])
);

AND2X2 _9840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(\datapath.meminstr [11]),
    .Y(\datapath._49_ [11])
);

AND2X2 _9841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(\datapath.meminstr [12]),
    .Y(\datapath._49_ [12])
);

INVX2 _9842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [13]),
    .Y(_261_)
);

NOR2X1 _9843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.flushsystem ),
    .B(_261_),
    .Y(\datapath._49_ [13])
);

AND2X2 _9844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(\datapath.meminstr [14]),
    .Y(\datapath._49_ [14])
);

AND2X2 _9845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(\controlunit.csrfile_trap_wen ),
    .Y(\datapath._50_ )
);

AND2X2 _9846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(\controlunit.mret ),
    .Y(\datapath._51_ )
);

NOR2X1 _9847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [4]),
    .B(_260_),
    .Y(_262_)
);

NAND2X1 _9848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [6]),
    .B(_262_),
    .Y(_263_)
);

NOR2X1 _9849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_256_),
    .B(_257_),
    .Y(_264_)
);

NAND2X1 _9850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_259_),
    .B(_264_),
    .Y(_265_)
);

NOR2X1 _9851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [2]),
    .B(_265_),
    .Y(_266_)
);

NAND2X1 _9852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.tkbranch ),
    .B(_266_),
    .Y(_267_)
);

NOR2X1 _9853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_263_),
    .B(_267_),
    .Y(branch)
);

INVX1 _9854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0__1_bF$buf4),
    .Y(_268_)
);

OAI21X1 _9855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [12]),
    .B(\datapath.meminstr [13]),
    .C(_0__0_bF$buf3),
    .Y(_269_)
);

OAI21X1 _9856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_261_),
    .B(_268_),
    .C(_269_),
    .Y(_270_)
);

NOR2X1 _9857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [4]),
    .B(\datapath.meminstr [6]),
    .Y(_271_)
);

NAND3X1 _9858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_270_),
    .B(_271_),
    .C(_266_),
    .Y(_272_)
);

NOR2X1 _9859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.jumps [1]),
    .B(\datapath.programcounter.jumps [0]),
    .Y(_273_)
);

INVX1 _9860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_263_),
    .Y(_274_)
);

INVX1 _9861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_265_),
    .Y(_275_)
);

NOR2X1 _9862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_258_),
    .B(_268_),
    .Y(_276_)
);

NAND3X1 _9863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_276_),
    .B(_274_),
    .C(_275_),
    .Y(_277_)
);

INVX1 _9864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_264_),
    .Y(_278_)
);

NAND2X1 _9865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.meminstr [2]),
    .B(\datapath.meminstr [3]),
    .Y(_279_)
);

OAI21X1 _9866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_278_),
    .B(_279_),
    .C(_267_),
    .Y(_280_)
);

NAND2X1 _9867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_274_),
    .B(_280_),
    .Y(_281_)
);

OAI21X1 _9868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_281_),
    .B(_273_),
    .C(_277_),
    .Y(_282_)
);

NOR2X1 _9869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memexecptions [0]),
    .B(\datapath.memexecptions [2]),
    .Y(_283_)
);

NOR2X1 _9870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_irq ),
    .B(\datapath.memexecptions [1]),
    .Y(_284_)
);

NAND2X1 _9871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_283_),
    .B(_284_),
    .Y(_285_)
);

NOR2X1 _9872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_285_),
    .B(_282_),
    .Y(\datapath.excpt_cause [2])
);

NAND2X1 _9873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_),
    .B(\datapath.excpt_cause [2]),
    .Y(\controlunit.csrfile_trap_wen )
);

AOI21X1 _9874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_),
    .B(\datapath.excpt_cause [2]),
    .C(\bypassandflushunit.flushsystem ),
    .Y(\datapath._52_ )
);

INVX1 _9875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.memexecptions [0]),
    .Y(_286_)
);

INVX1 _9876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_282_),
    .Y(_287_)
);

NAND3X1 _9877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_286_),
    .B(\datapath.memexecptions [2]),
    .C(_287_),
    .Y(_288_)
);

NAND2X1 _9878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_284_),
    .B(_288_),
    .Y(\datapath.excpt_cause [0])
);

INVX1 _9879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_285_),
    .Y(_289_)
);

OR2X2 _9880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_),
    .B(_260_),
    .Y(_290_)
);

AOI22X1 _9881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_289_),
    .B(_290_),
    .C(_282_),
    .D(_284_),
    .Y(\datapath.excpt_cause [1])
);

INVX1 _9882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.csr.csr_irq ),
    .Y(_291_)
);

OAI21X1 _9883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_288_),
    .B(\datapath.memexecptions [1]),
    .C(_291_),
    .Y(\datapath.excpt_cause [3])
);

INVX1 _9884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IMEM_DATA[0]),
    .Y(_292_)
);

AOI21X1 _9885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idinstr [0]),
    .B(\bypassandflushunit.stall_bF$buf5 ),
    .C(\bypassandflushunit.flushid ),
    .Y(_293_)
);

OAI21X1 _9886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_292_),
    .B(\bypassandflushunit.stall_bF$buf4 ),
    .C(_293_),
    .Y(\datapath._03_ [0])
);

INVX1 _9887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IMEM_DATA[1]),
    .Y(_294_)
);

AOI21X1 _9888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf3 ),
    .B(\datapath.idinstr [1]),
    .C(\bypassandflushunit.flushid ),
    .Y(_295_)
);

OAI21X1 _9889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf2 ),
    .B(_294_),
    .C(_295_),
    .Y(\datapath._03_ [1])
);

NOR2X1 _9890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf1 ),
    .B(IMEM_DATA[2]),
    .Y(_296_)
);

INVX8 _9891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf0 ),
    .Y(_297_)
);

INVX8 _9892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.flushid ),
    .Y(_298_)
);

OAI21X1 _9893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf0),
    .B(\datapath.idinstr [2]),
    .C(_298__bF$buf4),
    .Y(_299_)
);

NOR2X1 _9894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_296_),
    .B(_299_),
    .Y(\datapath._03_ [2])
);

NOR2X1 _9895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf9 ),
    .B(IMEM_DATA[3]),
    .Y(_300_)
);

OAI21X1 _9896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf8),
    .B(\datapath.idinstr [3]),
    .C(_298__bF$buf3),
    .Y(_301_)
);

NOR2X1 _9897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_300_),
    .B(_301_),
    .Y(\datapath._03_ [3])
);

INVX1 _9898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(IMEM_DATA[4]),
    .Y(_302_)
);

AOI21X1 _9899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf8 ),
    .B(\datapath.idinstr [4]),
    .C(\bypassandflushunit.flushid ),
    .Y(_303_)
);

OAI21X1 _9900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf7 ),
    .B(_302_),
    .C(_303_),
    .Y(\datapath._03_ [4])
);

NOR2X1 _9901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf6 ),
    .B(IMEM_DATA[5]),
    .Y(_304_)
);

OAI21X1 _9902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf7),
    .B(\datapath.idinstr [5]),
    .C(_298__bF$buf2),
    .Y(_305_)
);

NOR2X1 _9903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_304_),
    .B(_305_),
    .Y(\datapath._03_ [5])
);

NOR2X1 _9904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf5 ),
    .B(IMEM_DATA[6]),
    .Y(_306_)
);

OAI21X1 _9905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf6),
    .B(\datapath.idinstr [6]),
    .C(_298__bF$buf1),
    .Y(_307_)
);

NOR2X1 _9906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_306_),
    .B(_307_),
    .Y(\datapath._03_ [6])
);

NOR2X1 _9907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf4 ),
    .B(IMEM_DATA[7]),
    .Y(_308_)
);

OAI21X1 _9908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf5),
    .B(\datapath.idinstr [7]),
    .C(_298__bF$buf0),
    .Y(_309_)
);

NOR2X1 _9909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_308_),
    .B(_309_),
    .Y(\datapath._03_ [7])
);

NOR2X1 _9910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf3 ),
    .B(IMEM_DATA[8]),
    .Y(_310_)
);

OAI21X1 _9911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf4),
    .B(\datapath.idinstr [8]),
    .C(_298__bF$buf4),
    .Y(_311_)
);

NOR2X1 _9912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_310_),
    .B(_311_),
    .Y(\datapath._03_ [8])
);

NOR2X1 _9913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf2 ),
    .B(IMEM_DATA[9]),
    .Y(_312_)
);

OAI21X1 _9914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf3),
    .B(\datapath.idinstr [9]),
    .C(_298__bF$buf3),
    .Y(_313_)
);

NOR2X1 _9915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_312_),
    .B(_313_),
    .Y(\datapath._03_ [9])
);

NOR2X1 _9916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf1 ),
    .B(IMEM_DATA[10]),
    .Y(_314_)
);

OAI21X1 _9917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf2),
    .B(\datapath.idinstr [10]),
    .C(_298__bF$buf2),
    .Y(_315_)
);

NOR2X1 _9918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_314_),
    .B(_315_),
    .Y(\datapath._03_ [10])
);

NOR2X1 _9919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf0 ),
    .B(IMEM_DATA[11]),
    .Y(_316_)
);

OAI21X1 _9920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf1),
    .B(\datapath.idinstr [11]),
    .C(_298__bF$buf1),
    .Y(_317_)
);

NOR2X1 _9921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_316_),
    .B(_317_),
    .Y(\datapath._03_ [11])
);

NOR2X1 _9922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf9 ),
    .B(IMEM_DATA[12]),
    .Y(_318_)
);

OAI21X1 _9923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf0),
    .B(\datapath.idinstr [12]),
    .C(_298__bF$buf0),
    .Y(_319_)
);

NOR2X1 _9924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_318_),
    .B(_319_),
    .Y(\datapath._03_ [12])
);

NOR2X1 _9925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf8 ),
    .B(IMEM_DATA[13]),
    .Y(_320_)
);

OAI21X1 _9926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf8),
    .B(\datapath.idinstr [13]),
    .C(_298__bF$buf4),
    .Y(_321_)
);

NOR2X1 _9927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_320_),
    .B(_321_),
    .Y(\datapath._03_ [13])
);

NOR2X1 _9928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf7 ),
    .B(IMEM_DATA[14]),
    .Y(_322_)
);

OAI21X1 _9929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf7),
    .B(\datapath.idinstr [14]),
    .C(_298__bF$buf3),
    .Y(_323_)
);

NOR2X1 _9930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_322_),
    .B(_323_),
    .Y(\datapath._03_ [14])
);

NOR2X1 _9931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf6 ),
    .B(IMEM_DATA[15]),
    .Y(_324_)
);

OAI21X1 _9932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf6),
    .B(\datapath.idinstr_15_bF$buf25 ),
    .C(_298__bF$buf2),
    .Y(_325_)
);

NOR2X1 _9933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_324_),
    .B(_325_),
    .Y(\datapath._03_ [15])
);

NOR2X1 _9934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf5 ),
    .B(IMEM_DATA[16]),
    .Y(_326_)
);

OAI21X1 _9935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf5),
    .B(\datapath.idinstr_16_bF$buf8 ),
    .C(_298__bF$buf1),
    .Y(_327_)
);

NOR2X1 _9936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_326_),
    .B(_327_),
    .Y(\datapath._03_ [16])
);

NOR2X1 _9937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf4 ),
    .B(IMEM_DATA[17]),
    .Y(_328_)
);

OAI21X1 _9938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf4),
    .B(\datapath.idinstr_17_bF$buf18 ),
    .C(_298__bF$buf0),
    .Y(_329_)
);

NOR2X1 _9939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_328_),
    .B(_329_),
    .Y(\datapath._03_ [17])
);

NOR2X1 _9940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf3 ),
    .B(IMEM_DATA[18]),
    .Y(_330_)
);

OAI21X1 _9941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf3),
    .B(\datapath.idinstr_18_bF$buf5 ),
    .C(_298__bF$buf4),
    .Y(_331_)
);

NOR2X1 _9942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_330_),
    .B(_331_),
    .Y(\datapath._03_ [18])
);

NOR2X1 _9943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf2 ),
    .B(IMEM_DATA[19]),
    .Y(_332_)
);

OAI21X1 _9944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf2),
    .B(\datapath.idinstr_19_bF$buf0 ),
    .C(_298__bF$buf3),
    .Y(_333_)
);

NOR2X1 _9945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_332_),
    .B(_333_),
    .Y(\datapath._03_ [19])
);

NOR2X1 _9946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf1 ),
    .B(IMEM_DATA[20]),
    .Y(_334_)
);

OAI21X1 _9947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf1),
    .B(\datapath.idinstr_20_bF$buf26 ),
    .C(_298__bF$buf2),
    .Y(_335_)
);

NOR2X1 _9948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_334_),
    .B(_335_),
    .Y(\datapath._03_ [20])
);

NOR2X1 _9949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf0 ),
    .B(IMEM_DATA[21]),
    .Y(_336_)
);

OAI21X1 _9950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf0),
    .B(\datapath.idinstr_21_bF$buf5 ),
    .C(_298__bF$buf1),
    .Y(_337_)
);

NOR2X1 _9951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_336_),
    .B(_337_),
    .Y(\datapath._03_ [21])
);

NOR2X1 _9952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf9 ),
    .B(IMEM_DATA[22]),
    .Y(_338_)
);

OAI21X1 _9953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf8),
    .B(\datapath.idinstr_22_bF$buf15 ),
    .C(_298__bF$buf0),
    .Y(_339_)
);

NOR2X1 _9954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_338_),
    .B(_339_),
    .Y(\datapath._03_ [22])
);

NOR2X1 _9955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf8 ),
    .B(IMEM_DATA[23]),
    .Y(_340_)
);

OAI21X1 _9956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf7),
    .B(\datapath.idinstr_23_bF$buf4 ),
    .C(_298__bF$buf4),
    .Y(_341_)
);

NOR2X1 _9957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_340_),
    .B(_341_),
    .Y(\datapath._03_ [23])
);

NOR2X1 _9958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf7 ),
    .B(IMEM_DATA[24]),
    .Y(_342_)
);

OAI21X1 _9959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf6),
    .B(\datapath.idinstr_24_bF$buf0 ),
    .C(_298__bF$buf3),
    .Y(_343_)
);

NOR2X1 _9960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_342_),
    .B(_343_),
    .Y(\datapath._03_ [24])
);

NOR2X1 _9961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf6 ),
    .B(IMEM_DATA[25]),
    .Y(_344_)
);

OAI21X1 _9962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf5),
    .B(\datapath.idinstr [25]),
    .C(_298__bF$buf2),
    .Y(_345_)
);

NOR2X1 _9963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_344_),
    .B(_345_),
    .Y(\datapath._03_ [25])
);

NOR2X1 _9964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf5 ),
    .B(IMEM_DATA[26]),
    .Y(_346_)
);

OAI21X1 _9965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf4),
    .B(\datapath.idinstr [26]),
    .C(_298__bF$buf1),
    .Y(_347_)
);

NOR2X1 _9966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_346_),
    .B(_347_),
    .Y(\datapath._03_ [26])
);

NOR2X1 _9967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf4 ),
    .B(IMEM_DATA[27]),
    .Y(_348_)
);

OAI21X1 _9968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf3),
    .B(\datapath.idinstr [27]),
    .C(_298__bF$buf0),
    .Y(_349_)
);

NOR2X1 _9969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_348_),
    .B(_349_),
    .Y(\datapath._03_ [27])
);

NOR2X1 _9970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf3 ),
    .B(IMEM_DATA[28]),
    .Y(_350_)
);

OAI21X1 _9971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf2),
    .B(\datapath.idinstr [28]),
    .C(_298__bF$buf4),
    .Y(_351_)
);

NOR2X1 _9972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_350_),
    .B(_351_),
    .Y(\datapath._03_ [28])
);

NOR2X1 _9973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf2 ),
    .B(IMEM_DATA[29]),
    .Y(_352_)
);

OAI21X1 _9974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf1),
    .B(\datapath.idinstr [29]),
    .C(_298__bF$buf3),
    .Y(_353_)
);

NOR2X1 _9975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_352_),
    .B(_353_),
    .Y(\datapath._03_ [29])
);

NOR2X1 _9976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf1 ),
    .B(IMEM_DATA[30]),
    .Y(_354_)
);

OAI21X1 _9977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf0),
    .B(\datapath.idinstr [30]),
    .C(_298__bF$buf2),
    .Y(_355_)
);

NOR2X1 _9978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_354_),
    .B(_355_),
    .Y(\datapath._03_ [30])
);

NOR2X1 _9979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\bypassandflushunit.stall_bF$buf0 ),
    .B(IMEM_DATA[31]),
    .Y(_356_)
);

OAI21X1 _9980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf8),
    .B(\datapath.idinstr [31]),
    .C(_298__bF$buf1),
    .Y(_357_)
);

NOR2X1 _9981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_356_),
    .B(_357_),
    .Y(\datapath._03_ [31])
);

INVX1 _9982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [0]),
    .Y(_358_)
);

NAND2X1 _9983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [0]),
    .B(_297__bF$buf7),
    .Y(_359_)
);

OAI21X1 _9984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf6),
    .B(_358_),
    .C(_359_),
    .Y(\datapath._05_ [0])
);

INVX1 _9985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [1]),
    .Y(_360_)
);

NAND2X1 _9986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [1]),
    .B(_297__bF$buf5),
    .Y(_361_)
);

OAI21X1 _9987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf4),
    .B(_360_),
    .C(_361_),
    .Y(\datapath._05_ [1])
);

INVX1 _9988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [2]),
    .Y(_362_)
);

NAND2X1 _9989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [2]),
    .B(_297__bF$buf3),
    .Y(_363_)
);

OAI21X1 _9990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf2),
    .B(_362_),
    .C(_363_),
    .Y(\datapath._05_ [2])
);

INVX1 _9991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [3]),
    .Y(_364_)
);

NAND2X1 _9992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [3]),
    .B(_297__bF$buf1),
    .Y(_365_)
);

OAI21X1 _9993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf0),
    .B(_364_),
    .C(_365_),
    .Y(\datapath._05_ [3])
);

INVX1 _9994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [4]),
    .Y(_366_)
);

NAND2X1 _9995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [4]),
    .B(_297__bF$buf8),
    .Y(_367_)
);

OAI21X1 _9996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf7),
    .B(_366_),
    .C(_367_),
    .Y(\datapath._05_ [4])
);

INVX1 _9997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.idpc [5]),
    .Y(_368_)
);

NAND2X1 _9998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\datapath.programcounter.pc [5]),
    .B(_297__bF$buf6),
    .Y(_369_)
);

OAI21X1 _9999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297__bF$buf5),
    .B(_368_),
    .C(_369_),
    .Y(\datapath._05_ [5])
);

endmodule
