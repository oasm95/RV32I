/* Verilog module written by vlogFanout (qflow) */
/* With clock tree generation and fanout reduction */
/* and gate resizing */

module csr(
    output CSR_IRQ,
    output [31:0] CSR_PCaddr,
    input CSR_Ret,
    input [31:0] CSR_Wdata,
    input CSR_Wen,
    input CSR_Wen_traps,
    input [11:0] CSR_addr,
    output [31:0] CSR_data,
    input [3:0] CSR_mcause,
    input [31:0] CSR_mepc,
    input Extern_IRQ,
    input clk
);

wire _168_ ;
wire _60_ ;
wire _397_ ;
wire _19_ ;
wire _321_ ;
wire _57_ ;
wire _130_ ;
wire _415_ ;
wire _95_ ;
wire _224_ ;
wire _453_ ;
wire _262_ ;
wire _318_ ;
wire _127_ ;
wire _356_ ;
wire _165_ ;
wire _394_ ;
wire _259_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _412_ ;
wire _92_ ;
wire _221_ ;
wire _450_ ;
wire _315_ ;
wire _124_ ;
wire _353_ ;
wire _409_ ;
wire _89_ ;
wire _162_ ;
wire _218_ ;
wire _391_ ;
wire _447_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _159_ ;
wire _51_ ;
wire _388_ ;
wire _197_ ;
wire _7_ ;
wire _312_ ;
wire _48_ ;
wire _121_ ;
wire _350_ ;
wire _406_ ;
wire _86_ ;
wire _215_ ;
wire _444_ ;
wire _253_ ;
wire _309_ ;
wire _482_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _347_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire [31:0] _07_ ;
wire _45_ ;
wire _403_ ;
wire _83_ ;
wire _212_ ;
wire _441_ ;
wire _250_ ;
wire _306_ ;
wire _115_ ;
wire _344_ ;
wire _153_ ;
wire _209_ ;
wire _382_ ;
wire _438_ ;
wire _191_ ;
wire _247_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire _285_ ;
wire _1_ ;
wire [1:0] mstatus ;
wire _42_ ;
wire _379_ ;
wire _188_ ;
wire _400_ ;
wire _80_ ;
wire _303_ ;
wire _39_ ;
wire _112_ ;
wire _341_ ;
wire clk ;
wire _77_ ;
wire _150_ ;
wire _206_ ;
wire _435_ ;
wire _244_ ;
wire _473_ ;
wire _109_ ;
wire _282_ ;
wire _338_ ;
wire CSR_IRQ ;
wire _147_ ;
wire _376_ ;
wire _235__bF$buf0 ;
wire _235__bF$buf1 ;
wire _235__bF$buf2 ;
wire _235__bF$buf3 ;
wire _235__bF$buf4 ;
wire _185_ ;
wire _279_ ;
wire _300_ ;
wire _36_ ;
wire _74_ ;
wire _203_ ;
wire _432_ ;
wire _241_ ;
wire _470_ ;
wire _106_ ;
wire _335_ ;
wire _144_ ;
wire _373_ ;
wire _429_ ;
wire _182_ ;
wire _238_ ;
wire _467_ ;
wire _276_ ;
wire [1:0] _33_ ;
wire _179_ ;
wire _71_ ;
wire _200_ ;
wire _103_ ;
wire _332_ ;
wire _68_ ;
wire _141_ ;
wire _370_ ;
wire _426_ ;
wire _235_ ;
wire _464_ ;
wire _273_ ;
wire _329_ ;
wire _138_ ;
wire _30_ ;
wire _367_ ;
wire _176_ ;
wire _27_ ;
wire _100_ ;
wire _65_ ;
wire _423_ ;
wire _232_ ;
wire _461_ ;
wire _270_ ;
wire _326_ ;
wire _135_ ;
wire _364_ ;
wire CSR_Wen_traps ;
wire _114__bF$buf0 ;
wire _114__bF$buf1 ;
wire _114__bF$buf2 ;
wire _114__bF$buf3 ;
wire _114__bF$buf4 ;
wire _114__bF$buf5 ;
wire _114__bF$buf6 ;
wire _173_ ;
wire _229_ ;
wire _458_ ;
wire _267_ ;
wire _24_ ;
wire [31:0] CSR_mepc ;
wire _62_ ;
wire _399_ ;
wire _420_ ;
wire _323_ ;
wire _59_ ;
wire _132_ ;
wire _361_ ;
wire _417_ ;
wire _97_ ;
wire _170_ ;
wire _226_ ;
wire _455_ ;
wire _264_ ;
wire [11:0] CSR_addr ;
wire _129_ ;
wire [29:0] _21_ ;
wire _358_ ;
wire _167_ ;
wire _396_ ;
wire _299_ ;
wire _18_ ;
wire _320_ ;
wire _56_ ;
wire _414_ ;
wire _94_ ;
wire _223_ ;
wire _452_ ;
wire _261_ ;
wire _317_ ;
wire _126_ ;
wire _355_ ;
wire _164_ ;
wire _393_ ;
wire [31:0] CSR_PCaddr ;
wire _449_ ;
wire _258_ ;
wire [31:0] _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _199_ ;
wire _411_ ;
wire _91_ ;
wire _220_ ;
wire _9_ ;
wire _108__bF$buf0 ;
wire _108__bF$buf1 ;
wire _108__bF$buf2 ;
wire _108__bF$buf3 ;
wire _108__bF$buf4 ;
wire _314_ ;
wire _123_ ;
wire _352_ ;
wire _408_ ;
wire _88_ ;
wire _161_ ;
wire _217_ ;
wire _390_ ;
wire _446_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _349_ ;
wire _158_ ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _311_ ;
wire _47_ ;
wire _120_ ;
wire _405_ ;
wire _85_ ;
wire _214_ ;
wire _443_ ;
wire _252_ ;
wire CSR_Ret_bF$buf0 ;
wire CSR_Ret_bF$buf1 ;
wire CSR_Ret_bF$buf2 ;
wire CSR_Ret_bF$buf3 ;
wire CSR_Ret_bF$buf4 ;
wire CSR_Ret_bF$buf5 ;
wire _308_ ;
wire _481_ ;
wire _117_ ;
wire _290_ ;
wire _346_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _249_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _402_ ;
wire _82_ ;
wire _211_ ;
wire _440_ ;
wire _305_ ;
wire _114_ ;
wire _343_ ;
wire _79_ ;
wire _152_ ;
wire _208_ ;
wire _381_ ;
wire _437_ ;
wire _190_ ;
wire _246_ ;
wire _475_ ;
wire _284_ ;
wire _0_ ;
wire Extern_IRQ ;
wire _149_ ;
wire _41_ ;
wire _378_ ;
wire _187_ ;
wire _302_ ;
wire [3:0] CSR_mcause ;
wire _38_ ;
wire _111_ ;
wire _340_ ;
wire _76_ ;
wire _205_ ;
wire _434_ ;
wire _243_ ;
wire _472_ ;
wire _108_ ;
wire _281_ ;
wire _337_ ;
wire _146_ ;
wire _375_ ;
wire _184_ ;
wire _469_ ;
wire _278_ ;
wire _35_ ;
wire _73_ ;
wire _202_ ;
wire _431_ ;
wire _240_ ;
wire _105_ ;
wire _334_ ;
wire _143_ ;
wire _372_ ;
wire _428_ ;
wire _181_ ;
wire _237_ ;
wire _466_ ;
wire _275_ ;
wire [31:0] CSR_Wdata ;
wire _32_ ;
wire _369_ ;
wire _178_ ;
wire _70_ ;
wire _170__bF$buf0 ;
wire _170__bF$buf1 ;
wire _170__bF$buf2 ;
wire _170__bF$buf3 ;
wire _170__bF$buf4 ;
wire _170__bF$buf5 ;
wire _170__bF$buf6 ;
wire _29_ ;
wire _102_ ;
wire _331_ ;
wire _67_ ;
wire _140_ ;
wire _425_ ;
wire _234_ ;
wire _463_ ;
wire _272_ ;
wire _328_ ;
wire _137_ ;
wire _366_ ;
wire _175_ ;
wire _269_ ;
wire _26_ ;
wire _64_ ;
wire _422_ ;
wire _231_ ;
wire _460_ ;
wire _325_ ;
wire _134_ ;
wire _363_ ;
wire _419_ ;
wire _99_ ;
wire _172_ ;
wire _228_ ;
wire _457_ ;
wire [29:0] mepc ;
wire _266_ ;
wire _23_ ;
wire _169_ ;
wire _61_ ;
wire _398_ ;
wire meta_irq ;
wire _322_ ;
wire _58_ ;
wire _131_ ;
wire _360_ ;
wire _416_ ;
wire _96_ ;
wire _225_ ;
wire _454_ ;
wire _263_ ;
wire _319_ ;
wire _128_ ;
wire _20_ ;
wire _357_ ;
wire _166_ ;
wire _395_ ;
wire _298_ ;
wire _11__bF$buf0 ;
wire _11__bF$buf1 ;
wire _11__bF$buf2 ;
wire _11__bF$buf3 ;
wire _11__bF$buf4 ;
wire _17_ ;
wire _55_ ;
wire _413_ ;
wire _93_ ;
wire _222_ ;
wire _112__bF$buf0 ;
wire _112__bF$buf1 ;
wire _112__bF$buf2 ;
wire _112__bF$buf3 ;
wire _112__bF$buf4 ;
wire _112__bF$buf5 ;
wire _112__bF$buf6 ;
wire _451_ ;
wire _260_ ;
wire _316_ ;
wire _125_ ;
wire _354_ ;
wire _163_ ;
wire _219_ ;
wire _392_ ;
wire _448_ ;
wire _257_ ;
wire [31:0] _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _198_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _313_ ;
wire _49_ ;
wire _122_ ;
wire _351_ ;
wire _407_ ;
wire _87_ ;
wire _160_ ;
wire _216_ ;
wire CSR_Wen ;
wire _445_ ;
wire _254_ ;
wire _483_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _348_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire _289_ ;
wire _5_ ;
wire _310_ ;
wire _237__bF$buf0 ;
wire _237__bF$buf1 ;
wire _237__bF$buf2 ;
wire _237__bF$buf3 ;
wire _237__bF$buf4 ;
wire _46_ ;
wire _404_ ;
wire _84_ ;
wire _213_ ;
wire _442_ ;
wire _251_ ;
wire _307_ ;
wire _480_ ;
wire _116_ ;
wire _345_ ;
wire _154_ ;
wire _383_ ;
wire _439_ ;
wire _192_ ;
wire _248_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _24__bF$buf0 ;
wire _24__bF$buf1 ;
wire _24__bF$buf2 ;
wire _24__bF$buf3 ;
wire _24__bF$buf4 ;
wire _401_ ;
wire _81_ ;
wire _210_ ;
wire _304_ ;
wire _113_ ;
wire _342_ ;
wire _78_ ;
wire _151_ ;
wire _207_ ;
wire _380_ ;
wire _436_ ;
wire _245_ ;
wire _474_ ;
wire _283_ ;
wire _339_ ;
wire CSR_Wen_traps_bF$buf0 ;
wire CSR_Wen_traps_bF$buf1 ;
wire CSR_Wen_traps_bF$buf2 ;
wire CSR_Wen_traps_bF$buf3 ;
wire CSR_Wen_traps_bF$buf4 ;
wire CSR_Wen_traps_bF$buf5 ;
wire _148_ ;
wire _40_ ;
wire _377_ ;
wire _186_ ;
wire _31__bF$buf0 ;
wire _31__bF$buf1 ;
wire _31__bF$buf2 ;
wire _31__bF$buf3 ;
wire _31__bF$buf4 ;
wire _301_ ;
wire _37_ ;
wire _110_ ;
wire CSR_Ret ;
wire _75_ ;
wire _204_ ;
wire _433_ ;
wire _242_ ;
wire _471_ ;
wire _107_ ;
wire _280_ ;
wire _336_ ;
wire _145_ ;
wire _374_ ;
wire _183_ ;
wire _239_ ;
wire _468_ ;
wire _277_ ;
wire [31:0] mvect ;
wire _34_ ;
wire _72_ ;
wire _201_ ;
wire _430_ ;
wire _104_ ;
wire _333_ ;
wire _69_ ;
wire _142_ ;
wire _371_ ;
wire _427_ ;
wire _180_ ;
wire _236_ ;
wire _465_ ;
wire _274_ ;
wire _139_ ;
wire _31_ ;
wire _368_ ;
wire _177_ ;
wire [31:0] _28_ ;
wire _101_ ;
wire _330_ ;
wire _66_ ;
wire _424_ ;
wire _233_ ;
wire _462_ ;
wire _271_ ;
wire _327_ ;
wire _136_ ;
wire _365_ ;
wire _174_ ;
wire _459_ ;
wire _268_ ;
wire _25_ ;
wire _63_ ;
wire _421_ ;
wire _230_ ;
wire [31:0] CSR_data ;
wire [31:0] mcause ;
wire _324_ ;
wire _133_ ;
wire _362_ ;
wire _418_ ;
wire _98_ ;
wire _171_ ;
wire _227_ ;
wire _456_ ;
wire _265_ ;
wire mie ;
wire mip ;
wire _22_ ;
wire _359_ ;

BUFX2 BUFX2_insert71 (
    .A(_31_),
    .Y(_31__bF$buf0)
);

BUFX2 BUFX2_insert70 (
    .A(_31_),
    .Y(_31__bF$buf1)
);

BUFX2 BUFX2_insert69 (
    .A(_31_),
    .Y(_31__bF$buf2)
);

BUFX2 BUFX2_insert68 (
    .A(_31_),
    .Y(_31__bF$buf3)
);

BUFX2 BUFX2_insert67 (
    .A(_31_),
    .Y(_31__bF$buf4)
);

BUFX2 BUFX2_insert66 (
    .A(CSR_Ret),
    .Y(CSR_Ret_bF$buf0)
);

BUFX2 BUFX2_insert65 (
    .A(CSR_Ret),
    .Y(CSR_Ret_bF$buf1)
);

BUFX2 BUFX2_insert64 (
    .A(CSR_Ret),
    .Y(CSR_Ret_bF$buf2)
);

BUFX2 BUFX2_insert63 (
    .A(CSR_Ret),
    .Y(CSR_Ret_bF$buf3)
);

BUFX2 BUFX2_insert62 (
    .A(CSR_Ret),
    .Y(CSR_Ret_bF$buf4)
);

BUFX2 BUFX2_insert61 (
    .A(CSR_Ret),
    .Y(CSR_Ret_bF$buf5)
);

BUFX2 BUFX2_insert60 (
    .A(_11_),
    .Y(_11__bF$buf0)
);

BUFX2 BUFX2_insert59 (
    .A(_11_),
    .Y(_11__bF$buf1)
);

BUFX2 BUFX2_insert58 (
    .A(_11_),
    .Y(_11__bF$buf2)
);

BUFX2 BUFX2_insert57 (
    .A(_11_),
    .Y(_11__bF$buf3)
);

BUFX2 BUFX2_insert56 (
    .A(_11_),
    .Y(_11__bF$buf4)
);

BUFX2 BUFX2_insert55 (
    .A(_237_),
    .Y(_237__bF$buf0)
);

BUFX2 BUFX2_insert54 (
    .A(_237_),
    .Y(_237__bF$buf1)
);

BUFX2 BUFX2_insert53 (
    .A(_237_),
    .Y(_237__bF$buf2)
);

BUFX2 BUFX2_insert52 (
    .A(_237_),
    .Y(_237__bF$buf3)
);

BUFX2 BUFX2_insert51 (
    .A(_237_),
    .Y(_237__bF$buf4)
);

BUFX2 BUFX2_insert50 (
    .A(_108_),
    .Y(_108__bF$buf0)
);

BUFX2 BUFX2_insert49 (
    .A(_108_),
    .Y(_108__bF$buf1)
);

BUFX2 BUFX2_insert48 (
    .A(_108_),
    .Y(_108__bF$buf2)
);

BUFX2 BUFX2_insert47 (
    .A(_108_),
    .Y(_108__bF$buf3)
);

BUFX2 BUFX2_insert46 (
    .A(_108_),
    .Y(_108__bF$buf4)
);

BUFX2 BUFX2_insert45 (
    .A(_114_),
    .Y(_114__bF$buf0)
);

BUFX2 BUFX2_insert44 (
    .A(_114_),
    .Y(_114__bF$buf1)
);

BUFX2 BUFX2_insert43 (
    .A(_114_),
    .Y(_114__bF$buf2)
);

BUFX2 BUFX2_insert42 (
    .A(_114_),
    .Y(_114__bF$buf3)
);

BUFX2 BUFX2_insert41 (
    .A(_114_),
    .Y(_114__bF$buf4)
);

BUFX2 BUFX2_insert40 (
    .A(_114_),
    .Y(_114__bF$buf5)
);

BUFX2 BUFX2_insert39 (
    .A(_114_),
    .Y(_114__bF$buf6)
);

BUFX2 BUFX2_insert38 (
    .A(_170_),
    .Y(_170__bF$buf0)
);

BUFX2 BUFX2_insert37 (
    .A(_170_),
    .Y(_170__bF$buf1)
);

BUFX2 BUFX2_insert36 (
    .A(_170_),
    .Y(_170__bF$buf2)
);

BUFX2 BUFX2_insert35 (
    .A(_170_),
    .Y(_170__bF$buf3)
);

BUFX2 BUFX2_insert34 (
    .A(_170_),
    .Y(_170__bF$buf4)
);

BUFX2 BUFX2_insert33 (
    .A(_170_),
    .Y(_170__bF$buf5)
);

BUFX2 BUFX2_insert32 (
    .A(_170_),
    .Y(_170__bF$buf6)
);

BUFX2 BUFX2_insert31 (
    .A(_24_),
    .Y(_24__bF$buf0)
);

BUFX2 BUFX2_insert30 (
    .A(_24_),
    .Y(_24__bF$buf1)
);

BUFX2 BUFX2_insert29 (
    .A(_24_),
    .Y(_24__bF$buf2)
);

BUFX2 BUFX2_insert28 (
    .A(_24_),
    .Y(_24__bF$buf3)
);

BUFX2 BUFX2_insert27 (
    .A(_24_),
    .Y(_24__bF$buf4)
);

BUFX2 BUFX2_insert26 (
    .A(CSR_Wen_traps),
    .Y(CSR_Wen_traps_bF$buf0)
);

BUFX2 BUFX2_insert25 (
    .A(CSR_Wen_traps),
    .Y(CSR_Wen_traps_bF$buf1)
);

BUFX2 BUFX2_insert24 (
    .A(CSR_Wen_traps),
    .Y(CSR_Wen_traps_bF$buf2)
);

BUFX2 BUFX2_insert23 (
    .A(CSR_Wen_traps),
    .Y(CSR_Wen_traps_bF$buf3)
);

BUFX2 BUFX2_insert22 (
    .A(CSR_Wen_traps),
    .Y(CSR_Wen_traps_bF$buf4)
);

BUFX2 BUFX2_insert21 (
    .A(CSR_Wen_traps),
    .Y(CSR_Wen_traps_bF$buf5)
);

BUFX2 BUFX2_insert20 (
    .A(_235_),
    .Y(_235__bF$buf0)
);

BUFX2 BUFX2_insert19 (
    .A(_235_),
    .Y(_235__bF$buf1)
);

BUFX2 BUFX2_insert18 (
    .A(_235_),
    .Y(_235__bF$buf2)
);

BUFX2 BUFX2_insert17 (
    .A(_235_),
    .Y(_235__bF$buf3)
);

BUFX2 BUFX2_insert16 (
    .A(_235_),
    .Y(_235__bF$buf4)
);

CLKBUF1 CLKBUF1_insert15 (
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert14 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert13 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert12 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert11 (
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert10 (
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert9 (
    .A(clk),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert8 (
    .A(clk),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert7 (
    .A(clk),
    .Y(clk_bF$buf8)
);

BUFX2 BUFX2_insert6 (
    .A(_112_),
    .Y(_112__bF$buf0)
);

BUFX2 BUFX2_insert5 (
    .A(_112_),
    .Y(_112__bF$buf1)
);

BUFX2 BUFX2_insert4 (
    .A(_112_),
    .Y(_112__bF$buf2)
);

BUFX2 BUFX2_insert3 (
    .A(_112_),
    .Y(_112__bF$buf3)
);

BUFX2 BUFX2_insert2 (
    .A(_112_),
    .Y(_112__bF$buf4)
);

BUFX2 BUFX2_insert1 (
    .A(_112_),
    .Y(_112__bF$buf5)
);

BUFX2 BUFX2_insert0 (
    .A(_112_),
    .Y(_112__bF$buf6)
);

NAND2X1 _1000_ (
    .A(mepc[11]),
    .B(CSR_Ret_bF$buf5),
    .Y(_375_)
);

OAI21X1 _1001_ (
    .A(_372_),
    .B(_192_),
    .C(_194_),
    .Y(_376_)
);

INVX1 _1002_ (
    .A(_376_),
    .Y(_377_)
);

NAND2X1 _1003_ (
    .A(mvect[12]),
    .B(mvect[13]),
    .Y(_378_)
);

OAI21X1 _1004_ (
    .A(_372_),
    .B(_378_),
    .C(_108__bF$buf4),
    .Y(_379_)
);

OAI21X1 _1005_ (
    .A(_377_),
    .B(_379_),
    .C(_375_),
    .Y(_486_[13])
);

NAND2X1 _1006_ (
    .A(mepc[12]),
    .B(CSR_Ret_bF$buf4),
    .Y(_380_)
);

OAI21X1 _1007_ (
    .A(_372_),
    .B(_378_),
    .C(_196_),
    .Y(_381_)
);

INVX1 _1008_ (
    .A(_381_),
    .Y(_382_)
);

OR2X2 _1009_ (
    .A(_372_),
    .B(_378_),
    .Y(_383_)
);

OAI21X1 _1010_ (
    .A(_383_),
    .B(_196_),
    .C(_108__bF$buf3),
    .Y(_384_)
);

OAI21X1 _1011_ (
    .A(_384_),
    .B(_382_),
    .C(_380_),
    .Y(_486_[14])
);

NAND2X1 _1012_ (
    .A(mepc[13]),
    .B(CSR_Ret_bF$buf3),
    .Y(_385_)
);

OAI21X1 _1013_ (
    .A(_383_),
    .B(_196_),
    .C(_198_),
    .Y(_386_)
);

INVX1 _1014_ (
    .A(_386_),
    .Y(_387_)
);

NAND2X1 _1015_ (
    .A(mvect[14]),
    .B(mvect[15]),
    .Y(_388_)
);

OR2X2 _1016_ (
    .A(_378_),
    .B(_388_),
    .Y(_389_)
);

OAI21X1 _1017_ (
    .A(_372_),
    .B(_389_),
    .C(_108__bF$buf2),
    .Y(_390_)
);

OAI21X1 _1018_ (
    .A(_387_),
    .B(_390_),
    .C(_385_),
    .Y(_486_[15])
);

NAND2X1 _1019_ (
    .A(mepc[14]),
    .B(CSR_Ret_bF$buf2),
    .Y(_391_)
);

NOR2X1 _1020_ (
    .A(_389_),
    .B(_372_),
    .Y(_392_)
);

NOR2X1 _1021_ (
    .A(_378_),
    .B(_388_),
    .Y(_393_)
);

NAND3X1 _1022_ (
    .A(_371_),
    .B(_393_),
    .C(_350_),
    .Y(_394_)
);

NOR2X1 _1023_ (
    .A(_328_),
    .B(_394_),
    .Y(_395_)
);

NAND2X1 _1024_ (
    .A(mvect[16]),
    .B(_395_),
    .Y(_396_)
);

OAI21X1 _1025_ (
    .A(mvect[16]),
    .B(_392_),
    .C(_396_),
    .Y(_397_)
);

OAI21X1 _1026_ (
    .A(_397_),
    .B(CSR_Ret_bF$buf1),
    .C(_391_),
    .Y(_486_[16])
);

NAND2X1 _1027_ (
    .A(mepc[15]),
    .B(CSR_Ret_bF$buf0),
    .Y(_398_)
);

AOI21X1 _1028_ (
    .A(mvect[16]),
    .B(_395_),
    .C(mvect[17]),
    .Y(_399_)
);

INVX2 _1029_ (
    .A(_392_),
    .Y(_400_)
);

NAND2X1 _1030_ (
    .A(mvect[16]),
    .B(mvect[17]),
    .Y(_401_)
);

OAI21X1 _1031_ (
    .A(_400_),
    .B(_401_),
    .C(_108__bF$buf1),
    .Y(_402_)
);

OAI21X1 _1032_ (
    .A(_402_),
    .B(_399_),
    .C(_398_),
    .Y(_486_[17])
);

NAND2X1 _1033_ (
    .A(mepc[16]),
    .B(CSR_Ret_bF$buf5),
    .Y(_403_)
);

AND2X2 _1034_ (
    .A(mvect[16]),
    .B(mvect[17]),
    .Y(_404_)
);

AOI21X1 _1035_ (
    .A(_404_),
    .B(_392_),
    .C(mvect[18]),
    .Y(_405_)
);

NAND2X1 _1036_ (
    .A(mvect[18]),
    .B(_404_),
    .Y(_406_)
);

OAI21X1 _1037_ (
    .A(_400_),
    .B(_406_),
    .C(_108__bF$buf0),
    .Y(_407_)
);

OAI21X1 _1038_ (
    .A(_407_),
    .B(_405_),
    .C(_403_),
    .Y(_486_[18])
);

NAND2X1 _1039_ (
    .A(mepc[17]),
    .B(CSR_Ret_bF$buf4),
    .Y(_408_)
);

INVX1 _1040_ (
    .A(_406_),
    .Y(_409_)
);

AOI21X1 _1041_ (
    .A(_409_),
    .B(_395_),
    .C(mvect[19]),
    .Y(_410_)
);

AND2X2 _1042_ (
    .A(mvect[18]),
    .B(mvect[19]),
    .Y(_411_)
);

NAND2X1 _1043_ (
    .A(_404_),
    .B(_411_),
    .Y(_412_)
);

OAI21X1 _1044_ (
    .A(_400_),
    .B(_412_),
    .C(_108__bF$buf4),
    .Y(_413_)
);

OAI21X1 _1045_ (
    .A(_413_),
    .B(_410_),
    .C(_408_),
    .Y(_486_[19])
);

NAND2X1 _1046_ (
    .A(mepc[18]),
    .B(CSR_Ret_bF$buf3),
    .Y(_414_)
);

NAND3X1 _1047_ (
    .A(_404_),
    .B(_411_),
    .C(_392_),
    .Y(_415_)
);

AND2X2 _1048_ (
    .A(_415_),
    .B(_208_),
    .Y(_416_)
);

OAI21X1 _1049_ (
    .A(_415_),
    .B(_208_),
    .C(_108__bF$buf3),
    .Y(_417_)
);

OAI21X1 _1050_ (
    .A(_416_),
    .B(_417_),
    .C(_414_),
    .Y(_486_[20])
);

NAND2X1 _1051_ (
    .A(mepc[19]),
    .B(CSR_Ret_bF$buf2),
    .Y(_418_)
);

NOR2X1 _1052_ (
    .A(_208_),
    .B(_412_),
    .Y(_419_)
);

AOI21X1 _1053_ (
    .A(_419_),
    .B(_395_),
    .C(mvect[21]),
    .Y(_420_)
);

AND2X2 _1054_ (
    .A(mvect[20]),
    .B(mvect[21]),
    .Y(_421_)
);

NAND3X1 _1055_ (
    .A(_404_),
    .B(_411_),
    .C(_421_),
    .Y(_422_)
);

OAI21X1 _1056_ (
    .A(_400_),
    .B(_422_),
    .C(_108__bF$buf2),
    .Y(_423_)
);

OAI21X1 _1057_ (
    .A(_423_),
    .B(_420_),
    .C(_418_),
    .Y(_486_[21])
);

NAND2X1 _1058_ (
    .A(mepc[20]),
    .B(CSR_Ret_bF$buf1),
    .Y(_424_)
);

NAND2X1 _1059_ (
    .A(mvect[18]),
    .B(mvect[19]),
    .Y(_425_)
);

NAND2X1 _1060_ (
    .A(mvect[20]),
    .B(mvect[21]),
    .Y(_426_)
);

NOR3X1 _1061_ (
    .A(_401_),
    .B(_425_),
    .C(_426_),
    .Y(_427_)
);

NAND3X1 _1062_ (
    .A(_371_),
    .B(_393_),
    .C(_427_),
    .Y(_428_)
);

NOR2X1 _1063_ (
    .A(_356_),
    .B(_428_),
    .Y(_429_)
);

NOR2X1 _1064_ (
    .A(mvect[22]),
    .B(_429_),
    .Y(_430_)
);

NAND2X1 _1065_ (
    .A(mvect[22]),
    .B(_429_),
    .Y(_431_)
);

NAND2X1 _1066_ (
    .A(_108__bF$buf1),
    .B(_431_),
    .Y(_432_)
);

OAI21X1 _1067_ (
    .A(_432_),
    .B(_430_),
    .C(_424_),
    .Y(_486_[22])
);

NOR2X1 _1068_ (
    .A(mepc[21]),
    .B(_108__bF$buf0),
    .Y(_433_)
);

OR2X2 _1069_ (
    .A(_431_),
    .B(mvect[23]),
    .Y(_434_)
);

AOI21X1 _1070_ (
    .A(mvect[23]),
    .B(_431_),
    .C(CSR_Ret_bF$buf0),
    .Y(_435_)
);

AOI21X1 _1071_ (
    .A(_435_),
    .B(_434_),
    .C(_433_),
    .Y(_486_[23])
);

NAND2X1 _1072_ (
    .A(mepc[22]),
    .B(CSR_Ret_bF$buf5),
    .Y(_436_)
);

NAND2X1 _1073_ (
    .A(mvect[22]),
    .B(mvect[23]),
    .Y(_437_)
);

NOR3X1 _1074_ (
    .A(_356_),
    .B(_437_),
    .C(_428_),
    .Y(_438_)
);

NOR2X1 _1075_ (
    .A(mvect[24]),
    .B(_438_),
    .Y(_439_)
);

INVX1 _1076_ (
    .A(_438_),
    .Y(_440_)
);

OAI21X1 _1077_ (
    .A(_440_),
    .B(_216_),
    .C(_108__bF$buf4),
    .Y(_441_)
);

OAI21X1 _1078_ (
    .A(_441_),
    .B(_439_),
    .C(_436_),
    .Y(_486_[24])
);

NAND2X1 _1079_ (
    .A(mepc[23]),
    .B(CSR_Ret_bF$buf4),
    .Y(_442_)
);

AOI21X1 _1080_ (
    .A(mvect[24]),
    .B(_438_),
    .C(mvect[25]),
    .Y(_443_)
);

NAND2X1 _1081_ (
    .A(mvect[24]),
    .B(mvect[25]),
    .Y(_444_)
);

OAI21X1 _1082_ (
    .A(_440_),
    .B(_444_),
    .C(_108__bF$buf3),
    .Y(_445_)
);

OAI21X1 _1083_ (
    .A(_445_),
    .B(_443_),
    .C(_442_),
    .Y(_486_[25])
);

INVX1 _1084_ (
    .A(_444_),
    .Y(_446_)
);

AOI21X1 _1085_ (
    .A(_446_),
    .B(_438_),
    .C(mvect[26]),
    .Y(_447_)
);

NAND3X1 _1086_ (
    .A(mvect[26]),
    .B(_446_),
    .C(_438_),
    .Y(_448_)
);

NAND2X1 _1087_ (
    .A(_108__bF$buf2),
    .B(_448_),
    .Y(_449_)
);

NAND2X1 _1088_ (
    .A(mepc[24]),
    .B(CSR_Ret_bF$buf3),
    .Y(_450_)
);

OAI21X1 _1089_ (
    .A(_449_),
    .B(_447_),
    .C(_450_),
    .Y(_486_[26])
);

NAND3X1 _1090_ (
    .A(_222_),
    .B(_108__bF$buf1),
    .C(_448_),
    .Y(_451_)
);

NOR2X1 _1091_ (
    .A(mepc[25]),
    .B(_108__bF$buf0),
    .Y(_452_)
);

NAND2X1 _1092_ (
    .A(mvect[26]),
    .B(mvect[27]),
    .Y(_453_)
);

NOR2X1 _1093_ (
    .A(_444_),
    .B(_453_),
    .Y(_454_)
);

AND2X2 _1094_ (
    .A(_454_),
    .B(_108__bF$buf4),
    .Y(_455_)
);

AOI21X1 _1095_ (
    .A(_455_),
    .B(_438_),
    .C(_452_),
    .Y(_456_)
);

AND2X2 _1096_ (
    .A(_451_),
    .B(_456_),
    .Y(_486_[27])
);

NAND2X1 _1097_ (
    .A(mepc[26]),
    .B(CSR_Ret_bF$buf2),
    .Y(_457_)
);

NOR3X1 _1098_ (
    .A(_437_),
    .B(_444_),
    .C(_453_),
    .Y(_458_)
);

INVX1 _1099_ (
    .A(_458_),
    .Y(_459_)
);

NOR3X1 _1100_ (
    .A(_356_),
    .B(_459_),
    .C(_428_),
    .Y(_460_)
);

NOR2X1 _1101_ (
    .A(mvect[28]),
    .B(_460_),
    .Y(_461_)
);

NOR3X1 _1102_ (
    .A(_368_),
    .B(_389_),
    .C(_422_),
    .Y(_462_)
);

NAND3X1 _1103_ (
    .A(_351_),
    .B(_458_),
    .C(_462_),
    .Y(_463_)
);

OAI21X1 _1104_ (
    .A(_463_),
    .B(_224_),
    .C(_108__bF$buf3),
    .Y(_464_)
);

OAI21X1 _1105_ (
    .A(_464_),
    .B(_461_),
    .C(_457_),
    .Y(_486_[28])
);

NOR2X1 _1106_ (
    .A(mepc[27]),
    .B(_108__bF$buf2),
    .Y(_465_)
);

NAND2X1 _1107_ (
    .A(mvect[28]),
    .B(_460_),
    .Y(_466_)
);

OR2X2 _1108_ (
    .A(_466_),
    .B(mvect[29]),
    .Y(_467_)
);

AOI21X1 _1109_ (
    .A(mvect[29]),
    .B(_466_),
    .C(CSR_Ret_bF$buf1),
    .Y(_468_)
);

AOI21X1 _1110_ (
    .A(_468_),
    .B(_467_),
    .C(_465_),
    .Y(_486_[29])
);

INVX1 _1111_ (
    .A(mepc[28]),
    .Y(_469_)
);

NAND2X1 _1112_ (
    .A(mvect[28]),
    .B(mvect[29]),
    .Y(_470_)
);

NOR3X1 _1113_ (
    .A(_0_),
    .B(_470_),
    .C(_157_),
    .Y(_471_)
);

NAND3X1 _1114_ (
    .A(_350_),
    .B(_458_),
    .C(_471_),
    .Y(_472_)
);

OAI21X1 _1115_ (
    .A(_472_),
    .B(_428_),
    .C(mvect[30]),
    .Y(_473_)
);

INVX1 _1116_ (
    .A(_473_),
    .Y(_474_)
);

NOR2X1 _1117_ (
    .A(_428_),
    .B(_472_),
    .Y(_475_)
);

AND2X2 _1118_ (
    .A(_475_),
    .B(_228_),
    .Y(_476_)
);

OAI21X1 _1119_ (
    .A(_476_),
    .B(_474_),
    .C(_108__bF$buf1),
    .Y(_477_)
);

OAI21X1 _1120_ (
    .A(_469_),
    .B(_108__bF$buf0),
    .C(_477_),
    .Y(_486_[30])
);

INVX1 _1121_ (
    .A(_470_),
    .Y(_478_)
);

NAND2X1 _1122_ (
    .A(mvect[30]),
    .B(_478_),
    .Y(_479_)
);

INVX1 _1123_ (
    .A(_479_),
    .Y(_480_)
);

AOI21X1 _1124_ (
    .A(_480_),
    .B(_460_),
    .C(_230_),
    .Y(_481_)
);

NOR3X1 _1125_ (
    .A(mvect[31]),
    .B(_479_),
    .C(_463_),
    .Y(_482_)
);

OAI21X1 _1126_ (
    .A(_482_),
    .B(_481_),
    .C(_108__bF$buf4),
    .Y(_483_)
);

NAND2X1 _1127_ (
    .A(mepc[29]),
    .B(CSR_Ret_bF$buf0),
    .Y(_484_)
);

NAND2X1 _1128_ (
    .A(_484_),
    .B(_483_),
    .Y(_486_[31])
);

BUFX2 _1129_ (
    .A(_485_),
    .Y(CSR_IRQ)
);

BUFX2 _1130_ (
    .A(1'h0),
    .Y(CSR_PCaddr[0])
);

BUFX2 _1131_ (
    .A(1'h0),
    .Y(CSR_PCaddr[1])
);

BUFX2 _1132_ (
    .A(_486_[2]),
    .Y(CSR_PCaddr[2])
);

BUFX2 _1133_ (
    .A(_486_[3]),
    .Y(CSR_PCaddr[3])
);

BUFX2 _1134_ (
    .A(_486_[4]),
    .Y(CSR_PCaddr[4])
);

BUFX2 _1135_ (
    .A(_486_[5]),
    .Y(CSR_PCaddr[5])
);

BUFX2 _1136_ (
    .A(_486_[6]),
    .Y(CSR_PCaddr[6])
);

BUFX2 _1137_ (
    .A(_486_[7]),
    .Y(CSR_PCaddr[7])
);

BUFX2 _1138_ (
    .A(_486_[8]),
    .Y(CSR_PCaddr[8])
);

BUFX2 _1139_ (
    .A(_486_[9]),
    .Y(CSR_PCaddr[9])
);

BUFX2 _1140_ (
    .A(_486_[10]),
    .Y(CSR_PCaddr[10])
);

BUFX2 _1141_ (
    .A(_486_[11]),
    .Y(CSR_PCaddr[11])
);

BUFX2 _1142_ (
    .A(_486_[12]),
    .Y(CSR_PCaddr[12])
);

BUFX2 _1143_ (
    .A(_486_[13]),
    .Y(CSR_PCaddr[13])
);

BUFX2 _1144_ (
    .A(_486_[14]),
    .Y(CSR_PCaddr[14])
);

BUFX2 _1145_ (
    .A(_486_[15]),
    .Y(CSR_PCaddr[15])
);

BUFX2 _1146_ (
    .A(_486_[16]),
    .Y(CSR_PCaddr[16])
);

BUFX2 _1147_ (
    .A(_486_[17]),
    .Y(CSR_PCaddr[17])
);

BUFX2 _1148_ (
    .A(_486_[18]),
    .Y(CSR_PCaddr[18])
);

BUFX2 _1149_ (
    .A(_486_[19]),
    .Y(CSR_PCaddr[19])
);

BUFX2 _1150_ (
    .A(_486_[20]),
    .Y(CSR_PCaddr[20])
);

BUFX2 _1151_ (
    .A(_486_[21]),
    .Y(CSR_PCaddr[21])
);

BUFX2 _1152_ (
    .A(_486_[22]),
    .Y(CSR_PCaddr[22])
);

BUFX2 _1153_ (
    .A(_486_[23]),
    .Y(CSR_PCaddr[23])
);

BUFX2 _1154_ (
    .A(_486_[24]),
    .Y(CSR_PCaddr[24])
);

BUFX2 _1155_ (
    .A(_486_[25]),
    .Y(CSR_PCaddr[25])
);

BUFX2 _1156_ (
    .A(_486_[26]),
    .Y(CSR_PCaddr[26])
);

BUFX2 _1157_ (
    .A(_486_[27]),
    .Y(CSR_PCaddr[27])
);

BUFX2 _1158_ (
    .A(_486_[28]),
    .Y(CSR_PCaddr[28])
);

BUFX2 _1159_ (
    .A(_486_[29]),
    .Y(CSR_PCaddr[29])
);

BUFX2 _1160_ (
    .A(_486_[30]),
    .Y(CSR_PCaddr[30])
);

BUFX2 _1161_ (
    .A(_486_[31]),
    .Y(CSR_PCaddr[31])
);

BUFX2 _1162_ (
    .A(_487_[0]),
    .Y(CSR_data[0])
);

BUFX2 _1163_ (
    .A(_487_[1]),
    .Y(CSR_data[1])
);

BUFX2 _1164_ (
    .A(_487_[2]),
    .Y(CSR_data[2])
);

BUFX2 _1165_ (
    .A(_487_[3]),
    .Y(CSR_data[3])
);

BUFX2 _1166_ (
    .A(_487_[4]),
    .Y(CSR_data[4])
);

BUFX2 _1167_ (
    .A(_487_[5]),
    .Y(CSR_data[5])
);

BUFX2 _1168_ (
    .A(_487_[6]),
    .Y(CSR_data[6])
);

BUFX2 _1169_ (
    .A(_487_[7]),
    .Y(CSR_data[7])
);

BUFX2 _1170_ (
    .A(_487_[8]),
    .Y(CSR_data[8])
);

BUFX2 _1171_ (
    .A(_487_[9]),
    .Y(CSR_data[9])
);

BUFX2 _1172_ (
    .A(_487_[10]),
    .Y(CSR_data[10])
);

BUFX2 _1173_ (
    .A(_487_[11]),
    .Y(CSR_data[11])
);

BUFX2 _1174_ (
    .A(_487_[12]),
    .Y(CSR_data[12])
);

BUFX2 _1175_ (
    .A(_487_[13]),
    .Y(CSR_data[13])
);

BUFX2 _1176_ (
    .A(_487_[14]),
    .Y(CSR_data[14])
);

BUFX2 _1177_ (
    .A(_487_[15]),
    .Y(CSR_data[15])
);

BUFX2 _1178_ (
    .A(_487_[16]),
    .Y(CSR_data[16])
);

BUFX2 _1179_ (
    .A(_487_[17]),
    .Y(CSR_data[17])
);

BUFX2 _1180_ (
    .A(_487_[18]),
    .Y(CSR_data[18])
);

BUFX2 _1181_ (
    .A(_487_[19]),
    .Y(CSR_data[19])
);

BUFX2 _1182_ (
    .A(_487_[20]),
    .Y(CSR_data[20])
);

BUFX2 _1183_ (
    .A(_487_[21]),
    .Y(CSR_data[21])
);

BUFX2 _1184_ (
    .A(_487_[22]),
    .Y(CSR_data[22])
);

BUFX2 _1185_ (
    .A(_487_[23]),
    .Y(CSR_data[23])
);

BUFX2 _1186_ (
    .A(_487_[24]),
    .Y(CSR_data[24])
);

BUFX2 _1187_ (
    .A(_487_[25]),
    .Y(CSR_data[25])
);

BUFX2 _1188_ (
    .A(_487_[26]),
    .Y(CSR_data[26])
);

BUFX2 _1189_ (
    .A(_487_[27]),
    .Y(CSR_data[27])
);

BUFX2 _1190_ (
    .A(_487_[28]),
    .Y(CSR_data[28])
);

BUFX2 _1191_ (
    .A(_487_[29]),
    .Y(CSR_data[29])
);

BUFX2 _1192_ (
    .A(_487_[30]),
    .Y(CSR_data[30])
);

BUFX2 _1193_ (
    .A(_487_[31]),
    .Y(CSR_data[31])
);

DFFPOSX1 _1194_ (
    .CLK(clk_bF$buf8),
    .D(_21_[0]),
    .Q(mepc[0])
);

DFFPOSX1 _1195_ (
    .CLK(clk_bF$buf7),
    .D(_21_[1]),
    .Q(mepc[1])
);

DFFPOSX1 _1196_ (
    .CLK(clk_bF$buf6),
    .D(_21_[2]),
    .Q(mepc[2])
);

DFFPOSX1 _1197_ (
    .CLK(clk_bF$buf5),
    .D(_21_[3]),
    .Q(mepc[3])
);

DFFPOSX1 _1198_ (
    .CLK(clk_bF$buf4),
    .D(_21_[4]),
    .Q(mepc[4])
);

DFFPOSX1 _1199_ (
    .CLK(clk_bF$buf3),
    .D(_21_[5]),
    .Q(mepc[5])
);

DFFPOSX1 _1200_ (
    .CLK(clk_bF$buf2),
    .D(_21_[6]),
    .Q(mepc[6])
);

DFFPOSX1 _1201_ (
    .CLK(clk_bF$buf1),
    .D(_21_[7]),
    .Q(mepc[7])
);

DFFPOSX1 _1202_ (
    .CLK(clk_bF$buf0),
    .D(_21_[8]),
    .Q(mepc[8])
);

DFFPOSX1 _1203_ (
    .CLK(clk_bF$buf8),
    .D(_21_[9]),
    .Q(mepc[9])
);

DFFPOSX1 _1204_ (
    .CLK(clk_bF$buf7),
    .D(_21_[10]),
    .Q(mepc[10])
);

DFFPOSX1 _1205_ (
    .CLK(clk_bF$buf6),
    .D(_21_[11]),
    .Q(mepc[11])
);

DFFPOSX1 _1206_ (
    .CLK(clk_bF$buf5),
    .D(_21_[12]),
    .Q(mepc[12])
);

DFFPOSX1 _1207_ (
    .CLK(clk_bF$buf4),
    .D(_21_[13]),
    .Q(mepc[13])
);

DFFPOSX1 _1208_ (
    .CLK(clk_bF$buf3),
    .D(_21_[14]),
    .Q(mepc[14])
);

DFFPOSX1 _1209_ (
    .CLK(clk_bF$buf2),
    .D(_21_[15]),
    .Q(mepc[15])
);

DFFPOSX1 _1210_ (
    .CLK(clk_bF$buf1),
    .D(_21_[16]),
    .Q(mepc[16])
);

DFFPOSX1 _1211_ (
    .CLK(clk_bF$buf0),
    .D(_21_[17]),
    .Q(mepc[17])
);

DFFPOSX1 _1212_ (
    .CLK(clk_bF$buf8),
    .D(_21_[18]),
    .Q(mepc[18])
);

DFFPOSX1 _1213_ (
    .CLK(clk_bF$buf7),
    .D(_21_[19]),
    .Q(mepc[19])
);

DFFPOSX1 _1214_ (
    .CLK(clk_bF$buf6),
    .D(_21_[20]),
    .Q(mepc[20])
);

DFFPOSX1 _1215_ (
    .CLK(clk_bF$buf5),
    .D(_21_[21]),
    .Q(mepc[21])
);

DFFPOSX1 _1216_ (
    .CLK(clk_bF$buf4),
    .D(_21_[22]),
    .Q(mepc[22])
);

DFFPOSX1 _1217_ (
    .CLK(clk_bF$buf3),
    .D(_21_[23]),
    .Q(mepc[23])
);

DFFPOSX1 _1218_ (
    .CLK(clk_bF$buf2),
    .D(_21_[24]),
    .Q(mepc[24])
);

DFFPOSX1 _1219_ (
    .CLK(clk_bF$buf1),
    .D(_21_[25]),
    .Q(mepc[25])
);

DFFPOSX1 _1220_ (
    .CLK(clk_bF$buf0),
    .D(_21_[26]),
    .Q(mepc[26])
);

DFFPOSX1 _1221_ (
    .CLK(clk_bF$buf8),
    .D(_21_[27]),
    .Q(mepc[27])
);

DFFPOSX1 _1222_ (
    .CLK(clk_bF$buf7),
    .D(_21_[28]),
    .Q(mepc[28])
);

DFFPOSX1 _1223_ (
    .CLK(clk_bF$buf6),
    .D(_21_[29]),
    .Q(mepc[29])
);

DFFPOSX1 _1224_ (
    .CLK(clk_bF$buf5),
    .D(Extern_IRQ),
    .Q(meta_irq)
);

DFFPOSX1 _1225_ (
    .CLK(clk_bF$buf4),
    .D(meta_irq),
    .Q(mip)
);

DFFPOSX1 _1226_ (
    .CLK(clk_bF$buf3),
    .D(_14_),
    .Q(mie)
);

DFFPOSX1 _1227_ (
    .CLK(clk_bF$buf2),
    .D(_07_[0]),
    .Q(mvect[0])
);

DFFPOSX1 _1228_ (
    .CLK(clk_bF$buf1),
    .D(_07_[1]),
    .Q(mvect[1])
);

DFFPOSX1 _1229_ (
    .CLK(clk_bF$buf0),
    .D(_07_[2]),
    .Q(mvect[2])
);

DFFPOSX1 _1230_ (
    .CLK(clk_bF$buf8),
    .D(_07_[3]),
    .Q(mvect[3])
);

DFFPOSX1 _1231_ (
    .CLK(clk_bF$buf7),
    .D(_07_[4]),
    .Q(mvect[4])
);

DFFPOSX1 _1232_ (
    .CLK(clk_bF$buf6),
    .D(_07_[5]),
    .Q(mvect[5])
);

DFFPOSX1 _1233_ (
    .CLK(clk_bF$buf5),
    .D(_07_[6]),
    .Q(mvect[6])
);

DFFPOSX1 _1234_ (
    .CLK(clk_bF$buf4),
    .D(_07_[7]),
    .Q(mvect[7])
);

DFFPOSX1 _1235_ (
    .CLK(clk_bF$buf3),
    .D(_07_[8]),
    .Q(mvect[8])
);

DFFPOSX1 _1236_ (
    .CLK(clk_bF$buf2),
    .D(_07_[9]),
    .Q(mvect[9])
);

DFFPOSX1 _1237_ (
    .CLK(clk_bF$buf1),
    .D(_07_[10]),
    .Q(mvect[10])
);

DFFPOSX1 _1238_ (
    .CLK(clk_bF$buf0),
    .D(_07_[11]),
    .Q(mvect[11])
);

DFFPOSX1 _1239_ (
    .CLK(clk_bF$buf8),
    .D(_07_[12]),
    .Q(mvect[12])
);

DFFPOSX1 _1240_ (
    .CLK(clk_bF$buf7),
    .D(_07_[13]),
    .Q(mvect[13])
);

DFFPOSX1 _1241_ (
    .CLK(clk_bF$buf6),
    .D(_07_[14]),
    .Q(mvect[14])
);

DFFPOSX1 _1242_ (
    .CLK(clk_bF$buf5),
    .D(_07_[15]),
    .Q(mvect[15])
);

DFFPOSX1 _1243_ (
    .CLK(clk_bF$buf4),
    .D(_07_[16]),
    .Q(mvect[16])
);

DFFPOSX1 _1244_ (
    .CLK(clk_bF$buf3),
    .D(_07_[17]),
    .Q(mvect[17])
);

DFFPOSX1 _1245_ (
    .CLK(clk_bF$buf2),
    .D(_07_[18]),
    .Q(mvect[18])
);

DFFPOSX1 _1246_ (
    .CLK(clk_bF$buf1),
    .D(_07_[19]),
    .Q(mvect[19])
);

DFFPOSX1 _1247_ (
    .CLK(clk_bF$buf0),
    .D(_07_[20]),
    .Q(mvect[20])
);

DFFPOSX1 _1248_ (
    .CLK(clk_bF$buf8),
    .D(_07_[21]),
    .Q(mvect[21])
);

DFFPOSX1 _1249_ (
    .CLK(clk_bF$buf7),
    .D(_07_[22]),
    .Q(mvect[22])
);

DFFPOSX1 _1250_ (
    .CLK(clk_bF$buf6),
    .D(_07_[23]),
    .Q(mvect[23])
);

DFFPOSX1 _1251_ (
    .CLK(clk_bF$buf5),
    .D(_07_[24]),
    .Q(mvect[24])
);

DFFPOSX1 _1252_ (
    .CLK(clk_bF$buf4),
    .D(_07_[25]),
    .Q(mvect[25])
);

DFFPOSX1 _1253_ (
    .CLK(clk_bF$buf3),
    .D(_07_[26]),
    .Q(mvect[26])
);

DFFPOSX1 _1254_ (
    .CLK(clk_bF$buf2),
    .D(_07_[27]),
    .Q(mvect[27])
);

DFFPOSX1 _1255_ (
    .CLK(clk_bF$buf1),
    .D(_07_[28]),
    .Q(mvect[28])
);

DFFPOSX1 _1256_ (
    .CLK(clk_bF$buf0),
    .D(_07_[29]),
    .Q(mvect[29])
);

DFFPOSX1 _1257_ (
    .CLK(clk_bF$buf8),
    .D(_07_[30]),
    .Q(mvect[30])
);

DFFPOSX1 _1258_ (
    .CLK(clk_bF$buf7),
    .D(_07_[31]),
    .Q(mvect[31])
);

DFFPOSX1 _1259_ (
    .CLK(clk_bF$buf6),
    .D(_33_[0]),
    .Q(mstatus[0])
);

DFFPOSX1 _1260_ (
    .CLK(clk_bF$buf5),
    .D(_33_[1]),
    .Q(mstatus[1])
);

DFFPOSX1 _1261_ (
    .CLK(clk_bF$buf4),
    .D(_28_[0]),
    .Q(mcause[0])
);

DFFPOSX1 _1262_ (
    .CLK(clk_bF$buf3),
    .D(_28_[1]),
    .Q(mcause[1])
);

DFFPOSX1 _1263_ (
    .CLK(clk_bF$buf2),
    .D(_28_[2]),
    .Q(mcause[2])
);

DFFPOSX1 _1264_ (
    .CLK(clk_bF$buf1),
    .D(_28_[3]),
    .Q(mcause[3])
);

DFFPOSX1 _1265_ (
    .CLK(clk_bF$buf0),
    .D(_28_[4]),
    .Q(mcause[4])
);

DFFPOSX1 _1266_ (
    .CLK(clk_bF$buf8),
    .D(_28_[5]),
    .Q(mcause[5])
);

DFFPOSX1 _1267_ (
    .CLK(clk_bF$buf7),
    .D(_28_[6]),
    .Q(mcause[6])
);

DFFPOSX1 _1268_ (
    .CLK(clk_bF$buf6),
    .D(_28_[7]),
    .Q(mcause[7])
);

DFFPOSX1 _1269_ (
    .CLK(clk_bF$buf5),
    .D(_28_[8]),
    .Q(mcause[8])
);

DFFPOSX1 _1270_ (
    .CLK(clk_bF$buf4),
    .D(_28_[9]),
    .Q(mcause[9])
);

DFFPOSX1 _1271_ (
    .CLK(clk_bF$buf3),
    .D(_28_[10]),
    .Q(mcause[10])
);

DFFPOSX1 _1272_ (
    .CLK(clk_bF$buf2),
    .D(_28_[11]),
    .Q(mcause[11])
);

DFFPOSX1 _1273_ (
    .CLK(clk_bF$buf1),
    .D(_28_[12]),
    .Q(mcause[12])
);

DFFPOSX1 _1274_ (
    .CLK(clk_bF$buf0),
    .D(_28_[13]),
    .Q(mcause[13])
);

DFFPOSX1 _1275_ (
    .CLK(clk_bF$buf8),
    .D(_28_[14]),
    .Q(mcause[14])
);

DFFPOSX1 _1276_ (
    .CLK(clk_bF$buf7),
    .D(_28_[15]),
    .Q(mcause[15])
);

DFFPOSX1 _1277_ (
    .CLK(clk_bF$buf6),
    .D(_28_[16]),
    .Q(mcause[16])
);

DFFPOSX1 _1278_ (
    .CLK(clk_bF$buf5),
    .D(_28_[17]),
    .Q(mcause[17])
);

DFFPOSX1 _1279_ (
    .CLK(clk_bF$buf4),
    .D(_28_[18]),
    .Q(mcause[18])
);

DFFPOSX1 _1280_ (
    .CLK(clk_bF$buf3),
    .D(_28_[19]),
    .Q(mcause[19])
);

DFFPOSX1 _1281_ (
    .CLK(clk_bF$buf2),
    .D(_28_[20]),
    .Q(mcause[20])
);

DFFPOSX1 _1282_ (
    .CLK(clk_bF$buf1),
    .D(_28_[21]),
    .Q(mcause[21])
);

DFFPOSX1 _1283_ (
    .CLK(clk_bF$buf0),
    .D(_28_[22]),
    .Q(mcause[22])
);

DFFPOSX1 _1284_ (
    .CLK(clk_bF$buf8),
    .D(_28_[23]),
    .Q(mcause[23])
);

DFFPOSX1 _1285_ (
    .CLK(clk_bF$buf7),
    .D(_28_[24]),
    .Q(mcause[24])
);

DFFPOSX1 _1286_ (
    .CLK(clk_bF$buf6),
    .D(_28_[25]),
    .Q(mcause[25])
);

DFFPOSX1 _1287_ (
    .CLK(clk_bF$buf5),
    .D(_28_[26]),
    .Q(mcause[26])
);

DFFPOSX1 _1288_ (
    .CLK(clk_bF$buf4),
    .D(_28_[27]),
    .Q(mcause[27])
);

DFFPOSX1 _1289_ (
    .CLK(clk_bF$buf3),
    .D(_28_[28]),
    .Q(mcause[28])
);

DFFPOSX1 _1290_ (
    .CLK(clk_bF$buf2),
    .D(_28_[29]),
    .Q(mcause[29])
);

DFFPOSX1 _1291_ (
    .CLK(clk_bF$buf1),
    .D(_28_[30]),
    .Q(mcause[30])
);

DFFPOSX1 _1292_ (
    .CLK(clk_bF$buf0),
    .D(_28_[31]),
    .Q(mcause[31])
);

INVX2 _488_ (
    .A(mvect[0]),
    .Y(_0_)
);

NOR2X1 _489_ (
    .A(CSR_addr[11]),
    .B(CSR_addr[10]),
    .Y(_1_)
);

NAND3X1 _490_ (
    .A(CSR_addr[9]),
    .B(CSR_addr[8]),
    .C(_1_),
    .Y(_2_)
);

INVX1 _491_ (
    .A(CSR_addr[7]),
    .Y(_3_)
);

NOR2X1 _492_ (
    .A(CSR_addr[5]),
    .B(CSR_addr[4]),
    .Y(_4_)
);

NAND3X1 _493_ (
    .A(_3_),
    .B(CSR_addr[6]),
    .C(_4_),
    .Y(_5_)
);

NOR2X1 _494_ (
    .A(_2_),
    .B(_5_),
    .Y(_6_)
);

OR2X2 _495_ (
    .A(CSR_addr[3]),
    .B(CSR_addr[2]),
    .Y(_7_)
);

INVX1 _496_ (
    .A(CSR_addr[0]),
    .Y(_8_)
);

NAND2X1 _497_ (
    .A(CSR_addr[1]),
    .B(_8_),
    .Y(_9_)
);

NOR2X1 _498_ (
    .A(_7_),
    .B(_9_),
    .Y(_10_)
);

NAND2X1 _499_ (
    .A(_10_),
    .B(_6_),
    .Y(_11_)
);

INVX4 _500_ (
    .A(_11__bF$buf4),
    .Y(_12_)
);

NAND2X1 _501_ (
    .A(mcause[0]),
    .B(_12_),
    .Y(_13_)
);

NOR2X1 _502_ (
    .A(CSR_addr[7]),
    .B(CSR_addr[6]),
    .Y(_15_)
);

NAND2X1 _503_ (
    .A(_4_),
    .B(_15_),
    .Y(_16_)
);

NOR2X1 _504_ (
    .A(_16_),
    .B(_2_),
    .Y(_17_)
);

INVX1 _505_ (
    .A(CSR_addr[1]),
    .Y(_18_)
);

NAND2X1 _506_ (
    .A(CSR_addr[0]),
    .B(_18_),
    .Y(_19_)
);

INVX1 _507_ (
    .A(CSR_addr[3]),
    .Y(_20_)
);

NAND2X1 _508_ (
    .A(CSR_addr[2]),
    .B(_20_),
    .Y(_22_)
);

NOR2X1 _509_ (
    .A(_19_),
    .B(_22_),
    .Y(_23_)
);

AND2X2 _510_ (
    .A(_17_),
    .B(_23_),
    .Y(_24_)
);

INVX1 _511_ (
    .A(_24__bF$buf4),
    .Y(_25_)
);

OAI21X1 _512_ (
    .A(_0_),
    .B(_25_),
    .C(_13_),
    .Y(_487_[0])
);

INVX1 _513_ (
    .A(mvect[1]),
    .Y(_26_)
);

NAND2X1 _514_ (
    .A(mcause[1]),
    .B(_12_),
    .Y(_27_)
);

OAI21X1 _515_ (
    .A(_26_),
    .B(_25_),
    .C(_27_),
    .Y(_487_[1])
);

INVX1 _516_ (
    .A(mcause[2]),
    .Y(_29_)
);

NOR2X1 _517_ (
    .A(_7_),
    .B(_19_),
    .Y(_30_)
);

AND2X2 _518_ (
    .A(_6_),
    .B(_30_),
    .Y(_31_)
);

AOI22X1 _519_ (
    .A(_24__bF$buf3),
    .B(mvect[2]),
    .C(mepc[0]),
    .D(_31__bF$buf4),
    .Y(_32_)
);

OAI21X1 _520_ (
    .A(_29_),
    .B(_11__bF$buf3),
    .C(_32_),
    .Y(_487_[2])
);

INVX1 _521_ (
    .A(mstatus[0]),
    .Y(_34_)
);

NOR2X1 _522_ (
    .A(CSR_addr[1]),
    .B(CSR_addr[0]),
    .Y(_35_)
);

INVX1 _523_ (
    .A(_17_),
    .Y(_36_)
);

NOR2X1 _524_ (
    .A(_7_),
    .B(_36_),
    .Y(_37_)
);

NAND2X1 _525_ (
    .A(_35_),
    .B(_37_),
    .Y(_38_)
);

NAND2X1 _526_ (
    .A(mepc[1]),
    .B(_31__bF$buf3),
    .Y(_39_)
);

AOI22X1 _527_ (
    .A(mvect[3]),
    .B(_24__bF$buf2),
    .C(_12_),
    .D(mcause[3]),
    .Y(_40_)
);

AND2X2 _528_ (
    .A(_40_),
    .B(_39_),
    .Y(_41_)
);

OAI21X1 _529_ (
    .A(_34_),
    .B(_38_),
    .C(_41_),
    .Y(_487_[3])
);

INVX1 _530_ (
    .A(mcause[4]),
    .Y(_42_)
);

AOI22X1 _531_ (
    .A(_24__bF$buf1),
    .B(mvect[4]),
    .C(mepc[2]),
    .D(_31__bF$buf2),
    .Y(_43_)
);

OAI21X1 _532_ (
    .A(_42_),
    .B(_11__bF$buf2),
    .C(_43_),
    .Y(_487_[4])
);

INVX1 _533_ (
    .A(mcause[5]),
    .Y(_44_)
);

AOI22X1 _534_ (
    .A(_24__bF$buf0),
    .B(mvect[5]),
    .C(mepc[3]),
    .D(_31__bF$buf1),
    .Y(_45_)
);

OAI21X1 _535_ (
    .A(_44_),
    .B(_11__bF$buf1),
    .C(_45_),
    .Y(_487_[5])
);

INVX1 _536_ (
    .A(mcause[6]),
    .Y(_46_)
);

AOI22X1 _537_ (
    .A(_24__bF$buf4),
    .B(mvect[6]),
    .C(mepc[4]),
    .D(_31__bF$buf0),
    .Y(_47_)
);

OAI21X1 _538_ (
    .A(_46_),
    .B(_11__bF$buf0),
    .C(_47_),
    .Y(_487_[6])
);

INVX1 _539_ (
    .A(mstatus[1]),
    .Y(_48_)
);

NAND2X1 _540_ (
    .A(mepc[5]),
    .B(_31__bF$buf4),
    .Y(_49_)
);

AOI22X1 _541_ (
    .A(mvect[7]),
    .B(_24__bF$buf3),
    .C(_12_),
    .D(mcause[7]),
    .Y(_50_)
);

AND2X2 _542_ (
    .A(_50_),
    .B(_49_),
    .Y(_51_)
);

OAI21X1 _543_ (
    .A(_48_),
    .B(_38_),
    .C(_51_),
    .Y(_487_[7])
);

AND2X2 _544_ (
    .A(_17_),
    .B(_30_),
    .Y(_52_)
);

AOI21X1 _545_ (
    .A(mvect[8]),
    .B(_24__bF$buf2),
    .C(_52_),
    .Y(_53_)
);

AOI22X1 _546_ (
    .A(mepc[6]),
    .B(_31__bF$buf3),
    .C(_12_),
    .D(mcause[8]),
    .Y(_54_)
);

NAND2X1 _547_ (
    .A(_53_),
    .B(_54_),
    .Y(_487_[8])
);

INVX1 _548_ (
    .A(mcause[9]),
    .Y(_55_)
);

AOI22X1 _549_ (
    .A(_24__bF$buf1),
    .B(mvect[9]),
    .C(mepc[7]),
    .D(_31__bF$buf2),
    .Y(_56_)
);

OAI21X1 _550_ (
    .A(_55_),
    .B(_11__bF$buf4),
    .C(_56_),
    .Y(_487_[9])
);

INVX1 _551_ (
    .A(mcause[10]),
    .Y(_57_)
);

AOI22X1 _552_ (
    .A(_24__bF$buf0),
    .B(mvect[10]),
    .C(mepc[8]),
    .D(_31__bF$buf1),
    .Y(_58_)
);

OAI21X1 _553_ (
    .A(_57_),
    .B(_11__bF$buf3),
    .C(_58_),
    .Y(_487_[10])
);

INVX1 _554_ (
    .A(mip),
    .Y(_59_)
);

INVX1 _555_ (
    .A(_35_),
    .Y(_60_)
);

OR2X2 _556_ (
    .A(_60_),
    .B(_22_),
    .Y(_61_)
);

NOR2X1 _557_ (
    .A(_59_),
    .B(_61_),
    .Y(_62_)
);

AOI22X1 _558_ (
    .A(_6_),
    .B(_62_),
    .C(_37_),
    .D(_35_),
    .Y(_63_)
);

NOR2X1 _559_ (
    .A(_61_),
    .B(_36_),
    .Y(_64_)
);

AOI22X1 _560_ (
    .A(mcause[11]),
    .B(_12_),
    .C(_64_),
    .D(mie),
    .Y(_65_)
);

AOI22X1 _561_ (
    .A(_24__bF$buf4),
    .B(mvect[11]),
    .C(mepc[9]),
    .D(_31__bF$buf0),
    .Y(_66_)
);

NAND3X1 _562_ (
    .A(_66_),
    .B(_63_),
    .C(_65_),
    .Y(_487_[11])
);

NAND2X1 _563_ (
    .A(mepc[10]),
    .B(_31__bF$buf4),
    .Y(_67_)
);

AOI22X1 _564_ (
    .A(mvect[12]),
    .B(_24__bF$buf3),
    .C(_12_),
    .D(mcause[12]),
    .Y(_68_)
);

NAND3X1 _565_ (
    .A(_38_),
    .B(_67_),
    .C(_68_),
    .Y(_487_[12])
);

INVX1 _566_ (
    .A(mcause[13]),
    .Y(_69_)
);

AOI22X1 _567_ (
    .A(_24__bF$buf2),
    .B(mvect[13]),
    .C(mepc[11]),
    .D(_31__bF$buf3),
    .Y(_70_)
);

OAI21X1 _568_ (
    .A(_69_),
    .B(_11__bF$buf2),
    .C(_70_),
    .Y(_487_[13])
);

INVX1 _569_ (
    .A(mcause[14]),
    .Y(_71_)
);

AOI22X1 _570_ (
    .A(_24__bF$buf1),
    .B(mvect[14]),
    .C(mepc[12]),
    .D(_31__bF$buf2),
    .Y(_72_)
);

OAI21X1 _571_ (
    .A(_71_),
    .B(_11__bF$buf1),
    .C(_72_),
    .Y(_487_[14])
);

INVX1 _572_ (
    .A(mcause[15]),
    .Y(_73_)
);

AOI22X1 _573_ (
    .A(_24__bF$buf0),
    .B(mvect[15]),
    .C(mepc[13]),
    .D(_31__bF$buf1),
    .Y(_74_)
);

OAI21X1 _574_ (
    .A(_73_),
    .B(_11__bF$buf0),
    .C(_74_),
    .Y(_487_[15])
);

INVX1 _575_ (
    .A(mcause[16]),
    .Y(_75_)
);

AOI22X1 _576_ (
    .A(_24__bF$buf4),
    .B(mvect[16]),
    .C(mepc[14]),
    .D(_31__bF$buf0),
    .Y(_76_)
);

OAI21X1 _577_ (
    .A(_75_),
    .B(_11__bF$buf4),
    .C(_76_),
    .Y(_487_[16])
);

INVX1 _578_ (
    .A(mcause[17]),
    .Y(_77_)
);

AOI22X1 _579_ (
    .A(_24__bF$buf3),
    .B(mvect[17]),
    .C(mepc[15]),
    .D(_31__bF$buf4),
    .Y(_78_)
);

OAI21X1 _580_ (
    .A(_77_),
    .B(_11__bF$buf3),
    .C(_78_),
    .Y(_487_[17])
);

INVX1 _581_ (
    .A(mcause[18]),
    .Y(_79_)
);

AOI22X1 _582_ (
    .A(_24__bF$buf2),
    .B(mvect[18]),
    .C(mepc[16]),
    .D(_31__bF$buf3),
    .Y(_80_)
);

OAI21X1 _583_ (
    .A(_79_),
    .B(_11__bF$buf2),
    .C(_80_),
    .Y(_487_[18])
);

INVX1 _584_ (
    .A(mcause[19]),
    .Y(_81_)
);

AOI22X1 _585_ (
    .A(_24__bF$buf1),
    .B(mvect[19]),
    .C(mepc[17]),
    .D(_31__bF$buf2),
    .Y(_82_)
);

OAI21X1 _586_ (
    .A(_81_),
    .B(_11__bF$buf1),
    .C(_82_),
    .Y(_487_[19])
);

INVX1 _587_ (
    .A(mcause[20]),
    .Y(_83_)
);

AOI22X1 _588_ (
    .A(_24__bF$buf0),
    .B(mvect[20]),
    .C(mepc[18]),
    .D(_31__bF$buf1),
    .Y(_84_)
);

OAI21X1 _589_ (
    .A(_83_),
    .B(_11__bF$buf0),
    .C(_84_),
    .Y(_487_[20])
);

INVX1 _590_ (
    .A(mcause[21]),
    .Y(_85_)
);

AOI22X1 _591_ (
    .A(_24__bF$buf4),
    .B(mvect[21]),
    .C(mepc[19]),
    .D(_31__bF$buf0),
    .Y(_86_)
);

OAI21X1 _592_ (
    .A(_85_),
    .B(_11__bF$buf4),
    .C(_86_),
    .Y(_487_[21])
);

INVX1 _593_ (
    .A(mcause[22]),
    .Y(_87_)
);

AOI22X1 _594_ (
    .A(_24__bF$buf3),
    .B(mvect[22]),
    .C(mepc[20]),
    .D(_31__bF$buf4),
    .Y(_88_)
);

OAI21X1 _595_ (
    .A(_87_),
    .B(_11__bF$buf3),
    .C(_88_),
    .Y(_487_[22])
);

INVX1 _596_ (
    .A(mcause[23]),
    .Y(_89_)
);

AOI22X1 _597_ (
    .A(_24__bF$buf2),
    .B(mvect[23]),
    .C(mepc[21]),
    .D(_31__bF$buf3),
    .Y(_90_)
);

OAI21X1 _598_ (
    .A(_89_),
    .B(_11__bF$buf2),
    .C(_90_),
    .Y(_487_[23])
);

INVX1 _599_ (
    .A(mcause[24]),
    .Y(_91_)
);

AOI22X1 _600_ (
    .A(_24__bF$buf1),
    .B(mvect[24]),
    .C(mepc[22]),
    .D(_31__bF$buf2),
    .Y(_92_)
);

OAI21X1 _601_ (
    .A(_91_),
    .B(_11__bF$buf1),
    .C(_92_),
    .Y(_487_[24])
);

INVX1 _602_ (
    .A(mcause[25]),
    .Y(_93_)
);

AOI22X1 _603_ (
    .A(_24__bF$buf0),
    .B(mvect[25]),
    .C(mepc[23]),
    .D(_31__bF$buf1),
    .Y(_94_)
);

OAI21X1 _604_ (
    .A(_93_),
    .B(_11__bF$buf0),
    .C(_94_),
    .Y(_487_[25])
);

INVX1 _605_ (
    .A(mcause[26]),
    .Y(_95_)
);

AOI22X1 _606_ (
    .A(_24__bF$buf4),
    .B(mvect[26]),
    .C(mepc[24]),
    .D(_31__bF$buf0),
    .Y(_96_)
);

OAI21X1 _607_ (
    .A(_95_),
    .B(_11__bF$buf4),
    .C(_96_),
    .Y(_487_[26])
);

INVX1 _608_ (
    .A(mcause[27]),
    .Y(_97_)
);

AOI22X1 _609_ (
    .A(_24__bF$buf3),
    .B(mvect[27]),
    .C(mepc[25]),
    .D(_31__bF$buf4),
    .Y(_98_)
);

OAI21X1 _610_ (
    .A(_97_),
    .B(_11__bF$buf3),
    .C(_98_),
    .Y(_487_[27])
);

INVX1 _611_ (
    .A(mcause[28]),
    .Y(_99_)
);

AOI22X1 _612_ (
    .A(_24__bF$buf2),
    .B(mvect[28]),
    .C(mepc[26]),
    .D(_31__bF$buf3),
    .Y(_100_)
);

OAI21X1 _613_ (
    .A(_99_),
    .B(_11__bF$buf2),
    .C(_100_),
    .Y(_487_[28])
);

INVX1 _614_ (
    .A(mcause[29]),
    .Y(_101_)
);

AOI22X1 _615_ (
    .A(_24__bF$buf1),
    .B(mvect[29]),
    .C(mepc[27]),
    .D(_31__bF$buf2),
    .Y(_102_)
);

OAI21X1 _616_ (
    .A(_101_),
    .B(_11__bF$buf1),
    .C(_102_),
    .Y(_487_[29])
);

AOI21X1 _617_ (
    .A(mvect[30]),
    .B(_24__bF$buf0),
    .C(_52_),
    .Y(_103_)
);

AOI22X1 _618_ (
    .A(mepc[28]),
    .B(_31__bF$buf1),
    .C(_12_),
    .D(mcause[30]),
    .Y(_104_)
);

NAND2X1 _619_ (
    .A(_103_),
    .B(_104_),
    .Y(_487_[30])
);

INVX1 _620_ (
    .A(mcause[31]),
    .Y(_105_)
);

AOI22X1 _621_ (
    .A(_24__bF$buf4),
    .B(mvect[31]),
    .C(mepc[29]),
    .D(_31__bF$buf0),
    .Y(_106_)
);

OAI21X1 _622_ (
    .A(_105_),
    .B(_11__bF$buf0),
    .C(_106_),
    .Y(_487_[31])
);

NAND2X1 _623_ (
    .A(CSR_mcause[0]),
    .B(CSR_Wen_traps_bF$buf5),
    .Y(_107_)
);

INVX8 _624_ (
    .A(CSR_Ret_bF$buf5),
    .Y(_108_)
);

NAND2X1 _625_ (
    .A(CSR_Wen),
    .B(_108__bF$buf3),
    .Y(_109_)
);

NOR2X1 _626_ (
    .A(_109_),
    .B(_11__bF$buf4),
    .Y(_110_)
);

NOR2X1 _627_ (
    .A(mcause[0]),
    .B(_110_),
    .Y(_111_)
);

INVX8 _628_ (
    .A(CSR_Wen_traps_bF$buf4),
    .Y(_112_)
);

INVX1 _629_ (
    .A(_109_),
    .Y(_113_)
);

NAND2X1 _630_ (
    .A(_113_),
    .B(_12_),
    .Y(_114_)
);

OAI21X1 _631_ (
    .A(_114__bF$buf6),
    .B(CSR_Wdata[0]),
    .C(_112__bF$buf6),
    .Y(_115_)
);

OAI21X1 _632_ (
    .A(_115_),
    .B(_111_),
    .C(_107_),
    .Y(_28_[0])
);

NAND2X1 _633_ (
    .A(CSR_Wen_traps_bF$buf3),
    .B(CSR_mcause[1]),
    .Y(_116_)
);

NOR2X1 _634_ (
    .A(mcause[1]),
    .B(_110_),
    .Y(_117_)
);

OAI21X1 _635_ (
    .A(_114__bF$buf5),
    .B(CSR_Wdata[1]),
    .C(_112__bF$buf5),
    .Y(_118_)
);

OAI21X1 _636_ (
    .A(_118_),
    .B(_117_),
    .C(_116_),
    .Y(_28_[1])
);

NAND2X1 _637_ (
    .A(CSR_Wen_traps_bF$buf2),
    .B(CSR_mcause[2]),
    .Y(_119_)
);

OAI21X1 _638_ (
    .A(_11__bF$buf3),
    .B(_109_),
    .C(_29_),
    .Y(_120_)
);

OAI21X1 _639_ (
    .A(_114__bF$buf4),
    .B(CSR_Wdata[2]),
    .C(_120_),
    .Y(_121_)
);

OAI21X1 _640_ (
    .A(_121_),
    .B(CSR_Wen_traps_bF$buf1),
    .C(_119_),
    .Y(_28_[2])
);

NAND2X1 _641_ (
    .A(CSR_Wen_traps_bF$buf0),
    .B(CSR_mcause[3]),
    .Y(_122_)
);

NOR2X1 _642_ (
    .A(mcause[3]),
    .B(_110_),
    .Y(_123_)
);

OAI21X1 _643_ (
    .A(_114__bF$buf3),
    .B(CSR_Wdata[3]),
    .C(_112__bF$buf4),
    .Y(_124_)
);

OAI21X1 _644_ (
    .A(_124_),
    .B(_123_),
    .C(_122_),
    .Y(_28_[3])
);

OAI21X1 _645_ (
    .A(_114__bF$buf2),
    .B(CSR_Wdata[4]),
    .C(_112__bF$buf3),
    .Y(_125_)
);

AOI21X1 _646_ (
    .A(_42_),
    .B(_114__bF$buf1),
    .C(_125_),
    .Y(_28_[4])
);

OAI21X1 _647_ (
    .A(_114__bF$buf0),
    .B(CSR_Wdata[5]),
    .C(_112__bF$buf2),
    .Y(_126_)
);

AOI21X1 _648_ (
    .A(_44_),
    .B(_114__bF$buf6),
    .C(_126_),
    .Y(_28_[5])
);

OAI21X1 _649_ (
    .A(_114__bF$buf5),
    .B(CSR_Wdata[6]),
    .C(_112__bF$buf1),
    .Y(_127_)
);

AOI21X1 _650_ (
    .A(_46_),
    .B(_114__bF$buf4),
    .C(_127_),
    .Y(_28_[6])
);

NOR2X1 _651_ (
    .A(mcause[7]),
    .B(_110_),
    .Y(_128_)
);

OAI21X1 _652_ (
    .A(_114__bF$buf3),
    .B(CSR_Wdata[7]),
    .C(_112__bF$buf0),
    .Y(_129_)
);

NOR2X1 _653_ (
    .A(_128_),
    .B(_129_),
    .Y(_28_[7])
);

NOR2X1 _654_ (
    .A(mcause[8]),
    .B(_110_),
    .Y(_130_)
);

OAI21X1 _655_ (
    .A(_114__bF$buf2),
    .B(CSR_Wdata[8]),
    .C(_112__bF$buf6),
    .Y(_131_)
);

NOR2X1 _656_ (
    .A(_130_),
    .B(_131_),
    .Y(_28_[8])
);

OAI21X1 _657_ (
    .A(_114__bF$buf1),
    .B(CSR_Wdata[9]),
    .C(_112__bF$buf5),
    .Y(_132_)
);

AOI21X1 _658_ (
    .A(_55_),
    .B(_114__bF$buf0),
    .C(_132_),
    .Y(_28_[9])
);

OAI21X1 _659_ (
    .A(_114__bF$buf6),
    .B(CSR_Wdata[10]),
    .C(_112__bF$buf4),
    .Y(_133_)
);

AOI21X1 _660_ (
    .A(_57_),
    .B(_114__bF$buf5),
    .C(_133_),
    .Y(_28_[10])
);

NOR2X1 _661_ (
    .A(mcause[11]),
    .B(_110_),
    .Y(_134_)
);

OAI21X1 _662_ (
    .A(_114__bF$buf4),
    .B(CSR_Wdata[11]),
    .C(_112__bF$buf3),
    .Y(_135_)
);

NOR2X1 _663_ (
    .A(_134_),
    .B(_135_),
    .Y(_28_[11])
);

NOR2X1 _664_ (
    .A(mcause[12]),
    .B(_110_),
    .Y(_136_)
);

OAI21X1 _665_ (
    .A(_114__bF$buf3),
    .B(CSR_Wdata[12]),
    .C(_112__bF$buf2),
    .Y(_137_)
);

NOR2X1 _666_ (
    .A(_136_),
    .B(_137_),
    .Y(_28_[12])
);

OAI21X1 _667_ (
    .A(_114__bF$buf2),
    .B(CSR_Wdata[13]),
    .C(_112__bF$buf1),
    .Y(_138_)
);

AOI21X1 _668_ (
    .A(_69_),
    .B(_114__bF$buf1),
    .C(_138_),
    .Y(_28_[13])
);

OAI21X1 _669_ (
    .A(_114__bF$buf0),
    .B(CSR_Wdata[14]),
    .C(_112__bF$buf0),
    .Y(_139_)
);

AOI21X1 _670_ (
    .A(_71_),
    .B(_114__bF$buf6),
    .C(_139_),
    .Y(_28_[14])
);

OAI21X1 _671_ (
    .A(_114__bF$buf5),
    .B(CSR_Wdata[15]),
    .C(_112__bF$buf6),
    .Y(_140_)
);

AOI21X1 _672_ (
    .A(_73_),
    .B(_114__bF$buf4),
    .C(_140_),
    .Y(_28_[15])
);

OAI21X1 _673_ (
    .A(_114__bF$buf3),
    .B(CSR_Wdata[16]),
    .C(_112__bF$buf5),
    .Y(_141_)
);

AOI21X1 _674_ (
    .A(_75_),
    .B(_114__bF$buf2),
    .C(_141_),
    .Y(_28_[16])
);

OAI21X1 _675_ (
    .A(_114__bF$buf1),
    .B(CSR_Wdata[17]),
    .C(_112__bF$buf4),
    .Y(_142_)
);

AOI21X1 _676_ (
    .A(_77_),
    .B(_114__bF$buf0),
    .C(_142_),
    .Y(_28_[17])
);

OAI21X1 _677_ (
    .A(_114__bF$buf6),
    .B(CSR_Wdata[18]),
    .C(_112__bF$buf3),
    .Y(_143_)
);

AOI21X1 _678_ (
    .A(_79_),
    .B(_114__bF$buf5),
    .C(_143_),
    .Y(_28_[18])
);

OAI21X1 _679_ (
    .A(_114__bF$buf4),
    .B(CSR_Wdata[19]),
    .C(_112__bF$buf2),
    .Y(_144_)
);

AOI21X1 _680_ (
    .A(_81_),
    .B(_114__bF$buf3),
    .C(_144_),
    .Y(_28_[19])
);

OAI21X1 _681_ (
    .A(_114__bF$buf2),
    .B(CSR_Wdata[20]),
    .C(_112__bF$buf1),
    .Y(_145_)
);

AOI21X1 _682_ (
    .A(_83_),
    .B(_114__bF$buf1),
    .C(_145_),
    .Y(_28_[20])
);

OAI21X1 _683_ (
    .A(_114__bF$buf0),
    .B(CSR_Wdata[21]),
    .C(_112__bF$buf0),
    .Y(_146_)
);

AOI21X1 _684_ (
    .A(_85_),
    .B(_114__bF$buf6),
    .C(_146_),
    .Y(_28_[21])
);

OAI21X1 _685_ (
    .A(_114__bF$buf5),
    .B(CSR_Wdata[22]),
    .C(_112__bF$buf6),
    .Y(_147_)
);

AOI21X1 _686_ (
    .A(_87_),
    .B(_114__bF$buf4),
    .C(_147_),
    .Y(_28_[22])
);

OAI21X1 _687_ (
    .A(_114__bF$buf3),
    .B(CSR_Wdata[23]),
    .C(_112__bF$buf5),
    .Y(_148_)
);

AOI21X1 _688_ (
    .A(_89_),
    .B(_114__bF$buf2),
    .C(_148_),
    .Y(_28_[23])
);

OAI21X1 _689_ (
    .A(_114__bF$buf1),
    .B(CSR_Wdata[24]),
    .C(_112__bF$buf4),
    .Y(_149_)
);

AOI21X1 _690_ (
    .A(_91_),
    .B(_114__bF$buf0),
    .C(_149_),
    .Y(_28_[24])
);

OAI21X1 _691_ (
    .A(_114__bF$buf6),
    .B(CSR_Wdata[25]),
    .C(_112__bF$buf3),
    .Y(_150_)
);

AOI21X1 _692_ (
    .A(_93_),
    .B(_114__bF$buf5),
    .C(_150_),
    .Y(_28_[25])
);

OAI21X1 _693_ (
    .A(_114__bF$buf4),
    .B(CSR_Wdata[26]),
    .C(_112__bF$buf2),
    .Y(_151_)
);

AOI21X1 _694_ (
    .A(_95_),
    .B(_114__bF$buf3),
    .C(_151_),
    .Y(_28_[26])
);

OAI21X1 _695_ (
    .A(_114__bF$buf2),
    .B(CSR_Wdata[27]),
    .C(_112__bF$buf1),
    .Y(_152_)
);

AOI21X1 _696_ (
    .A(_97_),
    .B(_114__bF$buf1),
    .C(_152_),
    .Y(_28_[27])
);

OAI21X1 _697_ (
    .A(_114__bF$buf0),
    .B(CSR_Wdata[28]),
    .C(_112__bF$buf0),
    .Y(_153_)
);

AOI21X1 _698_ (
    .A(_99_),
    .B(_114__bF$buf6),
    .C(_153_),
    .Y(_28_[28])
);

OAI21X1 _699_ (
    .A(_114__bF$buf5),
    .B(CSR_Wdata[29]),
    .C(_112__bF$buf6),
    .Y(_154_)
);

AOI21X1 _700_ (
    .A(_101_),
    .B(_114__bF$buf4),
    .C(_154_),
    .Y(_28_[29])
);

NOR2X1 _701_ (
    .A(mcause[30]),
    .B(_110_),
    .Y(_155_)
);

OAI21X1 _702_ (
    .A(_114__bF$buf3),
    .B(CSR_Wdata[30]),
    .C(_112__bF$buf5),
    .Y(_156_)
);

NOR2X1 _703_ (
    .A(_155_),
    .B(_156_),
    .Y(_28_[30])
);

NAND3X1 _704_ (
    .A(mstatus[0]),
    .B(mie),
    .C(mip),
    .Y(_157_)
);

INVX1 _705_ (
    .A(_157_),
    .Y(_485_)
);

NAND2X1 _706_ (
    .A(mcause[31]),
    .B(_112__bF$buf4),
    .Y(_158_)
);

OAI22X1 _707_ (
    .A(_112__bF$buf3),
    .B(_157_),
    .C(_110_),
    .D(_158_),
    .Y(_28_[31])
);

INVX1 _708_ (
    .A(CSR_Wen),
    .Y(_159_)
);

NOR2X1 _709_ (
    .A(_7_),
    .B(_60_),
    .Y(_160_)
);

NAND2X1 _710_ (
    .A(_160_),
    .B(_17_),
    .Y(_161_)
);

NOR2X1 _711_ (
    .A(_159_),
    .B(_161_),
    .Y(_162_)
);

INVX1 _712_ (
    .A(CSR_Wdata[3]),
    .Y(_163_)
);

NAND2X1 _713_ (
    .A(_163_),
    .B(_162_),
    .Y(_164_)
);

OAI21X1 _714_ (
    .A(mstatus[0]),
    .B(_162_),
    .C(_164_),
    .Y(_165_)
);

OAI21X1 _715_ (
    .A(_108__bF$buf2),
    .B(mstatus[1]),
    .C(_112__bF$buf2),
    .Y(_166_)
);

AOI21X1 _716_ (
    .A(_108__bF$buf1),
    .B(_165_),
    .C(_166_),
    .Y(_33_[0])
);

MUX2X1 _717_ (
    .A(CSR_Wdata[7]),
    .B(mstatus[1]),
    .S(_162_),
    .Y(_167_)
);

NOR2X1 _718_ (
    .A(CSR_Ret_bF$buf4),
    .B(CSR_Wen_traps_bF$buf5),
    .Y(_168_)
);

AOI22X1 _719_ (
    .A(_34_),
    .B(CSR_Wen_traps_bF$buf4),
    .C(_167_),
    .D(_168_),
    .Y(_33_[1])
);

NOR2X1 _720_ (
    .A(CSR_Wen_traps_bF$buf3),
    .B(_109_),
    .Y(_169_)
);

NAND2X1 _721_ (
    .A(_169_),
    .B(_24__bF$buf3),
    .Y(_170_)
);

NOR2X1 _722_ (
    .A(CSR_Wdata[0]),
    .B(_170__bF$buf6),
    .Y(_171_)
);

AOI21X1 _723_ (
    .A(_0_),
    .B(_170__bF$buf5),
    .C(_171_),
    .Y(_07_[0])
);

NOR2X1 _724_ (
    .A(CSR_Wdata[1]),
    .B(_170__bF$buf4),
    .Y(_172_)
);

AOI21X1 _725_ (
    .A(_26_),
    .B(_170__bF$buf3),
    .C(_172_),
    .Y(_07_[1])
);

INVX1 _726_ (
    .A(mvect[2]),
    .Y(_173_)
);

NOR2X1 _727_ (
    .A(CSR_Wdata[2]),
    .B(_170__bF$buf2),
    .Y(_174_)
);

AOI21X1 _728_ (
    .A(_173_),
    .B(_170__bF$buf1),
    .C(_174_),
    .Y(_07_[2])
);

INVX2 _729_ (
    .A(mvect[3]),
    .Y(_175_)
);

MUX2X1 _730_ (
    .A(_175_),
    .B(_163_),
    .S(_170__bF$buf0),
    .Y(_07_[3])
);

INVX2 _731_ (
    .A(mvect[4]),
    .Y(_176_)
);

NOR2X1 _732_ (
    .A(CSR_Wdata[4]),
    .B(_170__bF$buf6),
    .Y(_177_)
);

AOI21X1 _733_ (
    .A(_176_),
    .B(_170__bF$buf5),
    .C(_177_),
    .Y(_07_[4])
);

INVX2 _734_ (
    .A(mvect[5]),
    .Y(_178_)
);

NOR2X1 _735_ (
    .A(CSR_Wdata[5]),
    .B(_170__bF$buf4),
    .Y(_179_)
);

AOI21X1 _736_ (
    .A(_178_),
    .B(_170__bF$buf3),
    .C(_179_),
    .Y(_07_[5])
);

INVX2 _737_ (
    .A(mvect[6]),
    .Y(_180_)
);

NOR2X1 _738_ (
    .A(CSR_Wdata[6]),
    .B(_170__bF$buf2),
    .Y(_181_)
);

AOI21X1 _739_ (
    .A(_180_),
    .B(_170__bF$buf1),
    .C(_181_),
    .Y(_07_[6])
);

INVX1 _740_ (
    .A(mvect[7]),
    .Y(_182_)
);

NOR2X1 _741_ (
    .A(CSR_Wdata[7]),
    .B(_170__bF$buf0),
    .Y(_183_)
);

AOI21X1 _742_ (
    .A(_182_),
    .B(_170__bF$buf6),
    .C(_183_),
    .Y(_07_[7])
);

INVX1 _743_ (
    .A(mvect[8]),
    .Y(_184_)
);

NOR2X1 _744_ (
    .A(CSR_Wdata[8]),
    .B(_170__bF$buf5),
    .Y(_185_)
);

AOI21X1 _745_ (
    .A(_184_),
    .B(_170__bF$buf4),
    .C(_185_),
    .Y(_07_[8])
);

INVX1 _746_ (
    .A(mvect[9]),
    .Y(_186_)
);

NOR2X1 _747_ (
    .A(CSR_Wdata[9]),
    .B(_170__bF$buf3),
    .Y(_187_)
);

AOI21X1 _748_ (
    .A(_186_),
    .B(_170__bF$buf2),
    .C(_187_),
    .Y(_07_[9])
);

INVX2 _749_ (
    .A(mvect[10]),
    .Y(_188_)
);

NOR2X1 _750_ (
    .A(CSR_Wdata[10]),
    .B(_170__bF$buf1),
    .Y(_189_)
);

AOI21X1 _751_ (
    .A(_188_),
    .B(_170__bF$buf0),
    .C(_189_),
    .Y(_07_[10])
);

INVX1 _752_ (
    .A(mvect[11]),
    .Y(_190_)
);

INVX1 _753_ (
    .A(CSR_Wdata[11]),
    .Y(_191_)
);

MUX2X1 _754_ (
    .A(_190_),
    .B(_191_),
    .S(_170__bF$buf6),
    .Y(_07_[11])
);

INVX2 _755_ (
    .A(mvect[12]),
    .Y(_192_)
);

NOR2X1 _756_ (
    .A(CSR_Wdata[12]),
    .B(_170__bF$buf5),
    .Y(_193_)
);

AOI21X1 _757_ (
    .A(_192_),
    .B(_170__bF$buf4),
    .C(_193_),
    .Y(_07_[12])
);

INVX1 _758_ (
    .A(mvect[13]),
    .Y(_194_)
);

NOR2X1 _759_ (
    .A(CSR_Wdata[13]),
    .B(_170__bF$buf3),
    .Y(_195_)
);

AOI21X1 _760_ (
    .A(_194_),
    .B(_170__bF$buf2),
    .C(_195_),
    .Y(_07_[13])
);

INVX2 _761_ (
    .A(mvect[14]),
    .Y(_196_)
);

NOR2X1 _762_ (
    .A(CSR_Wdata[14]),
    .B(_170__bF$buf1),
    .Y(_197_)
);

AOI21X1 _763_ (
    .A(_196_),
    .B(_170__bF$buf0),
    .C(_197_),
    .Y(_07_[14])
);

INVX1 _764_ (
    .A(mvect[15]),
    .Y(_198_)
);

NOR2X1 _765_ (
    .A(CSR_Wdata[15]),
    .B(_170__bF$buf6),
    .Y(_199_)
);

AOI21X1 _766_ (
    .A(_198_),
    .B(_170__bF$buf5),
    .C(_199_),
    .Y(_07_[15])
);

INVX1 _767_ (
    .A(mvect[16]),
    .Y(_200_)
);

NOR2X1 _768_ (
    .A(CSR_Wdata[16]),
    .B(_170__bF$buf4),
    .Y(_201_)
);

AOI21X1 _769_ (
    .A(_200_),
    .B(_170__bF$buf3),
    .C(_201_),
    .Y(_07_[16])
);

INVX1 _770_ (
    .A(mvect[17]),
    .Y(_202_)
);

NOR2X1 _771_ (
    .A(CSR_Wdata[17]),
    .B(_170__bF$buf2),
    .Y(_203_)
);

AOI21X1 _772_ (
    .A(_202_),
    .B(_170__bF$buf1),
    .C(_203_),
    .Y(_07_[17])
);

INVX1 _773_ (
    .A(mvect[18]),
    .Y(_204_)
);

NOR2X1 _774_ (
    .A(CSR_Wdata[18]),
    .B(_170__bF$buf0),
    .Y(_205_)
);

AOI21X1 _775_ (
    .A(_204_),
    .B(_170__bF$buf6),
    .C(_205_),
    .Y(_07_[18])
);

INVX1 _776_ (
    .A(mvect[19]),
    .Y(_206_)
);

NOR2X1 _777_ (
    .A(CSR_Wdata[19]),
    .B(_170__bF$buf5),
    .Y(_207_)
);

AOI21X1 _778_ (
    .A(_206_),
    .B(_170__bF$buf4),
    .C(_207_),
    .Y(_07_[19])
);

INVX2 _779_ (
    .A(mvect[20]),
    .Y(_208_)
);

NOR2X1 _780_ (
    .A(CSR_Wdata[20]),
    .B(_170__bF$buf3),
    .Y(_209_)
);

AOI21X1 _781_ (
    .A(_208_),
    .B(_170__bF$buf2),
    .C(_209_),
    .Y(_07_[20])
);

INVX1 _782_ (
    .A(mvect[21]),
    .Y(_210_)
);

NOR2X1 _783_ (
    .A(CSR_Wdata[21]),
    .B(_170__bF$buf1),
    .Y(_211_)
);

AOI21X1 _784_ (
    .A(_210_),
    .B(_170__bF$buf0),
    .C(_211_),
    .Y(_07_[21])
);

INVX1 _785_ (
    .A(mvect[22]),
    .Y(_212_)
);

NOR2X1 _786_ (
    .A(CSR_Wdata[22]),
    .B(_170__bF$buf6),
    .Y(_213_)
);

AOI21X1 _787_ (
    .A(_212_),
    .B(_170__bF$buf5),
    .C(_213_),
    .Y(_07_[22])
);

INVX1 _788_ (
    .A(mvect[23]),
    .Y(_214_)
);

NOR2X1 _789_ (
    .A(CSR_Wdata[23]),
    .B(_170__bF$buf4),
    .Y(_215_)
);

AOI21X1 _790_ (
    .A(_214_),
    .B(_170__bF$buf3),
    .C(_215_),
    .Y(_07_[23])
);

INVX1 _791_ (
    .A(mvect[24]),
    .Y(_216_)
);

NOR2X1 _792_ (
    .A(CSR_Wdata[24]),
    .B(_170__bF$buf2),
    .Y(_217_)
);

AOI21X1 _793_ (
    .A(_216_),
    .B(_170__bF$buf1),
    .C(_217_),
    .Y(_07_[24])
);

INVX1 _794_ (
    .A(mvect[25]),
    .Y(_218_)
);

NOR2X1 _795_ (
    .A(CSR_Wdata[25]),
    .B(_170__bF$buf0),
    .Y(_219_)
);

AOI21X1 _796_ (
    .A(_218_),
    .B(_170__bF$buf6),
    .C(_219_),
    .Y(_07_[25])
);

INVX1 _797_ (
    .A(mvect[26]),
    .Y(_220_)
);

NOR2X1 _798_ (
    .A(CSR_Wdata[26]),
    .B(_170__bF$buf5),
    .Y(_221_)
);

AOI21X1 _799_ (
    .A(_220_),
    .B(_170__bF$buf4),
    .C(_221_),
    .Y(_07_[26])
);

INVX1 _800_ (
    .A(mvect[27]),
    .Y(_222_)
);

NOR2X1 _801_ (
    .A(CSR_Wdata[27]),
    .B(_170__bF$buf3),
    .Y(_223_)
);

AOI21X1 _802_ (
    .A(_222_),
    .B(_170__bF$buf2),
    .C(_223_),
    .Y(_07_[27])
);

INVX1 _803_ (
    .A(mvect[28]),
    .Y(_224_)
);

NOR2X1 _804_ (
    .A(CSR_Wdata[28]),
    .B(_170__bF$buf1),
    .Y(_225_)
);

AOI21X1 _805_ (
    .A(_224_),
    .B(_170__bF$buf0),
    .C(_225_),
    .Y(_07_[28])
);

INVX1 _806_ (
    .A(mvect[29]),
    .Y(_226_)
);

NOR2X1 _807_ (
    .A(CSR_Wdata[29]),
    .B(_170__bF$buf6),
    .Y(_227_)
);

AOI21X1 _808_ (
    .A(_226_),
    .B(_170__bF$buf5),
    .C(_227_),
    .Y(_07_[29])
);

INVX1 _809_ (
    .A(mvect[30]),
    .Y(_228_)
);

NOR2X1 _810_ (
    .A(CSR_Wdata[30]),
    .B(_170__bF$buf4),
    .Y(_229_)
);

AOI21X1 _811_ (
    .A(_228_),
    .B(_170__bF$buf3),
    .C(_229_),
    .Y(_07_[30])
);

INVX1 _812_ (
    .A(mvect[31]),
    .Y(_230_)
);

NOR2X1 _813_ (
    .A(CSR_Wdata[31]),
    .B(_170__bF$buf2),
    .Y(_231_)
);

AOI21X1 _814_ (
    .A(_230_),
    .B(_170__bF$buf1),
    .C(_231_),
    .Y(_07_[31])
);

NAND2X1 _815_ (
    .A(_169_),
    .B(_64_),
    .Y(_232_)
);

NAND2X1 _816_ (
    .A(mie),
    .B(_232_),
    .Y(_233_)
);

OAI21X1 _817_ (
    .A(_191_),
    .B(_232_),
    .C(_233_),
    .Y(_14_)
);

NAND2X1 _818_ (
    .A(CSR_Wen_traps_bF$buf2),
    .B(CSR_mepc[2]),
    .Y(_234_)
);

AND2X2 _819_ (
    .A(_31__bF$buf4),
    .B(_113_),
    .Y(_235_)
);

NOR2X1 _820_ (
    .A(mepc[0]),
    .B(_235__bF$buf4),
    .Y(_236_)
);

NAND2X1 _821_ (
    .A(_113_),
    .B(_31__bF$buf3),
    .Y(_237_)
);

OAI21X1 _822_ (
    .A(_237__bF$buf4),
    .B(CSR_Wdata[2]),
    .C(_112__bF$buf1),
    .Y(_238_)
);

OAI21X1 _823_ (
    .A(_236_),
    .B(_238_),
    .C(_234_),
    .Y(_21_[0])
);

NAND2X1 _824_ (
    .A(CSR_Wen_traps_bF$buf1),
    .B(CSR_mepc[3]),
    .Y(_239_)
);

NOR2X1 _825_ (
    .A(mepc[1]),
    .B(_235__bF$buf3),
    .Y(_240_)
);

OAI21X1 _826_ (
    .A(_237__bF$buf3),
    .B(CSR_Wdata[3]),
    .C(_112__bF$buf0),
    .Y(_241_)
);

OAI21X1 _827_ (
    .A(_240_),
    .B(_241_),
    .C(_239_),
    .Y(_21_[1])
);

NAND2X1 _828_ (
    .A(CSR_Wen_traps_bF$buf0),
    .B(CSR_mepc[4]),
    .Y(_242_)
);

NOR2X1 _829_ (
    .A(mepc[2]),
    .B(_235__bF$buf2),
    .Y(_243_)
);

OAI21X1 _830_ (
    .A(_237__bF$buf2),
    .B(CSR_Wdata[4]),
    .C(_112__bF$buf6),
    .Y(_244_)
);

OAI21X1 _831_ (
    .A(_243_),
    .B(_244_),
    .C(_242_),
    .Y(_21_[2])
);

NAND2X1 _832_ (
    .A(CSR_Wen_traps_bF$buf5),
    .B(CSR_mepc[5]),
    .Y(_245_)
);

NOR2X1 _833_ (
    .A(mepc[3]),
    .B(_235__bF$buf1),
    .Y(_246_)
);

OAI21X1 _834_ (
    .A(_237__bF$buf1),
    .B(CSR_Wdata[5]),
    .C(_112__bF$buf5),
    .Y(_247_)
);

OAI21X1 _835_ (
    .A(_246_),
    .B(_247_),
    .C(_245_),
    .Y(_21_[3])
);

NAND2X1 _836_ (
    .A(CSR_Wen_traps_bF$buf4),
    .B(CSR_mepc[6]),
    .Y(_248_)
);

NOR2X1 _837_ (
    .A(mepc[4]),
    .B(_235__bF$buf0),
    .Y(_249_)
);

OAI21X1 _838_ (
    .A(_237__bF$buf0),
    .B(CSR_Wdata[6]),
    .C(_112__bF$buf4),
    .Y(_250_)
);

OAI21X1 _839_ (
    .A(_249_),
    .B(_250_),
    .C(_248_),
    .Y(_21_[4])
);

NAND2X1 _840_ (
    .A(CSR_Wen_traps_bF$buf3),
    .B(CSR_mepc[7]),
    .Y(_251_)
);

NOR2X1 _841_ (
    .A(mepc[5]),
    .B(_235__bF$buf4),
    .Y(_252_)
);

OAI21X1 _842_ (
    .A(_237__bF$buf4),
    .B(CSR_Wdata[7]),
    .C(_112__bF$buf3),
    .Y(_253_)
);

OAI21X1 _843_ (
    .A(_252_),
    .B(_253_),
    .C(_251_),
    .Y(_21_[5])
);

NAND2X1 _844_ (
    .A(CSR_Wen_traps_bF$buf2),
    .B(CSR_mepc[8]),
    .Y(_254_)
);

NOR2X1 _845_ (
    .A(mepc[6]),
    .B(_235__bF$buf3),
    .Y(_255_)
);

OAI21X1 _846_ (
    .A(_237__bF$buf3),
    .B(CSR_Wdata[8]),
    .C(_112__bF$buf2),
    .Y(_256_)
);

OAI21X1 _847_ (
    .A(_255_),
    .B(_256_),
    .C(_254_),
    .Y(_21_[6])
);

NAND2X1 _848_ (
    .A(CSR_Wen_traps_bF$buf1),
    .B(CSR_mepc[9]),
    .Y(_257_)
);

NOR2X1 _849_ (
    .A(mepc[7]),
    .B(_235__bF$buf2),
    .Y(_258_)
);

OAI21X1 _850_ (
    .A(_237__bF$buf2),
    .B(CSR_Wdata[9]),
    .C(_112__bF$buf1),
    .Y(_259_)
);

OAI21X1 _851_ (
    .A(_258_),
    .B(_259_),
    .C(_257_),
    .Y(_21_[7])
);

NAND2X1 _852_ (
    .A(CSR_Wen_traps_bF$buf0),
    .B(CSR_mepc[10]),
    .Y(_260_)
);

NOR2X1 _853_ (
    .A(mepc[8]),
    .B(_235__bF$buf1),
    .Y(_261_)
);

OAI21X1 _854_ (
    .A(_237__bF$buf1),
    .B(CSR_Wdata[10]),
    .C(_112__bF$buf0),
    .Y(_262_)
);

OAI21X1 _855_ (
    .A(_261_),
    .B(_262_),
    .C(_260_),
    .Y(_21_[8])
);

NAND2X1 _856_ (
    .A(CSR_Wen_traps_bF$buf5),
    .B(CSR_mepc[11]),
    .Y(_263_)
);

NOR2X1 _857_ (
    .A(mepc[9]),
    .B(_235__bF$buf0),
    .Y(_264_)
);

OAI21X1 _858_ (
    .A(_237__bF$buf0),
    .B(CSR_Wdata[11]),
    .C(_112__bF$buf6),
    .Y(_265_)
);

OAI21X1 _859_ (
    .A(_264_),
    .B(_265_),
    .C(_263_),
    .Y(_21_[9])
);

NAND2X1 _860_ (
    .A(CSR_Wen_traps_bF$buf4),
    .B(CSR_mepc[12]),
    .Y(_266_)
);

NOR2X1 _861_ (
    .A(mepc[10]),
    .B(_235__bF$buf4),
    .Y(_267_)
);

OAI21X1 _862_ (
    .A(_237__bF$buf4),
    .B(CSR_Wdata[12]),
    .C(_112__bF$buf5),
    .Y(_268_)
);

OAI21X1 _863_ (
    .A(_267_),
    .B(_268_),
    .C(_266_),
    .Y(_21_[10])
);

NAND2X1 _864_ (
    .A(CSR_Wen_traps_bF$buf3),
    .B(CSR_mepc[13]),
    .Y(_269_)
);

NOR2X1 _865_ (
    .A(mepc[11]),
    .B(_235__bF$buf3),
    .Y(_270_)
);

OAI21X1 _866_ (
    .A(_237__bF$buf3),
    .B(CSR_Wdata[13]),
    .C(_112__bF$buf4),
    .Y(_271_)
);

OAI21X1 _867_ (
    .A(_270_),
    .B(_271_),
    .C(_269_),
    .Y(_21_[11])
);

NAND2X1 _868_ (
    .A(CSR_Wen_traps_bF$buf2),
    .B(CSR_mepc[14]),
    .Y(_272_)
);

NOR2X1 _869_ (
    .A(mepc[12]),
    .B(_235__bF$buf2),
    .Y(_273_)
);

OAI21X1 _870_ (
    .A(_237__bF$buf2),
    .B(CSR_Wdata[14]),
    .C(_112__bF$buf3),
    .Y(_274_)
);

OAI21X1 _871_ (
    .A(_273_),
    .B(_274_),
    .C(_272_),
    .Y(_21_[12])
);

NAND2X1 _872_ (
    .A(CSR_Wen_traps_bF$buf1),
    .B(CSR_mepc[15]),
    .Y(_275_)
);

NOR2X1 _873_ (
    .A(mepc[13]),
    .B(_235__bF$buf1),
    .Y(_276_)
);

OAI21X1 _874_ (
    .A(_237__bF$buf1),
    .B(CSR_Wdata[15]),
    .C(_112__bF$buf2),
    .Y(_277_)
);

OAI21X1 _875_ (
    .A(_276_),
    .B(_277_),
    .C(_275_),
    .Y(_21_[13])
);

NAND2X1 _876_ (
    .A(CSR_Wen_traps_bF$buf0),
    .B(CSR_mepc[16]),
    .Y(_278_)
);

NOR2X1 _877_ (
    .A(mepc[14]),
    .B(_235__bF$buf0),
    .Y(_279_)
);

OAI21X1 _878_ (
    .A(_237__bF$buf0),
    .B(CSR_Wdata[16]),
    .C(_112__bF$buf1),
    .Y(_280_)
);

OAI21X1 _879_ (
    .A(_279_),
    .B(_280_),
    .C(_278_),
    .Y(_21_[14])
);

NAND2X1 _880_ (
    .A(CSR_Wen_traps_bF$buf5),
    .B(CSR_mepc[17]),
    .Y(_281_)
);

NOR2X1 _881_ (
    .A(mepc[15]),
    .B(_235__bF$buf4),
    .Y(_282_)
);

OAI21X1 _882_ (
    .A(_237__bF$buf4),
    .B(CSR_Wdata[17]),
    .C(_112__bF$buf0),
    .Y(_283_)
);

OAI21X1 _883_ (
    .A(_282_),
    .B(_283_),
    .C(_281_),
    .Y(_21_[15])
);

NAND2X1 _884_ (
    .A(CSR_Wen_traps_bF$buf4),
    .B(CSR_mepc[18]),
    .Y(_284_)
);

NOR2X1 _885_ (
    .A(mepc[16]),
    .B(_235__bF$buf3),
    .Y(_285_)
);

OAI21X1 _886_ (
    .A(_237__bF$buf3),
    .B(CSR_Wdata[18]),
    .C(_112__bF$buf6),
    .Y(_286_)
);

OAI21X1 _887_ (
    .A(_285_),
    .B(_286_),
    .C(_284_),
    .Y(_21_[16])
);

NAND2X1 _888_ (
    .A(CSR_Wen_traps_bF$buf3),
    .B(CSR_mepc[19]),
    .Y(_287_)
);

NOR2X1 _889_ (
    .A(mepc[17]),
    .B(_235__bF$buf2),
    .Y(_288_)
);

OAI21X1 _890_ (
    .A(_237__bF$buf2),
    .B(CSR_Wdata[19]),
    .C(_112__bF$buf5),
    .Y(_289_)
);

OAI21X1 _891_ (
    .A(_288_),
    .B(_289_),
    .C(_287_),
    .Y(_21_[17])
);

NAND2X1 _892_ (
    .A(CSR_Wen_traps_bF$buf2),
    .B(CSR_mepc[20]),
    .Y(_290_)
);

NOR2X1 _893_ (
    .A(mepc[18]),
    .B(_235__bF$buf1),
    .Y(_291_)
);

OAI21X1 _894_ (
    .A(_237__bF$buf1),
    .B(CSR_Wdata[20]),
    .C(_112__bF$buf4),
    .Y(_292_)
);

OAI21X1 _895_ (
    .A(_291_),
    .B(_292_),
    .C(_290_),
    .Y(_21_[18])
);

NAND2X1 _896_ (
    .A(CSR_Wen_traps_bF$buf1),
    .B(CSR_mepc[21]),
    .Y(_293_)
);

NOR2X1 _897_ (
    .A(mepc[19]),
    .B(_235__bF$buf0),
    .Y(_294_)
);

OAI21X1 _898_ (
    .A(_237__bF$buf0),
    .B(CSR_Wdata[21]),
    .C(_112__bF$buf3),
    .Y(_295_)
);

OAI21X1 _899_ (
    .A(_294_),
    .B(_295_),
    .C(_293_),
    .Y(_21_[19])
);

NAND2X1 _900_ (
    .A(CSR_Wen_traps_bF$buf0),
    .B(CSR_mepc[22]),
    .Y(_296_)
);

NOR2X1 _901_ (
    .A(mepc[20]),
    .B(_235__bF$buf4),
    .Y(_297_)
);

OAI21X1 _902_ (
    .A(_237__bF$buf4),
    .B(CSR_Wdata[22]),
    .C(_112__bF$buf2),
    .Y(_298_)
);

OAI21X1 _903_ (
    .A(_297_),
    .B(_298_),
    .C(_296_),
    .Y(_21_[20])
);

NAND2X1 _904_ (
    .A(CSR_Wen_traps_bF$buf5),
    .B(CSR_mepc[23]),
    .Y(_299_)
);

NOR2X1 _905_ (
    .A(mepc[21]),
    .B(_235__bF$buf3),
    .Y(_300_)
);

OAI21X1 _906_ (
    .A(_237__bF$buf3),
    .B(CSR_Wdata[23]),
    .C(_112__bF$buf1),
    .Y(_301_)
);

OAI21X1 _907_ (
    .A(_300_),
    .B(_301_),
    .C(_299_),
    .Y(_21_[21])
);

NAND2X1 _908_ (
    .A(CSR_Wen_traps_bF$buf4),
    .B(CSR_mepc[24]),
    .Y(_302_)
);

NOR2X1 _909_ (
    .A(mepc[22]),
    .B(_235__bF$buf2),
    .Y(_303_)
);

OAI21X1 _910_ (
    .A(_237__bF$buf2),
    .B(CSR_Wdata[24]),
    .C(_112__bF$buf0),
    .Y(_304_)
);

OAI21X1 _911_ (
    .A(_303_),
    .B(_304_),
    .C(_302_),
    .Y(_21_[22])
);

NAND2X1 _912_ (
    .A(CSR_Wen_traps_bF$buf3),
    .B(CSR_mepc[25]),
    .Y(_305_)
);

NOR2X1 _913_ (
    .A(mepc[23]),
    .B(_235__bF$buf1),
    .Y(_306_)
);

OAI21X1 _914_ (
    .A(_237__bF$buf1),
    .B(CSR_Wdata[25]),
    .C(_112__bF$buf6),
    .Y(_307_)
);

OAI21X1 _915_ (
    .A(_306_),
    .B(_307_),
    .C(_305_),
    .Y(_21_[23])
);

NAND2X1 _916_ (
    .A(CSR_Wen_traps_bF$buf2),
    .B(CSR_mepc[26]),
    .Y(_308_)
);

NOR2X1 _917_ (
    .A(mepc[24]),
    .B(_235__bF$buf0),
    .Y(_309_)
);

OAI21X1 _918_ (
    .A(_237__bF$buf0),
    .B(CSR_Wdata[26]),
    .C(_112__bF$buf5),
    .Y(_310_)
);

OAI21X1 _919_ (
    .A(_309_),
    .B(_310_),
    .C(_308_),
    .Y(_21_[24])
);

NAND2X1 _920_ (
    .A(CSR_Wen_traps_bF$buf1),
    .B(CSR_mepc[27]),
    .Y(_311_)
);

NOR2X1 _921_ (
    .A(mepc[25]),
    .B(_235__bF$buf4),
    .Y(_312_)
);

OAI21X1 _922_ (
    .A(_237__bF$buf4),
    .B(CSR_Wdata[27]),
    .C(_112__bF$buf4),
    .Y(_313_)
);

OAI21X1 _923_ (
    .A(_312_),
    .B(_313_),
    .C(_311_),
    .Y(_21_[25])
);

NAND2X1 _924_ (
    .A(CSR_Wen_traps_bF$buf0),
    .B(CSR_mepc[28]),
    .Y(_314_)
);

NOR2X1 _925_ (
    .A(mepc[26]),
    .B(_235__bF$buf3),
    .Y(_315_)
);

OAI21X1 _926_ (
    .A(_237__bF$buf3),
    .B(CSR_Wdata[28]),
    .C(_112__bF$buf3),
    .Y(_316_)
);

OAI21X1 _927_ (
    .A(_315_),
    .B(_316_),
    .C(_314_),
    .Y(_21_[26])
);

NAND2X1 _928_ (
    .A(CSR_Wen_traps_bF$buf5),
    .B(CSR_mepc[29]),
    .Y(_317_)
);

NOR2X1 _929_ (
    .A(mepc[27]),
    .B(_235__bF$buf2),
    .Y(_318_)
);

OAI21X1 _930_ (
    .A(_237__bF$buf2),
    .B(CSR_Wdata[29]),
    .C(_112__bF$buf2),
    .Y(_319_)
);

OAI21X1 _931_ (
    .A(_318_),
    .B(_319_),
    .C(_317_),
    .Y(_21_[27])
);

NAND2X1 _932_ (
    .A(CSR_Wen_traps_bF$buf4),
    .B(CSR_mepc[30]),
    .Y(_320_)
);

NOR2X1 _933_ (
    .A(mepc[28]),
    .B(_235__bF$buf1),
    .Y(_321_)
);

OAI21X1 _934_ (
    .A(_237__bF$buf1),
    .B(CSR_Wdata[30]),
    .C(_112__bF$buf1),
    .Y(_322_)
);

OAI21X1 _935_ (
    .A(_321_),
    .B(_322_),
    .C(_320_),
    .Y(_21_[28])
);

NAND2X1 _936_ (
    .A(CSR_Wen_traps_bF$buf3),
    .B(CSR_mepc[31]),
    .Y(_323_)
);

NOR2X1 _937_ (
    .A(mepc[29]),
    .B(_235__bF$buf0),
    .Y(_324_)
);

OAI21X1 _938_ (
    .A(_237__bF$buf0),
    .B(CSR_Wdata[31]),
    .C(_112__bF$buf0),
    .Y(_325_)
);

OAI21X1 _939_ (
    .A(_324_),
    .B(_325_),
    .C(_323_),
    .Y(_21_[29])
);

NOR2X1 _940_ (
    .A(_0_),
    .B(_157_),
    .Y(_326_)
);

NAND2X1 _941_ (
    .A(_173_),
    .B(_326_),
    .Y(_327_)
);

INVX2 _942_ (
    .A(_326_),
    .Y(_328_)
);

AOI21X1 _943_ (
    .A(mvect[2]),
    .B(_328_),
    .C(CSR_Ret_bF$buf3),
    .Y(_329_)
);

NOR2X1 _944_ (
    .A(mepc[0]),
    .B(_108__bF$buf0),
    .Y(_330_)
);

AOI21X1 _945_ (
    .A(_327_),
    .B(_329_),
    .C(_330_),
    .Y(_486_[2])
);

XNOR2X1 _946_ (
    .A(_327_),
    .B(_175_),
    .Y(_331_)
);

NAND2X1 _947_ (
    .A(mepc[1]),
    .B(CSR_Ret_bF$buf2),
    .Y(_332_)
);

OAI21X1 _948_ (
    .A(_331_),
    .B(CSR_Ret_bF$buf1),
    .C(_332_),
    .Y(_486_[3])
);

NOR2X1 _949_ (
    .A(mvect[2]),
    .B(mvect[3]),
    .Y(_333_)
);

OAI21X1 _950_ (
    .A(_328_),
    .B(_333_),
    .C(_176_),
    .Y(_334_)
);

OAI21X1 _951_ (
    .A(mvect[2]),
    .B(mvect[3]),
    .C(mvect[4]),
    .Y(_335_)
);

OAI21X1 _952_ (
    .A(_328_),
    .B(_335_),
    .C(_334_),
    .Y(_336_)
);

NAND2X1 _953_ (
    .A(mepc[2]),
    .B(CSR_Ret_bF$buf0),
    .Y(_337_)
);

OAI21X1 _954_ (
    .A(_336_),
    .B(CSR_Ret_bF$buf5),
    .C(_337_),
    .Y(_486_[4])
);

OAI21X1 _955_ (
    .A(_176_),
    .B(_333_),
    .C(_326_),
    .Y(_338_)
);

XNOR2X1 _956_ (
    .A(_338_),
    .B(_178_),
    .Y(_339_)
);

NAND2X1 _957_ (
    .A(mepc[3]),
    .B(CSR_Ret_bF$buf4),
    .Y(_340_)
);

OAI21X1 _958_ (
    .A(_339_),
    .B(CSR_Ret_bF$buf3),
    .C(_340_),
    .Y(_486_[5])
);

OAI21X1 _959_ (
    .A(_333_),
    .B(_176_),
    .C(_178_),
    .Y(_341_)
);

AOI21X1 _960_ (
    .A(_326_),
    .B(_341_),
    .C(mvect[6]),
    .Y(_342_)
);

NAND2X1 _961_ (
    .A(_326_),
    .B(_341_),
    .Y(_343_)
);

OAI21X1 _962_ (
    .A(_343_),
    .B(_180_),
    .C(_108__bF$buf4),
    .Y(_344_)
);

NAND2X1 _963_ (
    .A(mepc[4]),
    .B(CSR_Ret_bF$buf2),
    .Y(_345_)
);

OAI21X1 _964_ (
    .A(_344_),
    .B(_342_),
    .C(_345_),
    .Y(_486_[6])
);

OAI21X1 _965_ (
    .A(_343_),
    .B(_180_),
    .C(_182_),
    .Y(_346_)
);

NAND2X1 _966_ (
    .A(mvect[6]),
    .B(mvect[7]),
    .Y(_347_)
);

OAI21X1 _967_ (
    .A(_343_),
    .B(_347_),
    .C(_346_),
    .Y(_348_)
);

NAND2X1 _968_ (
    .A(mepc[5]),
    .B(CSR_Ret_bF$buf1),
    .Y(_349_)
);

OAI21X1 _969_ (
    .A(_348_),
    .B(CSR_Ret_bF$buf0),
    .C(_349_),
    .Y(_486_[7])
);

AOI21X1 _970_ (
    .A(_178_),
    .B(_335_),
    .C(_347_),
    .Y(_350_)
);

AND2X2 _971_ (
    .A(_350_),
    .B(_326_),
    .Y(_351_)
);

NAND2X1 _972_ (
    .A(mvect[8]),
    .B(_351_),
    .Y(_352_)
);

INVX1 _973_ (
    .A(_352_),
    .Y(_353_)
);

OAI21X1 _974_ (
    .A(_351_),
    .B(mvect[8]),
    .C(_108__bF$buf3),
    .Y(_354_)
);

NAND2X1 _975_ (
    .A(mepc[6]),
    .B(CSR_Ret_bF$buf5),
    .Y(_355_)
);

OAI21X1 _976_ (
    .A(_353_),
    .B(_354_),
    .C(_355_),
    .Y(_486_[8])
);

NAND2X1 _977_ (
    .A(_326_),
    .B(_350_),
    .Y(_356_)
);

OAI21X1 _978_ (
    .A(_356_),
    .B(_184_),
    .C(_186_),
    .Y(_357_)
);

NAND2X1 _979_ (
    .A(mvect[8]),
    .B(mvect[9]),
    .Y(_358_)
);

OAI21X1 _980_ (
    .A(_356_),
    .B(_358_),
    .C(_357_),
    .Y(_359_)
);

NAND2X1 _981_ (
    .A(mepc[7]),
    .B(CSR_Ret_bF$buf4),
    .Y(_360_)
);

OAI21X1 _982_ (
    .A(_359_),
    .B(CSR_Ret_bF$buf3),
    .C(_360_),
    .Y(_486_[9])
);

INVX1 _983_ (
    .A(_358_),
    .Y(_361_)
);

NAND2X1 _984_ (
    .A(_361_),
    .B(_351_),
    .Y(_362_)
);

XNOR2X1 _985_ (
    .A(_362_),
    .B(_188_),
    .Y(_363_)
);

NAND2X1 _986_ (
    .A(mepc[8]),
    .B(CSR_Ret_bF$buf2),
    .Y(_364_)
);

OAI21X1 _987_ (
    .A(_363_),
    .B(CSR_Ret_bF$buf1),
    .C(_364_),
    .Y(_486_[10])
);

NAND2X1 _988_ (
    .A(mvect[10]),
    .B(_361_),
    .Y(_365_)
);

OAI21X1 _989_ (
    .A(_356_),
    .B(_365_),
    .C(_190_),
    .Y(_366_)
);

NAND2X1 _990_ (
    .A(mvect[10]),
    .B(mvect[11]),
    .Y(_367_)
);

OR2X2 _991_ (
    .A(_358_),
    .B(_367_),
    .Y(_368_)
);

OAI21X1 _992_ (
    .A(_356_),
    .B(_368_),
    .C(_366_),
    .Y(_369_)
);

NAND2X1 _993_ (
    .A(mepc[9]),
    .B(CSR_Ret_bF$buf0),
    .Y(_370_)
);

OAI21X1 _994_ (
    .A(_369_),
    .B(CSR_Ret_bF$buf5),
    .C(_370_),
    .Y(_486_[11])
);

NOR2X1 _995_ (
    .A(_358_),
    .B(_367_),
    .Y(_371_)
);

NAND3X1 _996_ (
    .A(_326_),
    .B(_371_),
    .C(_350_),
    .Y(_372_)
);

XNOR2X1 _997_ (
    .A(_372_),
    .B(_192_),
    .Y(_373_)
);

NAND2X1 _998_ (
    .A(mepc[10]),
    .B(CSR_Ret_bF$buf4),
    .Y(_374_)
);

OAI21X1 _999_ (
    .A(_373_),
    .B(CSR_Ret_bF$buf3),
    .C(_374_),
    .Y(_486_[12])
);

endmodule
