/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */

module csr(
    inout vdd,
    inout gnd,
    output CSR_IRQ,
    output [31:0] CSR_PCaddr,
    input CSR_Ret,
    input [31:0] CSR_Wdata,
    input CSR_Wen,
    input CSR_Wen_traps,
    input [11:0] CSR_addr,
    output [31:0] CSR_data,
    input [3:0] CSR_mcause,
    input [31:0] CSR_mepc,
    input Extern_IRQ,
    input clk
);

wire _168_ ;
wire _60_ ;
wire _397_ ;
wire _19_ ;
wire _321_ ;
wire _57_ ;
wire _130_ ;
wire _415_ ;
wire _95_ ;
wire _224_ ;
wire _453_ ;
wire _262_ ;
wire _318_ ;
wire _127_ ;
wire _356_ ;
wire _165_ ;
wire _394_ ;
wire _259_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _412_ ;
wire _92_ ;
wire _221_ ;
wire _450_ ;
wire _315_ ;
wire _124_ ;
wire _353_ ;
wire _409_ ;
wire _89_ ;
wire _162_ ;
wire _218_ ;
wire _391_ ;
wire _447_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _159_ ;
wire _51_ ;
wire _388_ ;
wire _197_ ;
wire _7_ ;
wire _312_ ;
wire _48_ ;
wire _121_ ;
wire _350_ ;
wire _406_ ;
wire _86_ ;
wire _215_ ;
wire _444_ ;
wire _253_ ;
wire _309_ ;
wire _482_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _347_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire [31:0] _07_ ;
wire _45_ ;
wire _403_ ;
wire _83_ ;
wire _212_ ;
wire _441_ ;
wire _250_ ;
wire _306_ ;
wire _115_ ;
wire _344_ ;
wire _153_ ;
wire _209_ ;
wire _382_ ;
wire _438_ ;
wire _191_ ;
wire _247_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire _285_ ;
wire _1_ ;
wire [1:0] mstatus ;
wire _42_ ;
wire _379_ ;
wire _188_ ;
wire _400_ ;
wire _80_ ;
wire _303_ ;
wire _39_ ;
wire _112_ ;
wire _341_ ;
wire clk ;
wire _77_ ;
wire _150_ ;
wire _206_ ;
wire _435_ ;
wire _244_ ;
wire _473_ ;
wire _109_ ;
wire _282_ ;
wire _338_ ;
wire CSR_IRQ ;
wire _147_ ;
wire _376_ ;
wire _235__bF$buf0 ;
wire _235__bF$buf1 ;
wire _235__bF$buf2 ;
wire _235__bF$buf3 ;
wire _235__bF$buf4 ;
wire _185_ ;
wire _279_ ;
wire _300_ ;
wire _36_ ;
wire _74_ ;
wire _203_ ;
wire _432_ ;
wire _241_ ;
wire _470_ ;
wire _106_ ;
wire _335_ ;
wire _144_ ;
wire _373_ ;
wire _429_ ;
wire _182_ ;
wire _238_ ;
wire _467_ ;
wire _276_ ;
wire [1:0] _33_ ;
wire _179_ ;
wire _71_ ;
wire _200_ ;
wire _103_ ;
wire _332_ ;
wire _68_ ;
wire _141_ ;
wire _370_ ;
wire _426_ ;
wire _235_ ;
wire _464_ ;
wire _273_ ;
wire _329_ ;
wire _138_ ;
wire _30_ ;
wire _367_ ;
wire _176_ ;
wire _27_ ;
wire _100_ ;
wire _65_ ;
wire _423_ ;
wire _232_ ;
wire _461_ ;
wire _270_ ;
wire _326_ ;
wire _135_ ;
wire _364_ ;
wire CSR_Wen_traps ;
wire _114__bF$buf0 ;
wire _114__bF$buf1 ;
wire _114__bF$buf2 ;
wire _114__bF$buf3 ;
wire _114__bF$buf4 ;
wire _114__bF$buf5 ;
wire _114__bF$buf6 ;
wire _173_ ;
wire _229_ ;
wire _458_ ;
wire _267_ ;
wire _24_ ;
wire [31:0] CSR_mepc ;
wire _62_ ;
wire _399_ ;
wire _420_ ;
wire _323_ ;
wire _59_ ;
wire _132_ ;
wire _361_ ;
wire _417_ ;
wire _97_ ;
wire _170_ ;
wire _226_ ;
wire _455_ ;
wire _264_ ;
wire [11:0] CSR_addr ;
wire _129_ ;
wire [29:0] _21_ ;
wire _358_ ;
wire _167_ ;
wire _396_ ;
wire _299_ ;
wire _18_ ;
wire _320_ ;
wire _56_ ;
wire _414_ ;
wire _94_ ;
wire _223_ ;
wire _452_ ;
wire _261_ ;
wire _317_ ;
wire _126_ ;
wire _355_ ;
wire _164_ ;
wire _393_ ;
wire [31:0] CSR_PCaddr ;
wire _449_ ;
wire _258_ ;
wire [31:0] _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _199_ ;
wire _411_ ;
wire _91_ ;
wire _220_ ;
wire _9_ ;
wire _108__bF$buf0 ;
wire _108__bF$buf1 ;
wire _108__bF$buf2 ;
wire _108__bF$buf3 ;
wire _108__bF$buf4 ;
wire _314_ ;
wire _123_ ;
wire _352_ ;
wire _408_ ;
wire _88_ ;
wire _161_ ;
wire _217_ ;
wire _390_ ;
wire _446_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _349_ ;
wire _158_ ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _311_ ;
wire _47_ ;
wire _120_ ;
wire _405_ ;
wire _85_ ;
wire _214_ ;
wire _443_ ;
wire _252_ ;
wire CSR_Ret_bF$buf0 ;
wire CSR_Ret_bF$buf1 ;
wire CSR_Ret_bF$buf2 ;
wire CSR_Ret_bF$buf3 ;
wire CSR_Ret_bF$buf4 ;
wire CSR_Ret_bF$buf5 ;
wire _308_ ;
wire _481_ ;
wire _117_ ;
wire _290_ ;
wire _346_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _249_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _402_ ;
wire _82_ ;
wire _211_ ;
wire _440_ ;
wire _305_ ;
wire _114_ ;
wire _343_ ;
wire _79_ ;
wire _152_ ;
wire _208_ ;
wire _381_ ;
wire _437_ ;
wire _190_ ;
wire _246_ ;
wire _475_ ;
wire _284_ ;
wire _0_ ;
wire Extern_IRQ ;
wire _149_ ;
wire _41_ ;
wire _378_ ;
wire _187_ ;
wire _302_ ;
wire [3:0] CSR_mcause ;
wire _38_ ;
wire _111_ ;
wire _340_ ;
wire _76_ ;
wire _205_ ;
wire _434_ ;
wire _243_ ;
wire _472_ ;
wire _108_ ;
wire _281_ ;
wire _337_ ;
wire _146_ ;
wire _375_ ;
wire _184_ ;
wire _469_ ;
wire _278_ ;
wire _35_ ;
wire _73_ ;
wire _202_ ;
wire _431_ ;
wire _240_ ;
wire _105_ ;
wire _334_ ;
wire _143_ ;
wire _372_ ;
wire _428_ ;
wire _181_ ;
wire _237_ ;
wire _466_ ;
wire _275_ ;
wire [31:0] CSR_Wdata ;
wire _32_ ;
wire _369_ ;
wire _178_ ;
wire _70_ ;
wire _170__bF$buf0 ;
wire _170__bF$buf1 ;
wire _170__bF$buf2 ;
wire _170__bF$buf3 ;
wire _170__bF$buf4 ;
wire _170__bF$buf5 ;
wire _170__bF$buf6 ;
wire _29_ ;
wire _102_ ;
wire _331_ ;
wire _67_ ;
wire _140_ ;
wire _425_ ;
wire _234_ ;
wire _463_ ;
wire _272_ ;
wire _328_ ;
wire _137_ ;
wire _366_ ;
wire _175_ ;
wire _269_ ;
wire _26_ ;
wire _64_ ;
wire _422_ ;
wire _231_ ;
wire _460_ ;
wire _325_ ;
wire _134_ ;
wire _363_ ;
wire _419_ ;
wire _99_ ;
wire _172_ ;
wire _228_ ;
wire _457_ ;
wire [29:0] mepc ;
wire _266_ ;
wire _23_ ;
wire _169_ ;
wire _61_ ;
wire _398_ ;
wire meta_irq ;
wire _322_ ;
wire _58_ ;
wire _131_ ;
wire _360_ ;
wire _416_ ;
wire _96_ ;
wire _225_ ;
wire _454_ ;
wire _263_ ;
wire _319_ ;
wire _128_ ;
wire _20_ ;
wire _357_ ;
wire _166_ ;
wire _395_ ;
wire _298_ ;
wire _11__bF$buf0 ;
wire _11__bF$buf1 ;
wire _11__bF$buf2 ;
wire _11__bF$buf3 ;
wire _11__bF$buf4 ;
wire _17_ ;
wire _55_ ;
wire _413_ ;
wire _93_ ;
wire _222_ ;
wire _112__bF$buf0 ;
wire _112__bF$buf1 ;
wire _112__bF$buf2 ;
wire _112__bF$buf3 ;
wire _112__bF$buf4 ;
wire _112__bF$buf5 ;
wire _112__bF$buf6 ;
wire _451_ ;
wire _260_ ;
wire _316_ ;
wire _125_ ;
wire _354_ ;
wire _163_ ;
wire _219_ ;
wire _392_ ;
wire _448_ ;
wire _257_ ;
wire [31:0] _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _198_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _313_ ;
wire _49_ ;
wire _122_ ;
wire _351_ ;
wire _407_ ;
wire _87_ ;
wire _160_ ;
wire _216_ ;
wire CSR_Wen ;
wire _445_ ;
wire _254_ ;
wire _483_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _348_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire _289_ ;
wire _5_ ;
wire _310_ ;
wire _237__bF$buf0 ;
wire _237__bF$buf1 ;
wire _237__bF$buf2 ;
wire _237__bF$buf3 ;
wire _237__bF$buf4 ;
wire _46_ ;
wire _404_ ;
wire _84_ ;
wire _213_ ;
wire _442_ ;
wire _251_ ;
wire _307_ ;
wire _480_ ;
wire _116_ ;
wire _345_ ;
wire _154_ ;
wire _383_ ;
wire _439_ ;
wire _192_ ;
wire _248_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _24__bF$buf0 ;
wire _24__bF$buf1 ;
wire _24__bF$buf2 ;
wire _24__bF$buf3 ;
wire _24__bF$buf4 ;
wire _401_ ;
wire _81_ ;
wire _210_ ;
wire _304_ ;
wire _113_ ;
wire _342_ ;
wire _78_ ;
wire _151_ ;
wire _207_ ;
wire _380_ ;
wire _436_ ;
wire _245_ ;
wire _474_ ;
wire _283_ ;
wire _339_ ;
wire CSR_Wen_traps_bF$buf0 ;
wire CSR_Wen_traps_bF$buf1 ;
wire CSR_Wen_traps_bF$buf2 ;
wire CSR_Wen_traps_bF$buf3 ;
wire CSR_Wen_traps_bF$buf4 ;
wire CSR_Wen_traps_bF$buf5 ;
wire _148_ ;
wire _40_ ;
wire _377_ ;
wire _186_ ;
wire _31__bF$buf0 ;
wire _31__bF$buf1 ;
wire _31__bF$buf2 ;
wire _31__bF$buf3 ;
wire _31__bF$buf4 ;
wire _301_ ;
wire _37_ ;
wire _110_ ;
wire CSR_Ret ;
wire _75_ ;
wire _204_ ;
wire _433_ ;
wire _242_ ;
wire _471_ ;
wire _107_ ;
wire _280_ ;
wire _336_ ;
wire _145_ ;
wire _374_ ;
wire _183_ ;
wire _239_ ;
wire _468_ ;
wire _277_ ;
wire [31:0] mvect ;
wire _34_ ;
wire _72_ ;
wire _201_ ;
wire _430_ ;
wire _104_ ;
wire _333_ ;
wire _69_ ;
wire _142_ ;
wire _371_ ;
wire _427_ ;
wire _180_ ;
wire _236_ ;
wire _465_ ;
wire _274_ ;
wire _139_ ;
wire _31_ ;
wire _368_ ;
wire _177_ ;
wire [31:0] _28_ ;
wire _101_ ;
wire _330_ ;
wire _66_ ;
wire _424_ ;
wire _233_ ;
wire _462_ ;
wire _271_ ;
wire _327_ ;
wire _136_ ;
wire _365_ ;
wire _174_ ;
wire _459_ ;
wire _268_ ;
wire _25_ ;
wire _63_ ;
wire _421_ ;
wire _230_ ;
wire [31:0] CSR_data ;
wire [31:0] mcause ;
wire _324_ ;
wire _133_ ;
wire _362_ ;
wire _418_ ;
wire _98_ ;
wire _171_ ;
wire _227_ ;
wire _456_ ;
wire _265_ ;
wire mie ;
wire mip ;
wire _22_ ;
wire _359_ ;

BUFX2 BUFX2_insert71 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_31_),
    .Y(_31__bF$buf0)
);

BUFX2 BUFX2_insert70 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_31_),
    .Y(_31__bF$buf1)
);

BUFX2 BUFX2_insert69 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_31_),
    .Y(_31__bF$buf2)
);

BUFX2 BUFX2_insert68 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_31_),
    .Y(_31__bF$buf3)
);

BUFX2 BUFX2_insert67 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_31_),
    .Y(_31__bF$buf4)
);

BUFX2 BUFX2_insert66 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Ret),
    .Y(CSR_Ret_bF$buf0)
);

BUFX2 BUFX2_insert65 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Ret),
    .Y(CSR_Ret_bF$buf1)
);

BUFX2 BUFX2_insert64 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Ret),
    .Y(CSR_Ret_bF$buf2)
);

BUFX2 BUFX2_insert63 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Ret),
    .Y(CSR_Ret_bF$buf3)
);

BUFX2 BUFX2_insert62 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Ret),
    .Y(CSR_Ret_bF$buf4)
);

BUFX2 BUFX2_insert61 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Ret),
    .Y(CSR_Ret_bF$buf5)
);

BUFX2 BUFX2_insert60 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11_),
    .Y(_11__bF$buf0)
);

BUFX2 BUFX2_insert59 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11_),
    .Y(_11__bF$buf1)
);

BUFX2 BUFX2_insert58 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11_),
    .Y(_11__bF$buf2)
);

BUFX2 BUFX2_insert57 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11_),
    .Y(_11__bF$buf3)
);

BUFX2 BUFX2_insert56 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11_),
    .Y(_11__bF$buf4)
);

BUFX2 BUFX2_insert55 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237_),
    .Y(_237__bF$buf0)
);

BUFX2 BUFX2_insert54 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237_),
    .Y(_237__bF$buf1)
);

BUFX2 BUFX2_insert53 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237_),
    .Y(_237__bF$buf2)
);

BUFX2 BUFX2_insert52 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237_),
    .Y(_237__bF$buf3)
);

BUFX2 BUFX2_insert51 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237_),
    .Y(_237__bF$buf4)
);

BUFX2 BUFX2_insert50 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_108_),
    .Y(_108__bF$buf0)
);

BUFX2 BUFX2_insert49 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_108_),
    .Y(_108__bF$buf1)
);

BUFX2 BUFX2_insert48 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_108_),
    .Y(_108__bF$buf2)
);

BUFX2 BUFX2_insert47 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_108_),
    .Y(_108__bF$buf3)
);

BUFX2 BUFX2_insert46 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_108_),
    .Y(_108__bF$buf4)
);

BUFX2 BUFX2_insert45 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114_),
    .Y(_114__bF$buf0)
);

BUFX2 BUFX2_insert44 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114_),
    .Y(_114__bF$buf1)
);

BUFX2 BUFX2_insert43 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114_),
    .Y(_114__bF$buf2)
);

BUFX2 BUFX2_insert42 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114_),
    .Y(_114__bF$buf3)
);

BUFX2 BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114_),
    .Y(_114__bF$buf4)
);

BUFX2 BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114_),
    .Y(_114__bF$buf5)
);

BUFX2 BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114_),
    .Y(_114__bF$buf6)
);

BUFX2 BUFX2_insert38 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .Y(_170__bF$buf0)
);

BUFX2 BUFX2_insert37 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .Y(_170__bF$buf1)
);

BUFX2 BUFX2_insert36 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .Y(_170__bF$buf2)
);

BUFX2 BUFX2_insert35 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .Y(_170__bF$buf3)
);

BUFX2 BUFX2_insert34 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .Y(_170__bF$buf4)
);

BUFX2 BUFX2_insert33 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .Y(_170__bF$buf5)
);

BUFX2 BUFX2_insert32 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .Y(_170__bF$buf6)
);

BUFX2 BUFX2_insert31 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24_),
    .Y(_24__bF$buf0)
);

BUFX2 BUFX2_insert30 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24_),
    .Y(_24__bF$buf1)
);

BUFX2 BUFX2_insert29 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24_),
    .Y(_24__bF$buf2)
);

BUFX2 BUFX2_insert28 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24_),
    .Y(_24__bF$buf3)
);

BUFX2 BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24_),
    .Y(_24__bF$buf4)
);

BUFX2 BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps),
    .Y(CSR_Wen_traps_bF$buf0)
);

BUFX2 BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps),
    .Y(CSR_Wen_traps_bF$buf1)
);

BUFX2 BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps),
    .Y(CSR_Wen_traps_bF$buf2)
);

BUFX2 BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps),
    .Y(CSR_Wen_traps_bF$buf3)
);

BUFX2 BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps),
    .Y(CSR_Wen_traps_bF$buf4)
);

BUFX2 BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps),
    .Y(CSR_Wen_traps_bF$buf5)
);

BUFX2 BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_235_),
    .Y(_235__bF$buf0)
);

BUFX2 BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_235_),
    .Y(_235__bF$buf1)
);

BUFX2 BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_235_),
    .Y(_235__bF$buf2)
);

BUFX2 BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_235_),
    .Y(_235__bF$buf3)
);

BUFX2 BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_235_),
    .Y(_235__bF$buf4)
);

CLKBUF1 CLKBUF1_insert15 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert14 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert13 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert12 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert11 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert10 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert9 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert8 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert7 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf8)
);

BUFX2 BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112_),
    .Y(_112__bF$buf0)
);

BUFX2 BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112_),
    .Y(_112__bF$buf1)
);

BUFX2 BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112_),
    .Y(_112__bF$buf2)
);

BUFX2 BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112_),
    .Y(_112__bF$buf3)
);

BUFX2 BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112_),
    .Y(_112__bF$buf4)
);

BUFX2 BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112_),
    .Y(_112__bF$buf5)
);

BUFX2 BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112_),
    .Y(_112__bF$buf6)
);

NAND2X1 _1000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[11]),
    .B(CSR_Ret_bF$buf5),
    .Y(_375_)
);

OAI21X1 _1001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_372_),
    .B(_192_),
    .C(_194_),
    .Y(_376_)
);

INVX1 _1002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_376_),
    .Y(_377_)
);

NAND2X1 _1003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[12]),
    .B(mvect[13]),
    .Y(_378_)
);

OAI21X1 _1004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_372_),
    .B(_378_),
    .C(_108__bF$buf4),
    .Y(_379_)
);

OAI21X1 _1005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_377_),
    .B(_379_),
    .C(_375_),
    .Y(_486_[13])
);

NAND2X1 _1006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[12]),
    .B(CSR_Ret_bF$buf4),
    .Y(_380_)
);

OAI21X1 _1007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_372_),
    .B(_378_),
    .C(_196_),
    .Y(_381_)
);

INVX1 _1008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_381_),
    .Y(_382_)
);

OR2X2 _1009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_372_),
    .B(_378_),
    .Y(_383_)
);

OAI21X1 _1010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_383_),
    .B(_196_),
    .C(_108__bF$buf3),
    .Y(_384_)
);

OAI21X1 _1011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_384_),
    .B(_382_),
    .C(_380_),
    .Y(_486_[14])
);

NAND2X1 _1012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[13]),
    .B(CSR_Ret_bF$buf3),
    .Y(_385_)
);

OAI21X1 _1013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_383_),
    .B(_196_),
    .C(_198_),
    .Y(_386_)
);

INVX1 _1014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_386_),
    .Y(_387_)
);

NAND2X1 _1015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[14]),
    .B(mvect[15]),
    .Y(_388_)
);

OR2X2 _1016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_378_),
    .B(_388_),
    .Y(_389_)
);

OAI21X1 _1017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_372_),
    .B(_389_),
    .C(_108__bF$buf2),
    .Y(_390_)
);

OAI21X1 _1018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_387_),
    .B(_390_),
    .C(_385_),
    .Y(_486_[15])
);

NAND2X1 _1019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[14]),
    .B(CSR_Ret_bF$buf2),
    .Y(_391_)
);

NOR2X1 _1020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_389_),
    .B(_372_),
    .Y(_392_)
);

NOR2X1 _1021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_378_),
    .B(_388_),
    .Y(_393_)
);

NAND3X1 _1022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_371_),
    .B(_393_),
    .C(_350_),
    .Y(_394_)
);

NOR2X1 _1023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_328_),
    .B(_394_),
    .Y(_395_)
);

NAND2X1 _1024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[16]),
    .B(_395_),
    .Y(_396_)
);

OAI21X1 _1025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[16]),
    .B(_392_),
    .C(_396_),
    .Y(_397_)
);

OAI21X1 _1026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_397_),
    .B(CSR_Ret_bF$buf1),
    .C(_391_),
    .Y(_486_[16])
);

NAND2X1 _1027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[15]),
    .B(CSR_Ret_bF$buf0),
    .Y(_398_)
);

AOI21X1 _1028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[16]),
    .B(_395_),
    .C(mvect[17]),
    .Y(_399_)
);

INVX2 _1029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_392_),
    .Y(_400_)
);

NAND2X1 _1030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[16]),
    .B(mvect[17]),
    .Y(_401_)
);

OAI21X1 _1031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_400_),
    .B(_401_),
    .C(_108__bF$buf1),
    .Y(_402_)
);

OAI21X1 _1032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_402_),
    .B(_399_),
    .C(_398_),
    .Y(_486_[17])
);

NAND2X1 _1033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[16]),
    .B(CSR_Ret_bF$buf5),
    .Y(_403_)
);

AND2X2 _1034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[16]),
    .B(mvect[17]),
    .Y(_404_)
);

AOI21X1 _1035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_404_),
    .B(_392_),
    .C(mvect[18]),
    .Y(_405_)
);

NAND2X1 _1036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[18]),
    .B(_404_),
    .Y(_406_)
);

OAI21X1 _1037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_400_),
    .B(_406_),
    .C(_108__bF$buf0),
    .Y(_407_)
);

OAI21X1 _1038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_407_),
    .B(_405_),
    .C(_403_),
    .Y(_486_[18])
);

NAND2X1 _1039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[17]),
    .B(CSR_Ret_bF$buf4),
    .Y(_408_)
);

INVX1 _1040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_406_),
    .Y(_409_)
);

AOI21X1 _1041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_409_),
    .B(_395_),
    .C(mvect[19]),
    .Y(_410_)
);

AND2X2 _1042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[18]),
    .B(mvect[19]),
    .Y(_411_)
);

NAND2X1 _1043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_404_),
    .B(_411_),
    .Y(_412_)
);

OAI21X1 _1044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_400_),
    .B(_412_),
    .C(_108__bF$buf4),
    .Y(_413_)
);

OAI21X1 _1045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_413_),
    .B(_410_),
    .C(_408_),
    .Y(_486_[19])
);

NAND2X1 _1046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[18]),
    .B(CSR_Ret_bF$buf3),
    .Y(_414_)
);

NAND3X1 _1047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_404_),
    .B(_411_),
    .C(_392_),
    .Y(_415_)
);

AND2X2 _1048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_415_),
    .B(_208_),
    .Y(_416_)
);

OAI21X1 _1049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_415_),
    .B(_208_),
    .C(_108__bF$buf3),
    .Y(_417_)
);

OAI21X1 _1050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_416_),
    .B(_417_),
    .C(_414_),
    .Y(_486_[20])
);

NAND2X1 _1051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[19]),
    .B(CSR_Ret_bF$buf2),
    .Y(_418_)
);

NOR2X1 _1052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_208_),
    .B(_412_),
    .Y(_419_)
);

AOI21X1 _1053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_419_),
    .B(_395_),
    .C(mvect[21]),
    .Y(_420_)
);

AND2X2 _1054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[20]),
    .B(mvect[21]),
    .Y(_421_)
);

NAND3X1 _1055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_404_),
    .B(_411_),
    .C(_421_),
    .Y(_422_)
);

OAI21X1 _1056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_400_),
    .B(_422_),
    .C(_108__bF$buf2),
    .Y(_423_)
);

OAI21X1 _1057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_423_),
    .B(_420_),
    .C(_418_),
    .Y(_486_[21])
);

NAND2X1 _1058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[20]),
    .B(CSR_Ret_bF$buf1),
    .Y(_424_)
);

NAND2X1 _1059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[18]),
    .B(mvect[19]),
    .Y(_425_)
);

NAND2X1 _1060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[20]),
    .B(mvect[21]),
    .Y(_426_)
);

NOR3X1 _1061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_401_),
    .B(_425_),
    .C(_426_),
    .Y(_427_)
);

NAND3X1 _1062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_371_),
    .B(_393_),
    .C(_427_),
    .Y(_428_)
);

NOR2X1 _1063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_356_),
    .B(_428_),
    .Y(_429_)
);

NOR2X1 _1064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[22]),
    .B(_429_),
    .Y(_430_)
);

NAND2X1 _1065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[22]),
    .B(_429_),
    .Y(_431_)
);

NAND2X1 _1066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_108__bF$buf1),
    .B(_431_),
    .Y(_432_)
);

OAI21X1 _1067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_432_),
    .B(_430_),
    .C(_424_),
    .Y(_486_[22])
);

NOR2X1 _1068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[21]),
    .B(_108__bF$buf0),
    .Y(_433_)
);

OR2X2 _1069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_431_),
    .B(mvect[23]),
    .Y(_434_)
);

AOI21X1 _1070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[23]),
    .B(_431_),
    .C(CSR_Ret_bF$buf0),
    .Y(_435_)
);

AOI21X1 _1071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_435_),
    .B(_434_),
    .C(_433_),
    .Y(_486_[23])
);

NAND2X1 _1072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[22]),
    .B(CSR_Ret_bF$buf5),
    .Y(_436_)
);

NAND2X1 _1073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[22]),
    .B(mvect[23]),
    .Y(_437_)
);

NOR3X1 _1074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_356_),
    .B(_437_),
    .C(_428_),
    .Y(_438_)
);

NOR2X1 _1075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[24]),
    .B(_438_),
    .Y(_439_)
);

INVX1 _1076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_438_),
    .Y(_440_)
);

OAI21X1 _1077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_440_),
    .B(_216_),
    .C(_108__bF$buf4),
    .Y(_441_)
);

OAI21X1 _1078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_441_),
    .B(_439_),
    .C(_436_),
    .Y(_486_[24])
);

NAND2X1 _1079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[23]),
    .B(CSR_Ret_bF$buf4),
    .Y(_442_)
);

AOI21X1 _1080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[24]),
    .B(_438_),
    .C(mvect[25]),
    .Y(_443_)
);

NAND2X1 _1081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[24]),
    .B(mvect[25]),
    .Y(_444_)
);

OAI21X1 _1082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_440_),
    .B(_444_),
    .C(_108__bF$buf3),
    .Y(_445_)
);

OAI21X1 _1083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_445_),
    .B(_443_),
    .C(_442_),
    .Y(_486_[25])
);

INVX1 _1084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_444_),
    .Y(_446_)
);

AOI21X1 _1085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_446_),
    .B(_438_),
    .C(mvect[26]),
    .Y(_447_)
);

NAND3X1 _1086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[26]),
    .B(_446_),
    .C(_438_),
    .Y(_448_)
);

NAND2X1 _1087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_108__bF$buf2),
    .B(_448_),
    .Y(_449_)
);

NAND2X1 _1088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[24]),
    .B(CSR_Ret_bF$buf3),
    .Y(_450_)
);

OAI21X1 _1089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_449_),
    .B(_447_),
    .C(_450_),
    .Y(_486_[26])
);

NAND3X1 _1090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_222_),
    .B(_108__bF$buf1),
    .C(_448_),
    .Y(_451_)
);

NOR2X1 _1091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[25]),
    .B(_108__bF$buf0),
    .Y(_452_)
);

NAND2X1 _1092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[26]),
    .B(mvect[27]),
    .Y(_453_)
);

NOR2X1 _1093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_444_),
    .B(_453_),
    .Y(_454_)
);

AND2X2 _1094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_454_),
    .B(_108__bF$buf4),
    .Y(_455_)
);

AOI21X1 _1095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_455_),
    .B(_438_),
    .C(_452_),
    .Y(_456_)
);

AND2X2 _1096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_451_),
    .B(_456_),
    .Y(_486_[27])
);

NAND2X1 _1097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[26]),
    .B(CSR_Ret_bF$buf2),
    .Y(_457_)
);

NOR3X1 _1098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_437_),
    .B(_444_),
    .C(_453_),
    .Y(_458_)
);

INVX1 _1099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_458_),
    .Y(_459_)
);

NOR3X1 _1100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_356_),
    .B(_459_),
    .C(_428_),
    .Y(_460_)
);

NOR2X1 _1101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[28]),
    .B(_460_),
    .Y(_461_)
);

NOR3X1 _1102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_368_),
    .B(_389_),
    .C(_422_),
    .Y(_462_)
);

NAND3X1 _1103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_351_),
    .B(_458_),
    .C(_462_),
    .Y(_463_)
);

OAI21X1 _1104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_463_),
    .B(_224_),
    .C(_108__bF$buf3),
    .Y(_464_)
);

OAI21X1 _1105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_464_),
    .B(_461_),
    .C(_457_),
    .Y(_486_[28])
);

NOR2X1 _1106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[27]),
    .B(_108__bF$buf2),
    .Y(_465_)
);

NAND2X1 _1107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[28]),
    .B(_460_),
    .Y(_466_)
);

OR2X2 _1108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_466_),
    .B(mvect[29]),
    .Y(_467_)
);

AOI21X1 _1109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[29]),
    .B(_466_),
    .C(CSR_Ret_bF$buf1),
    .Y(_468_)
);

AOI21X1 _1110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_468_),
    .B(_467_),
    .C(_465_),
    .Y(_486_[29])
);

INVX1 _1111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[28]),
    .Y(_469_)
);

NAND2X1 _1112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[28]),
    .B(mvect[29]),
    .Y(_470_)
);

NOR3X1 _1113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_),
    .B(_470_),
    .C(_157_),
    .Y(_471_)
);

NAND3X1 _1114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_350_),
    .B(_458_),
    .C(_471_),
    .Y(_472_)
);

OAI21X1 _1115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_472_),
    .B(_428_),
    .C(mvect[30]),
    .Y(_473_)
);

INVX1 _1116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_473_),
    .Y(_474_)
);

NOR2X1 _1117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_428_),
    .B(_472_),
    .Y(_475_)
);

AND2X2 _1118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_475_),
    .B(_228_),
    .Y(_476_)
);

OAI21X1 _1119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_476_),
    .B(_474_),
    .C(_108__bF$buf1),
    .Y(_477_)
);

OAI21X1 _1120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_469_),
    .B(_108__bF$buf0),
    .C(_477_),
    .Y(_486_[30])
);

INVX1 _1121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_470_),
    .Y(_478_)
);

NAND2X1 _1122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[30]),
    .B(_478_),
    .Y(_479_)
);

INVX1 _1123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_479_),
    .Y(_480_)
);

AOI21X1 _1124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_480_),
    .B(_460_),
    .C(_230_),
    .Y(_481_)
);

NOR3X1 _1125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[31]),
    .B(_479_),
    .C(_463_),
    .Y(_482_)
);

OAI21X1 _1126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_482_),
    .B(_481_),
    .C(_108__bF$buf4),
    .Y(_483_)
);

NAND2X1 _1127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[29]),
    .B(CSR_Ret_bF$buf0),
    .Y(_484_)
);

NAND2X1 _1128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_484_),
    .B(_483_),
    .Y(_486_[31])
);

BUFX2 _1129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_485_),
    .Y(CSR_IRQ)
);

BUFX2 _1130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .Y(CSR_PCaddr[0])
);

BUFX2 _1131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(gnd),
    .Y(CSR_PCaddr[1])
);

BUFX2 _1132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[2]),
    .Y(CSR_PCaddr[2])
);

BUFX2 _1133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[3]),
    .Y(CSR_PCaddr[3])
);

BUFX2 _1134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[4]),
    .Y(CSR_PCaddr[4])
);

BUFX2 _1135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[5]),
    .Y(CSR_PCaddr[5])
);

BUFX2 _1136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[6]),
    .Y(CSR_PCaddr[6])
);

BUFX2 _1137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[7]),
    .Y(CSR_PCaddr[7])
);

BUFX2 _1138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[8]),
    .Y(CSR_PCaddr[8])
);

BUFX2 _1139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[9]),
    .Y(CSR_PCaddr[9])
);

BUFX2 _1140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[10]),
    .Y(CSR_PCaddr[10])
);

BUFX2 _1141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[11]),
    .Y(CSR_PCaddr[11])
);

BUFX2 _1142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[12]),
    .Y(CSR_PCaddr[12])
);

BUFX2 _1143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[13]),
    .Y(CSR_PCaddr[13])
);

BUFX2 _1144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[14]),
    .Y(CSR_PCaddr[14])
);

BUFX2 _1145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[15]),
    .Y(CSR_PCaddr[15])
);

BUFX2 _1146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[16]),
    .Y(CSR_PCaddr[16])
);

BUFX2 _1147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[17]),
    .Y(CSR_PCaddr[17])
);

BUFX2 _1148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[18]),
    .Y(CSR_PCaddr[18])
);

BUFX2 _1149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[19]),
    .Y(CSR_PCaddr[19])
);

BUFX2 _1150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[20]),
    .Y(CSR_PCaddr[20])
);

BUFX2 _1151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[21]),
    .Y(CSR_PCaddr[21])
);

BUFX2 _1152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[22]),
    .Y(CSR_PCaddr[22])
);

BUFX2 _1153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[23]),
    .Y(CSR_PCaddr[23])
);

BUFX2 _1154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[24]),
    .Y(CSR_PCaddr[24])
);

BUFX2 _1155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[25]),
    .Y(CSR_PCaddr[25])
);

BUFX2 _1156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[26]),
    .Y(CSR_PCaddr[26])
);

BUFX2 _1157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[27]),
    .Y(CSR_PCaddr[27])
);

BUFX2 _1158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[28]),
    .Y(CSR_PCaddr[28])
);

BUFX2 _1159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[29]),
    .Y(CSR_PCaddr[29])
);

BUFX2 _1160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[30]),
    .Y(CSR_PCaddr[30])
);

BUFX2 _1161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_[31]),
    .Y(CSR_PCaddr[31])
);

BUFX2 _1162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[0]),
    .Y(CSR_data[0])
);

BUFX2 _1163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[1]),
    .Y(CSR_data[1])
);

BUFX2 _1164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[2]),
    .Y(CSR_data[2])
);

BUFX2 _1165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[3]),
    .Y(CSR_data[3])
);

BUFX2 _1166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[4]),
    .Y(CSR_data[4])
);

BUFX2 _1167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[5]),
    .Y(CSR_data[5])
);

BUFX2 _1168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[6]),
    .Y(CSR_data[6])
);

BUFX2 _1169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[7]),
    .Y(CSR_data[7])
);

BUFX2 _1170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[8]),
    .Y(CSR_data[8])
);

BUFX2 _1171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[9]),
    .Y(CSR_data[9])
);

BUFX2 _1172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[10]),
    .Y(CSR_data[10])
);

BUFX2 _1173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[11]),
    .Y(CSR_data[11])
);

BUFX2 _1174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[12]),
    .Y(CSR_data[12])
);

BUFX2 _1175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[13]),
    .Y(CSR_data[13])
);

BUFX2 _1176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[14]),
    .Y(CSR_data[14])
);

BUFX2 _1177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[15]),
    .Y(CSR_data[15])
);

BUFX2 _1178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[16]),
    .Y(CSR_data[16])
);

BUFX2 _1179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[17]),
    .Y(CSR_data[17])
);

BUFX2 _1180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[18]),
    .Y(CSR_data[18])
);

BUFX2 _1181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[19]),
    .Y(CSR_data[19])
);

BUFX2 _1182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[20]),
    .Y(CSR_data[20])
);

BUFX2 _1183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[21]),
    .Y(CSR_data[21])
);

BUFX2 _1184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[22]),
    .Y(CSR_data[22])
);

BUFX2 _1185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[23]),
    .Y(CSR_data[23])
);

BUFX2 _1186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[24]),
    .Y(CSR_data[24])
);

BUFX2 _1187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[25]),
    .Y(CSR_data[25])
);

BUFX2 _1188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[26]),
    .Y(CSR_data[26])
);

BUFX2 _1189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[27]),
    .Y(CSR_data[27])
);

BUFX2 _1190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[28]),
    .Y(CSR_data[28])
);

BUFX2 _1191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[29]),
    .Y(CSR_data[29])
);

BUFX2 _1192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[30]),
    .Y(CSR_data[30])
);

BUFX2 _1193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_[31]),
    .Y(CSR_data[31])
);

DFFPOSX1 _1194_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_21_[0]),
    .Q(mepc[0])
);

DFFPOSX1 _1195_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_21_[1]),
    .Q(mepc[1])
);

DFFPOSX1 _1196_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_21_[2]),
    .Q(mepc[2])
);

DFFPOSX1 _1197_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_21_[3]),
    .Q(mepc[3])
);

DFFPOSX1 _1198_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_21_[4]),
    .Q(mepc[4])
);

DFFPOSX1 _1199_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_21_[5]),
    .Q(mepc[5])
);

DFFPOSX1 _1200_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_21_[6]),
    .Q(mepc[6])
);

DFFPOSX1 _1201_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_21_[7]),
    .Q(mepc[7])
);

DFFPOSX1 _1202_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_21_[8]),
    .Q(mepc[8])
);

DFFPOSX1 _1203_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_21_[9]),
    .Q(mepc[9])
);

DFFPOSX1 _1204_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_21_[10]),
    .Q(mepc[10])
);

DFFPOSX1 _1205_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_21_[11]),
    .Q(mepc[11])
);

DFFPOSX1 _1206_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_21_[12]),
    .Q(mepc[12])
);

DFFPOSX1 _1207_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_21_[13]),
    .Q(mepc[13])
);

DFFPOSX1 _1208_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_21_[14]),
    .Q(mepc[14])
);

DFFPOSX1 _1209_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_21_[15]),
    .Q(mepc[15])
);

DFFPOSX1 _1210_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_21_[16]),
    .Q(mepc[16])
);

DFFPOSX1 _1211_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_21_[17]),
    .Q(mepc[17])
);

DFFPOSX1 _1212_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_21_[18]),
    .Q(mepc[18])
);

DFFPOSX1 _1213_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_21_[19]),
    .Q(mepc[19])
);

DFFPOSX1 _1214_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_21_[20]),
    .Q(mepc[20])
);

DFFPOSX1 _1215_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_21_[21]),
    .Q(mepc[21])
);

DFFPOSX1 _1216_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_21_[22]),
    .Q(mepc[22])
);

DFFPOSX1 _1217_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_21_[23]),
    .Q(mepc[23])
);

DFFPOSX1 _1218_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_21_[24]),
    .Q(mepc[24])
);

DFFPOSX1 _1219_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_21_[25]),
    .Q(mepc[25])
);

DFFPOSX1 _1220_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_21_[26]),
    .Q(mepc[26])
);

DFFPOSX1 _1221_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_21_[27]),
    .Q(mepc[27])
);

DFFPOSX1 _1222_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_21_[28]),
    .Q(mepc[28])
);

DFFPOSX1 _1223_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_21_[29]),
    .Q(mepc[29])
);

DFFPOSX1 _1224_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(Extern_IRQ),
    .Q(meta_irq)
);

DFFPOSX1 _1225_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(meta_irq),
    .Q(mip)
);

DFFPOSX1 _1226_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_14_),
    .Q(mie)
);

DFFPOSX1 _1227_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_07_[0]),
    .Q(mvect[0])
);

DFFPOSX1 _1228_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_07_[1]),
    .Q(mvect[1])
);

DFFPOSX1 _1229_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_07_[2]),
    .Q(mvect[2])
);

DFFPOSX1 _1230_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_07_[3]),
    .Q(mvect[3])
);

DFFPOSX1 _1231_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_07_[4]),
    .Q(mvect[4])
);

DFFPOSX1 _1232_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_07_[5]),
    .Q(mvect[5])
);

DFFPOSX1 _1233_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_07_[6]),
    .Q(mvect[6])
);

DFFPOSX1 _1234_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_07_[7]),
    .Q(mvect[7])
);

DFFPOSX1 _1235_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_07_[8]),
    .Q(mvect[8])
);

DFFPOSX1 _1236_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_07_[9]),
    .Q(mvect[9])
);

DFFPOSX1 _1237_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_07_[10]),
    .Q(mvect[10])
);

DFFPOSX1 _1238_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_07_[11]),
    .Q(mvect[11])
);

DFFPOSX1 _1239_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_07_[12]),
    .Q(mvect[12])
);

DFFPOSX1 _1240_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_07_[13]),
    .Q(mvect[13])
);

DFFPOSX1 _1241_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_07_[14]),
    .Q(mvect[14])
);

DFFPOSX1 _1242_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_07_[15]),
    .Q(mvect[15])
);

DFFPOSX1 _1243_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_07_[16]),
    .Q(mvect[16])
);

DFFPOSX1 _1244_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_07_[17]),
    .Q(mvect[17])
);

DFFPOSX1 _1245_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_07_[18]),
    .Q(mvect[18])
);

DFFPOSX1 _1246_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_07_[19]),
    .Q(mvect[19])
);

DFFPOSX1 _1247_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_07_[20]),
    .Q(mvect[20])
);

DFFPOSX1 _1248_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_07_[21]),
    .Q(mvect[21])
);

DFFPOSX1 _1249_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_07_[22]),
    .Q(mvect[22])
);

DFFPOSX1 _1250_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_07_[23]),
    .Q(mvect[23])
);

DFFPOSX1 _1251_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_07_[24]),
    .Q(mvect[24])
);

DFFPOSX1 _1252_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_07_[25]),
    .Q(mvect[25])
);

DFFPOSX1 _1253_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_07_[26]),
    .Q(mvect[26])
);

DFFPOSX1 _1254_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_07_[27]),
    .Q(mvect[27])
);

DFFPOSX1 _1255_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_07_[28]),
    .Q(mvect[28])
);

DFFPOSX1 _1256_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_07_[29]),
    .Q(mvect[29])
);

DFFPOSX1 _1257_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_07_[30]),
    .Q(mvect[30])
);

DFFPOSX1 _1258_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_07_[31]),
    .Q(mvect[31])
);

DFFPOSX1 _1259_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_33_[0]),
    .Q(mstatus[0])
);

DFFPOSX1 _1260_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_33_[1]),
    .Q(mstatus[1])
);

DFFPOSX1 _1261_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_28_[0]),
    .Q(mcause[0])
);

DFFPOSX1 _1262_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_28_[1]),
    .Q(mcause[1])
);

DFFPOSX1 _1263_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_28_[2]),
    .Q(mcause[2])
);

DFFPOSX1 _1264_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_28_[3]),
    .Q(mcause[3])
);

DFFPOSX1 _1265_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_28_[4]),
    .Q(mcause[4])
);

DFFPOSX1 _1266_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_28_[5]),
    .Q(mcause[5])
);

DFFPOSX1 _1267_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_28_[6]),
    .Q(mcause[6])
);

DFFPOSX1 _1268_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_28_[7]),
    .Q(mcause[7])
);

DFFPOSX1 _1269_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_28_[8]),
    .Q(mcause[8])
);

DFFPOSX1 _1270_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_28_[9]),
    .Q(mcause[9])
);

DFFPOSX1 _1271_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_28_[10]),
    .Q(mcause[10])
);

DFFPOSX1 _1272_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_28_[11]),
    .Q(mcause[11])
);

DFFPOSX1 _1273_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_28_[12]),
    .Q(mcause[12])
);

DFFPOSX1 _1274_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_28_[13]),
    .Q(mcause[13])
);

DFFPOSX1 _1275_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_28_[14]),
    .Q(mcause[14])
);

DFFPOSX1 _1276_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_28_[15]),
    .Q(mcause[15])
);

DFFPOSX1 _1277_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_28_[16]),
    .Q(mcause[16])
);

DFFPOSX1 _1278_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_28_[17]),
    .Q(mcause[17])
);

DFFPOSX1 _1279_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_28_[18]),
    .Q(mcause[18])
);

DFFPOSX1 _1280_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_28_[19]),
    .Q(mcause[19])
);

DFFPOSX1 _1281_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_28_[20]),
    .Q(mcause[20])
);

DFFPOSX1 _1282_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_28_[21]),
    .Q(mcause[21])
);

DFFPOSX1 _1283_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_28_[22]),
    .Q(mcause[22])
);

DFFPOSX1 _1284_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(_28_[23]),
    .Q(mcause[23])
);

DFFPOSX1 _1285_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_28_[24]),
    .Q(mcause[24])
);

DFFPOSX1 _1286_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_28_[25]),
    .Q(mcause[25])
);

DFFPOSX1 _1287_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_28_[26]),
    .Q(mcause[26])
);

DFFPOSX1 _1288_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_28_[27]),
    .Q(mcause[27])
);

DFFPOSX1 _1289_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_28_[28]),
    .Q(mcause[28])
);

DFFPOSX1 _1290_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_28_[29]),
    .Q(mcause[29])
);

DFFPOSX1 _1291_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_28_[30]),
    .Q(mcause[30])
);

DFFPOSX1 _1292_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_28_[31]),
    .Q(mcause[31])
);

INVX2 _488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[0]),
    .Y(_0_)
);

NOR2X1 _489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_addr[11]),
    .B(CSR_addr[10]),
    .Y(_1_)
);

NAND3X1 _490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_addr[9]),
    .B(CSR_addr[8]),
    .C(_1_),
    .Y(_2_)
);

INVX1 _491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_addr[7]),
    .Y(_3_)
);

NOR2X1 _492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_addr[5]),
    .B(CSR_addr[4]),
    .Y(_4_)
);

NAND3X1 _493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3_),
    .B(CSR_addr[6]),
    .C(_4_),
    .Y(_5_)
);

NOR2X1 _494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_),
    .B(_5_),
    .Y(_6_)
);

OR2X2 _495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_addr[3]),
    .B(CSR_addr[2]),
    .Y(_7_)
);

INVX1 _496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_addr[0]),
    .Y(_8_)
);

NAND2X1 _497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_addr[1]),
    .B(_8_),
    .Y(_9_)
);

NOR2X1 _498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7_),
    .B(_9_),
    .Y(_10_)
);

NAND2X1 _499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10_),
    .B(_6_),
    .Y(_11_)
);

INVX4 _500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11__bF$buf4),
    .Y(_12_)
);

NAND2X1 _501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[0]),
    .B(_12_),
    .Y(_13_)
);

NOR2X1 _502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_addr[7]),
    .B(CSR_addr[6]),
    .Y(_15_)
);

NAND2X1 _503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4_),
    .B(_15_),
    .Y(_16_)
);

NOR2X1 _504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_16_),
    .B(_2_),
    .Y(_17_)
);

INVX1 _505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_addr[1]),
    .Y(_18_)
);

NAND2X1 _506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_addr[0]),
    .B(_18_),
    .Y(_19_)
);

INVX1 _507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_addr[3]),
    .Y(_20_)
);

NAND2X1 _508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_addr[2]),
    .B(_20_),
    .Y(_22_)
);

NOR2X1 _509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_19_),
    .B(_22_),
    .Y(_23_)
);

AND2X2 _510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_17_),
    .B(_23_),
    .Y(_24_)
);

INVX1 _511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf4),
    .Y(_25_)
);

OAI21X1 _512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_),
    .B(_25_),
    .C(_13_),
    .Y(_487_[0])
);

INVX1 _513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[1]),
    .Y(_26_)
);

NAND2X1 _514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[1]),
    .B(_12_),
    .Y(_27_)
);

OAI21X1 _515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_26_),
    .B(_25_),
    .C(_27_),
    .Y(_487_[1])
);

INVX1 _516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[2]),
    .Y(_29_)
);

NOR2X1 _517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7_),
    .B(_19_),
    .Y(_30_)
);

AND2X2 _518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6_),
    .B(_30_),
    .Y(_31_)
);

AOI22X1 _519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf3),
    .B(mvect[2]),
    .C(mepc[0]),
    .D(_31__bF$buf4),
    .Y(_32_)
);

OAI21X1 _520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_29_),
    .B(_11__bF$buf3),
    .C(_32_),
    .Y(_487_[2])
);

INVX1 _521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mstatus[0]),
    .Y(_34_)
);

NOR2X1 _522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_addr[1]),
    .B(CSR_addr[0]),
    .Y(_35_)
);

INVX1 _523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_17_),
    .Y(_36_)
);

NOR2X1 _524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7_),
    .B(_36_),
    .Y(_37_)
);

NAND2X1 _525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_35_),
    .B(_37_),
    .Y(_38_)
);

NAND2X1 _526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[1]),
    .B(_31__bF$buf3),
    .Y(_39_)
);

AOI22X1 _527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[3]),
    .B(_24__bF$buf2),
    .C(_12_),
    .D(mcause[3]),
    .Y(_40_)
);

AND2X2 _528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_40_),
    .B(_39_),
    .Y(_41_)
);

OAI21X1 _529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_34_),
    .B(_38_),
    .C(_41_),
    .Y(_487_[3])
);

INVX1 _530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[4]),
    .Y(_42_)
);

AOI22X1 _531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf1),
    .B(mvect[4]),
    .C(mepc[2]),
    .D(_31__bF$buf2),
    .Y(_43_)
);

OAI21X1 _532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_42_),
    .B(_11__bF$buf2),
    .C(_43_),
    .Y(_487_[4])
);

INVX1 _533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[5]),
    .Y(_44_)
);

AOI22X1 _534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf0),
    .B(mvect[5]),
    .C(mepc[3]),
    .D(_31__bF$buf1),
    .Y(_45_)
);

OAI21X1 _535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_44_),
    .B(_11__bF$buf1),
    .C(_45_),
    .Y(_487_[5])
);

INVX1 _536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[6]),
    .Y(_46_)
);

AOI22X1 _537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf4),
    .B(mvect[6]),
    .C(mepc[4]),
    .D(_31__bF$buf0),
    .Y(_47_)
);

OAI21X1 _538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_46_),
    .B(_11__bF$buf0),
    .C(_47_),
    .Y(_487_[6])
);

INVX1 _539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mstatus[1]),
    .Y(_48_)
);

NAND2X1 _540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[5]),
    .B(_31__bF$buf4),
    .Y(_49_)
);

AOI22X1 _541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[7]),
    .B(_24__bF$buf3),
    .C(_12_),
    .D(mcause[7]),
    .Y(_50_)
);

AND2X2 _542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_50_),
    .B(_49_),
    .Y(_51_)
);

OAI21X1 _543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_48_),
    .B(_38_),
    .C(_51_),
    .Y(_487_[7])
);

AND2X2 _544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_17_),
    .B(_30_),
    .Y(_52_)
);

AOI21X1 _545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[8]),
    .B(_24__bF$buf2),
    .C(_52_),
    .Y(_53_)
);

AOI22X1 _546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[6]),
    .B(_31__bF$buf3),
    .C(_12_),
    .D(mcause[8]),
    .Y(_54_)
);

NAND2X1 _547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_53_),
    .B(_54_),
    .Y(_487_[8])
);

INVX1 _548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[9]),
    .Y(_55_)
);

AOI22X1 _549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf1),
    .B(mvect[9]),
    .C(mepc[7]),
    .D(_31__bF$buf2),
    .Y(_56_)
);

OAI21X1 _550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_55_),
    .B(_11__bF$buf4),
    .C(_56_),
    .Y(_487_[9])
);

INVX1 _551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[10]),
    .Y(_57_)
);

AOI22X1 _552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf0),
    .B(mvect[10]),
    .C(mepc[8]),
    .D(_31__bF$buf1),
    .Y(_58_)
);

OAI21X1 _553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_57_),
    .B(_11__bF$buf3),
    .C(_58_),
    .Y(_487_[10])
);

INVX1 _554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mip),
    .Y(_59_)
);

INVX1 _555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_35_),
    .Y(_60_)
);

OR2X2 _556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_60_),
    .B(_22_),
    .Y(_61_)
);

NOR2X1 _557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_59_),
    .B(_61_),
    .Y(_62_)
);

AOI22X1 _558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6_),
    .B(_62_),
    .C(_37_),
    .D(_35_),
    .Y(_63_)
);

NOR2X1 _559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_61_),
    .B(_36_),
    .Y(_64_)
);

AOI22X1 _560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[11]),
    .B(_12_),
    .C(_64_),
    .D(mie),
    .Y(_65_)
);

AOI22X1 _561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf4),
    .B(mvect[11]),
    .C(mepc[9]),
    .D(_31__bF$buf0),
    .Y(_66_)
);

NAND3X1 _562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_66_),
    .B(_63_),
    .C(_65_),
    .Y(_487_[11])
);

NAND2X1 _563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[10]),
    .B(_31__bF$buf4),
    .Y(_67_)
);

AOI22X1 _564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[12]),
    .B(_24__bF$buf3),
    .C(_12_),
    .D(mcause[12]),
    .Y(_68_)
);

NAND3X1 _565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_38_),
    .B(_67_),
    .C(_68_),
    .Y(_487_[12])
);

INVX1 _566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[13]),
    .Y(_69_)
);

AOI22X1 _567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf2),
    .B(mvect[13]),
    .C(mepc[11]),
    .D(_31__bF$buf3),
    .Y(_70_)
);

OAI21X1 _568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_69_),
    .B(_11__bF$buf2),
    .C(_70_),
    .Y(_487_[13])
);

INVX1 _569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[14]),
    .Y(_71_)
);

AOI22X1 _570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf1),
    .B(mvect[14]),
    .C(mepc[12]),
    .D(_31__bF$buf2),
    .Y(_72_)
);

OAI21X1 _571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_71_),
    .B(_11__bF$buf1),
    .C(_72_),
    .Y(_487_[14])
);

INVX1 _572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[15]),
    .Y(_73_)
);

AOI22X1 _573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf0),
    .B(mvect[15]),
    .C(mepc[13]),
    .D(_31__bF$buf1),
    .Y(_74_)
);

OAI21X1 _574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73_),
    .B(_11__bF$buf0),
    .C(_74_),
    .Y(_487_[15])
);

INVX1 _575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[16]),
    .Y(_75_)
);

AOI22X1 _576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf4),
    .B(mvect[16]),
    .C(mepc[14]),
    .D(_31__bF$buf0),
    .Y(_76_)
);

OAI21X1 _577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_75_),
    .B(_11__bF$buf4),
    .C(_76_),
    .Y(_487_[16])
);

INVX1 _578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[17]),
    .Y(_77_)
);

AOI22X1 _579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf3),
    .B(mvect[17]),
    .C(mepc[15]),
    .D(_31__bF$buf4),
    .Y(_78_)
);

OAI21X1 _580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_77_),
    .B(_11__bF$buf3),
    .C(_78_),
    .Y(_487_[17])
);

INVX1 _581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[18]),
    .Y(_79_)
);

AOI22X1 _582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf2),
    .B(mvect[18]),
    .C(mepc[16]),
    .D(_31__bF$buf3),
    .Y(_80_)
);

OAI21X1 _583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_79_),
    .B(_11__bF$buf2),
    .C(_80_),
    .Y(_487_[18])
);

INVX1 _584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[19]),
    .Y(_81_)
);

AOI22X1 _585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf1),
    .B(mvect[19]),
    .C(mepc[17]),
    .D(_31__bF$buf2),
    .Y(_82_)
);

OAI21X1 _586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_81_),
    .B(_11__bF$buf1),
    .C(_82_),
    .Y(_487_[19])
);

INVX1 _587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[20]),
    .Y(_83_)
);

AOI22X1 _588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf0),
    .B(mvect[20]),
    .C(mepc[18]),
    .D(_31__bF$buf1),
    .Y(_84_)
);

OAI21X1 _589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_83_),
    .B(_11__bF$buf0),
    .C(_84_),
    .Y(_487_[20])
);

INVX1 _590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[21]),
    .Y(_85_)
);

AOI22X1 _591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf4),
    .B(mvect[21]),
    .C(mepc[19]),
    .D(_31__bF$buf0),
    .Y(_86_)
);

OAI21X1 _592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(_11__bF$buf4),
    .C(_86_),
    .Y(_487_[21])
);

INVX1 _593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[22]),
    .Y(_87_)
);

AOI22X1 _594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf3),
    .B(mvect[22]),
    .C(mepc[20]),
    .D(_31__bF$buf4),
    .Y(_88_)
);

OAI21X1 _595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_87_),
    .B(_11__bF$buf3),
    .C(_88_),
    .Y(_487_[22])
);

INVX1 _596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[23]),
    .Y(_89_)
);

AOI22X1 _597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf2),
    .B(mvect[23]),
    .C(mepc[21]),
    .D(_31__bF$buf3),
    .Y(_90_)
);

OAI21X1 _598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_89_),
    .B(_11__bF$buf2),
    .C(_90_),
    .Y(_487_[23])
);

INVX1 _599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[24]),
    .Y(_91_)
);

AOI22X1 _600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf1),
    .B(mvect[24]),
    .C(mepc[22]),
    .D(_31__bF$buf2),
    .Y(_92_)
);

OAI21X1 _601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_91_),
    .B(_11__bF$buf1),
    .C(_92_),
    .Y(_487_[24])
);

INVX1 _602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[25]),
    .Y(_93_)
);

AOI22X1 _603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf0),
    .B(mvect[25]),
    .C(mepc[23]),
    .D(_31__bF$buf1),
    .Y(_94_)
);

OAI21X1 _604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_11__bF$buf0),
    .C(_94_),
    .Y(_487_[25])
);

INVX1 _605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[26]),
    .Y(_95_)
);

AOI22X1 _606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf4),
    .B(mvect[26]),
    .C(mepc[24]),
    .D(_31__bF$buf0),
    .Y(_96_)
);

OAI21X1 _607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_95_),
    .B(_11__bF$buf4),
    .C(_96_),
    .Y(_487_[26])
);

INVX1 _608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[27]),
    .Y(_97_)
);

AOI22X1 _609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf3),
    .B(mvect[27]),
    .C(mepc[25]),
    .D(_31__bF$buf4),
    .Y(_98_)
);

OAI21X1 _610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_97_),
    .B(_11__bF$buf3),
    .C(_98_),
    .Y(_487_[27])
);

INVX1 _611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[28]),
    .Y(_99_)
);

AOI22X1 _612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf2),
    .B(mvect[28]),
    .C(mepc[26]),
    .D(_31__bF$buf3),
    .Y(_100_)
);

OAI21X1 _613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_99_),
    .B(_11__bF$buf2),
    .C(_100_),
    .Y(_487_[28])
);

INVX1 _614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[29]),
    .Y(_101_)
);

AOI22X1 _615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf1),
    .B(mvect[29]),
    .C(mepc[27]),
    .D(_31__bF$buf2),
    .Y(_102_)
);

OAI21X1 _616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_101_),
    .B(_11__bF$buf1),
    .C(_102_),
    .Y(_487_[29])
);

AOI21X1 _617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[30]),
    .B(_24__bF$buf0),
    .C(_52_),
    .Y(_103_)
);

AOI22X1 _618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[28]),
    .B(_31__bF$buf1),
    .C(_12_),
    .D(mcause[30]),
    .Y(_104_)
);

NAND2X1 _619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_103_),
    .B(_104_),
    .Y(_487_[30])
);

INVX1 _620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[31]),
    .Y(_105_)
);

AOI22X1 _621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24__bF$buf4),
    .B(mvect[31]),
    .C(mepc[29]),
    .D(_31__bF$buf0),
    .Y(_106_)
);

OAI21X1 _622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_105_),
    .B(_11__bF$buf0),
    .C(_106_),
    .Y(_487_[31])
);

NAND2X1 _623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_mcause[0]),
    .B(CSR_Wen_traps_bF$buf5),
    .Y(_107_)
);

INVX8 _624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Ret_bF$buf5),
    .Y(_108_)
);

NAND2X1 _625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen),
    .B(_108__bF$buf3),
    .Y(_109_)
);

NOR2X1 _626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_109_),
    .B(_11__bF$buf4),
    .Y(_110_)
);

NOR2X1 _627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[0]),
    .B(_110_),
    .Y(_111_)
);

INVX8 _628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf4),
    .Y(_112_)
);

INVX1 _629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_109_),
    .Y(_113_)
);

NAND2X1 _630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_113_),
    .B(_12_),
    .Y(_114_)
);

OAI21X1 _631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf6),
    .B(CSR_Wdata[0]),
    .C(_112__bF$buf6),
    .Y(_115_)
);

OAI21X1 _632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_115_),
    .B(_111_),
    .C(_107_),
    .Y(_28_[0])
);

NAND2X1 _633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf3),
    .B(CSR_mcause[1]),
    .Y(_116_)
);

NOR2X1 _634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[1]),
    .B(_110_),
    .Y(_117_)
);

OAI21X1 _635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf5),
    .B(CSR_Wdata[1]),
    .C(_112__bF$buf5),
    .Y(_118_)
);

OAI21X1 _636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_118_),
    .B(_117_),
    .C(_116_),
    .Y(_28_[1])
);

NAND2X1 _637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf2),
    .B(CSR_mcause[2]),
    .Y(_119_)
);

OAI21X1 _638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11__bF$buf3),
    .B(_109_),
    .C(_29_),
    .Y(_120_)
);

OAI21X1 _639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf4),
    .B(CSR_Wdata[2]),
    .C(_120_),
    .Y(_121_)
);

OAI21X1 _640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_121_),
    .B(CSR_Wen_traps_bF$buf1),
    .C(_119_),
    .Y(_28_[2])
);

NAND2X1 _641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf0),
    .B(CSR_mcause[3]),
    .Y(_122_)
);

NOR2X1 _642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[3]),
    .B(_110_),
    .Y(_123_)
);

OAI21X1 _643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf3),
    .B(CSR_Wdata[3]),
    .C(_112__bF$buf4),
    .Y(_124_)
);

OAI21X1 _644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_124_),
    .B(_123_),
    .C(_122_),
    .Y(_28_[3])
);

OAI21X1 _645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf2),
    .B(CSR_Wdata[4]),
    .C(_112__bF$buf3),
    .Y(_125_)
);

AOI21X1 _646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_42_),
    .B(_114__bF$buf1),
    .C(_125_),
    .Y(_28_[4])
);

OAI21X1 _647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf0),
    .B(CSR_Wdata[5]),
    .C(_112__bF$buf2),
    .Y(_126_)
);

AOI21X1 _648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_44_),
    .B(_114__bF$buf6),
    .C(_126_),
    .Y(_28_[5])
);

OAI21X1 _649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf5),
    .B(CSR_Wdata[6]),
    .C(_112__bF$buf1),
    .Y(_127_)
);

AOI21X1 _650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_46_),
    .B(_114__bF$buf4),
    .C(_127_),
    .Y(_28_[6])
);

NOR2X1 _651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[7]),
    .B(_110_),
    .Y(_128_)
);

OAI21X1 _652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf3),
    .B(CSR_Wdata[7]),
    .C(_112__bF$buf0),
    .Y(_129_)
);

NOR2X1 _653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_128_),
    .B(_129_),
    .Y(_28_[7])
);

NOR2X1 _654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[8]),
    .B(_110_),
    .Y(_130_)
);

OAI21X1 _655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf2),
    .B(CSR_Wdata[8]),
    .C(_112__bF$buf6),
    .Y(_131_)
);

NOR2X1 _656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_130_),
    .B(_131_),
    .Y(_28_[8])
);

OAI21X1 _657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf1),
    .B(CSR_Wdata[9]),
    .C(_112__bF$buf5),
    .Y(_132_)
);

AOI21X1 _658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_55_),
    .B(_114__bF$buf0),
    .C(_132_),
    .Y(_28_[9])
);

OAI21X1 _659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf6),
    .B(CSR_Wdata[10]),
    .C(_112__bF$buf4),
    .Y(_133_)
);

AOI21X1 _660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_57_),
    .B(_114__bF$buf5),
    .C(_133_),
    .Y(_28_[10])
);

NOR2X1 _661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[11]),
    .B(_110_),
    .Y(_134_)
);

OAI21X1 _662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf4),
    .B(CSR_Wdata[11]),
    .C(_112__bF$buf3),
    .Y(_135_)
);

NOR2X1 _663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_134_),
    .B(_135_),
    .Y(_28_[11])
);

NOR2X1 _664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[12]),
    .B(_110_),
    .Y(_136_)
);

OAI21X1 _665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf3),
    .B(CSR_Wdata[12]),
    .C(_112__bF$buf2),
    .Y(_137_)
);

NOR2X1 _666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_136_),
    .B(_137_),
    .Y(_28_[12])
);

OAI21X1 _667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf2),
    .B(CSR_Wdata[13]),
    .C(_112__bF$buf1),
    .Y(_138_)
);

AOI21X1 _668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_69_),
    .B(_114__bF$buf1),
    .C(_138_),
    .Y(_28_[13])
);

OAI21X1 _669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf0),
    .B(CSR_Wdata[14]),
    .C(_112__bF$buf0),
    .Y(_139_)
);

AOI21X1 _670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_71_),
    .B(_114__bF$buf6),
    .C(_139_),
    .Y(_28_[14])
);

OAI21X1 _671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf5),
    .B(CSR_Wdata[15]),
    .C(_112__bF$buf6),
    .Y(_140_)
);

AOI21X1 _672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73_),
    .B(_114__bF$buf4),
    .C(_140_),
    .Y(_28_[15])
);

OAI21X1 _673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf3),
    .B(CSR_Wdata[16]),
    .C(_112__bF$buf5),
    .Y(_141_)
);

AOI21X1 _674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_75_),
    .B(_114__bF$buf2),
    .C(_141_),
    .Y(_28_[16])
);

OAI21X1 _675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf1),
    .B(CSR_Wdata[17]),
    .C(_112__bF$buf4),
    .Y(_142_)
);

AOI21X1 _676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_77_),
    .B(_114__bF$buf0),
    .C(_142_),
    .Y(_28_[17])
);

OAI21X1 _677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf6),
    .B(CSR_Wdata[18]),
    .C(_112__bF$buf3),
    .Y(_143_)
);

AOI21X1 _678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_79_),
    .B(_114__bF$buf5),
    .C(_143_),
    .Y(_28_[18])
);

OAI21X1 _679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf4),
    .B(CSR_Wdata[19]),
    .C(_112__bF$buf2),
    .Y(_144_)
);

AOI21X1 _680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_81_),
    .B(_114__bF$buf3),
    .C(_144_),
    .Y(_28_[19])
);

OAI21X1 _681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf2),
    .B(CSR_Wdata[20]),
    .C(_112__bF$buf1),
    .Y(_145_)
);

AOI21X1 _682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_83_),
    .B(_114__bF$buf1),
    .C(_145_),
    .Y(_28_[20])
);

OAI21X1 _683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf0),
    .B(CSR_Wdata[21]),
    .C(_112__bF$buf0),
    .Y(_146_)
);

AOI21X1 _684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(_114__bF$buf6),
    .C(_146_),
    .Y(_28_[21])
);

OAI21X1 _685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf5),
    .B(CSR_Wdata[22]),
    .C(_112__bF$buf6),
    .Y(_147_)
);

AOI21X1 _686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_87_),
    .B(_114__bF$buf4),
    .C(_147_),
    .Y(_28_[22])
);

OAI21X1 _687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf3),
    .B(CSR_Wdata[23]),
    .C(_112__bF$buf5),
    .Y(_148_)
);

AOI21X1 _688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_89_),
    .B(_114__bF$buf2),
    .C(_148_),
    .Y(_28_[23])
);

OAI21X1 _689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf1),
    .B(CSR_Wdata[24]),
    .C(_112__bF$buf4),
    .Y(_149_)
);

AOI21X1 _690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_91_),
    .B(_114__bF$buf0),
    .C(_149_),
    .Y(_28_[24])
);

OAI21X1 _691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf6),
    .B(CSR_Wdata[25]),
    .C(_112__bF$buf3),
    .Y(_150_)
);

AOI21X1 _692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_114__bF$buf5),
    .C(_150_),
    .Y(_28_[25])
);

OAI21X1 _693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf4),
    .B(CSR_Wdata[26]),
    .C(_112__bF$buf2),
    .Y(_151_)
);

AOI21X1 _694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_95_),
    .B(_114__bF$buf3),
    .C(_151_),
    .Y(_28_[26])
);

OAI21X1 _695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf2),
    .B(CSR_Wdata[27]),
    .C(_112__bF$buf1),
    .Y(_152_)
);

AOI21X1 _696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_97_),
    .B(_114__bF$buf1),
    .C(_152_),
    .Y(_28_[27])
);

OAI21X1 _697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf0),
    .B(CSR_Wdata[28]),
    .C(_112__bF$buf0),
    .Y(_153_)
);

AOI21X1 _698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_99_),
    .B(_114__bF$buf6),
    .C(_153_),
    .Y(_28_[28])
);

OAI21X1 _699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf5),
    .B(CSR_Wdata[29]),
    .C(_112__bF$buf6),
    .Y(_154_)
);

AOI21X1 _700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_101_),
    .B(_114__bF$buf4),
    .C(_154_),
    .Y(_28_[29])
);

NOR2X1 _701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[30]),
    .B(_110_),
    .Y(_155_)
);

OAI21X1 _702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114__bF$buf3),
    .B(CSR_Wdata[30]),
    .C(_112__bF$buf5),
    .Y(_156_)
);

NOR2X1 _703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_155_),
    .B(_156_),
    .Y(_28_[30])
);

NAND3X1 _704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mstatus[0]),
    .B(mie),
    .C(mip),
    .Y(_157_)
);

INVX1 _705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_157_),
    .Y(_485_)
);

NAND2X1 _706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mcause[31]),
    .B(_112__bF$buf4),
    .Y(_158_)
);

OAI22X1 _707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112__bF$buf3),
    .B(_157_),
    .C(_110_),
    .D(_158_),
    .Y(_28_[31])
);

INVX1 _708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen),
    .Y(_159_)
);

NOR2X1 _709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7_),
    .B(_60_),
    .Y(_160_)
);

NAND2X1 _710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_160_),
    .B(_17_),
    .Y(_161_)
);

NOR2X1 _711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_159_),
    .B(_161_),
    .Y(_162_)
);

INVX1 _712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[3]),
    .Y(_163_)
);

NAND2X1 _713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_163_),
    .B(_162_),
    .Y(_164_)
);

OAI21X1 _714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mstatus[0]),
    .B(_162_),
    .C(_164_),
    .Y(_165_)
);

OAI21X1 _715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_108__bF$buf2),
    .B(mstatus[1]),
    .C(_112__bF$buf2),
    .Y(_166_)
);

AOI21X1 _716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_108__bF$buf1),
    .B(_165_),
    .C(_166_),
    .Y(_33_[0])
);

MUX2X1 _717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[7]),
    .B(mstatus[1]),
    .S(_162_),
    .Y(_167_)
);

NOR2X1 _718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Ret_bF$buf4),
    .B(CSR_Wen_traps_bF$buf5),
    .Y(_168_)
);

AOI22X1 _719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_34_),
    .B(CSR_Wen_traps_bF$buf4),
    .C(_167_),
    .D(_168_),
    .Y(_33_[1])
);

NOR2X1 _720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf3),
    .B(_109_),
    .Y(_169_)
);

NAND2X1 _721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_169_),
    .B(_24__bF$buf3),
    .Y(_170_)
);

NOR2X1 _722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[0]),
    .B(_170__bF$buf6),
    .Y(_171_)
);

AOI21X1 _723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_),
    .B(_170__bF$buf5),
    .C(_171_),
    .Y(_07_[0])
);

NOR2X1 _724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[1]),
    .B(_170__bF$buf4),
    .Y(_172_)
);

AOI21X1 _725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_26_),
    .B(_170__bF$buf3),
    .C(_172_),
    .Y(_07_[1])
);

INVX1 _726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[2]),
    .Y(_173_)
);

NOR2X1 _727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[2]),
    .B(_170__bF$buf2),
    .Y(_174_)
);

AOI21X1 _728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_173_),
    .B(_170__bF$buf1),
    .C(_174_),
    .Y(_07_[2])
);

INVX2 _729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[3]),
    .Y(_175_)
);

MUX2X1 _730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_175_),
    .B(_163_),
    .S(_170__bF$buf0),
    .Y(_07_[3])
);

INVX2 _731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[4]),
    .Y(_176_)
);

NOR2X1 _732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[4]),
    .B(_170__bF$buf6),
    .Y(_177_)
);

AOI21X1 _733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_176_),
    .B(_170__bF$buf5),
    .C(_177_),
    .Y(_07_[4])
);

INVX2 _734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[5]),
    .Y(_178_)
);

NOR2X1 _735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[5]),
    .B(_170__bF$buf4),
    .Y(_179_)
);

AOI21X1 _736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_178_),
    .B(_170__bF$buf3),
    .C(_179_),
    .Y(_07_[5])
);

INVX2 _737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[6]),
    .Y(_180_)
);

NOR2X1 _738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[6]),
    .B(_170__bF$buf2),
    .Y(_181_)
);

AOI21X1 _739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_180_),
    .B(_170__bF$buf1),
    .C(_181_),
    .Y(_07_[6])
);

INVX1 _740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[7]),
    .Y(_182_)
);

NOR2X1 _741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[7]),
    .B(_170__bF$buf0),
    .Y(_183_)
);

AOI21X1 _742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_182_),
    .B(_170__bF$buf6),
    .C(_183_),
    .Y(_07_[7])
);

INVX1 _743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[8]),
    .Y(_184_)
);

NOR2X1 _744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[8]),
    .B(_170__bF$buf5),
    .Y(_185_)
);

AOI21X1 _745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_184_),
    .B(_170__bF$buf4),
    .C(_185_),
    .Y(_07_[8])
);

INVX1 _746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[9]),
    .Y(_186_)
);

NOR2X1 _747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[9]),
    .B(_170__bF$buf3),
    .Y(_187_)
);

AOI21X1 _748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_186_),
    .B(_170__bF$buf2),
    .C(_187_),
    .Y(_07_[9])
);

INVX2 _749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[10]),
    .Y(_188_)
);

NOR2X1 _750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[10]),
    .B(_170__bF$buf1),
    .Y(_189_)
);

AOI21X1 _751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_188_),
    .B(_170__bF$buf0),
    .C(_189_),
    .Y(_07_[10])
);

INVX1 _752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[11]),
    .Y(_190_)
);

INVX1 _753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[11]),
    .Y(_191_)
);

MUX2X1 _754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(_191_),
    .S(_170__bF$buf6),
    .Y(_07_[11])
);

INVX2 _755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[12]),
    .Y(_192_)
);

NOR2X1 _756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[12]),
    .B(_170__bF$buf5),
    .Y(_193_)
);

AOI21X1 _757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_192_),
    .B(_170__bF$buf4),
    .C(_193_),
    .Y(_07_[12])
);

INVX1 _758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[13]),
    .Y(_194_)
);

NOR2X1 _759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[13]),
    .B(_170__bF$buf3),
    .Y(_195_)
);

AOI21X1 _760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_194_),
    .B(_170__bF$buf2),
    .C(_195_),
    .Y(_07_[13])
);

INVX2 _761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[14]),
    .Y(_196_)
);

NOR2X1 _762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[14]),
    .B(_170__bF$buf1),
    .Y(_197_)
);

AOI21X1 _763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_196_),
    .B(_170__bF$buf0),
    .C(_197_),
    .Y(_07_[14])
);

INVX1 _764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[15]),
    .Y(_198_)
);

NOR2X1 _765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[15]),
    .B(_170__bF$buf6),
    .Y(_199_)
);

AOI21X1 _766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_198_),
    .B(_170__bF$buf5),
    .C(_199_),
    .Y(_07_[15])
);

INVX1 _767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[16]),
    .Y(_200_)
);

NOR2X1 _768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[16]),
    .B(_170__bF$buf4),
    .Y(_201_)
);

AOI21X1 _769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_200_),
    .B(_170__bF$buf3),
    .C(_201_),
    .Y(_07_[16])
);

INVX1 _770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[17]),
    .Y(_202_)
);

NOR2X1 _771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[17]),
    .B(_170__bF$buf2),
    .Y(_203_)
);

AOI21X1 _772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_202_),
    .B(_170__bF$buf1),
    .C(_203_),
    .Y(_07_[17])
);

INVX1 _773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[18]),
    .Y(_204_)
);

NOR2X1 _774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[18]),
    .B(_170__bF$buf0),
    .Y(_205_)
);

AOI21X1 _775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_204_),
    .B(_170__bF$buf6),
    .C(_205_),
    .Y(_07_[18])
);

INVX1 _776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[19]),
    .Y(_206_)
);

NOR2X1 _777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[19]),
    .B(_170__bF$buf5),
    .Y(_207_)
);

AOI21X1 _778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_206_),
    .B(_170__bF$buf4),
    .C(_207_),
    .Y(_07_[19])
);

INVX2 _779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[20]),
    .Y(_208_)
);

NOR2X1 _780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[20]),
    .B(_170__bF$buf3),
    .Y(_209_)
);

AOI21X1 _781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_208_),
    .B(_170__bF$buf2),
    .C(_209_),
    .Y(_07_[20])
);

INVX1 _782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[21]),
    .Y(_210_)
);

NOR2X1 _783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[21]),
    .B(_170__bF$buf1),
    .Y(_211_)
);

AOI21X1 _784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_210_),
    .B(_170__bF$buf0),
    .C(_211_),
    .Y(_07_[21])
);

INVX1 _785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[22]),
    .Y(_212_)
);

NOR2X1 _786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[22]),
    .B(_170__bF$buf6),
    .Y(_213_)
);

AOI21X1 _787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_212_),
    .B(_170__bF$buf5),
    .C(_213_),
    .Y(_07_[22])
);

INVX1 _788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[23]),
    .Y(_214_)
);

NOR2X1 _789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[23]),
    .B(_170__bF$buf4),
    .Y(_215_)
);

AOI21X1 _790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_214_),
    .B(_170__bF$buf3),
    .C(_215_),
    .Y(_07_[23])
);

INVX1 _791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[24]),
    .Y(_216_)
);

NOR2X1 _792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[24]),
    .B(_170__bF$buf2),
    .Y(_217_)
);

AOI21X1 _793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_216_),
    .B(_170__bF$buf1),
    .C(_217_),
    .Y(_07_[24])
);

INVX1 _794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[25]),
    .Y(_218_)
);

NOR2X1 _795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[25]),
    .B(_170__bF$buf0),
    .Y(_219_)
);

AOI21X1 _796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_218_),
    .B(_170__bF$buf6),
    .C(_219_),
    .Y(_07_[25])
);

INVX1 _797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[26]),
    .Y(_220_)
);

NOR2X1 _798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[26]),
    .B(_170__bF$buf5),
    .Y(_221_)
);

AOI21X1 _799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_220_),
    .B(_170__bF$buf4),
    .C(_221_),
    .Y(_07_[26])
);

INVX1 _800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[27]),
    .Y(_222_)
);

NOR2X1 _801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[27]),
    .B(_170__bF$buf3),
    .Y(_223_)
);

AOI21X1 _802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_222_),
    .B(_170__bF$buf2),
    .C(_223_),
    .Y(_07_[27])
);

INVX1 _803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[28]),
    .Y(_224_)
);

NOR2X1 _804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[28]),
    .B(_170__bF$buf1),
    .Y(_225_)
);

AOI21X1 _805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_224_),
    .B(_170__bF$buf0),
    .C(_225_),
    .Y(_07_[28])
);

INVX1 _806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[29]),
    .Y(_226_)
);

NOR2X1 _807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[29]),
    .B(_170__bF$buf6),
    .Y(_227_)
);

AOI21X1 _808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_226_),
    .B(_170__bF$buf5),
    .C(_227_),
    .Y(_07_[29])
);

INVX1 _809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[30]),
    .Y(_228_)
);

NOR2X1 _810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[30]),
    .B(_170__bF$buf4),
    .Y(_229_)
);

AOI21X1 _811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_228_),
    .B(_170__bF$buf3),
    .C(_229_),
    .Y(_07_[30])
);

INVX1 _812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[31]),
    .Y(_230_)
);

NOR2X1 _813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wdata[31]),
    .B(_170__bF$buf2),
    .Y(_231_)
);

AOI21X1 _814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_230_),
    .B(_170__bF$buf1),
    .C(_231_),
    .Y(_07_[31])
);

NAND2X1 _815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_169_),
    .B(_64_),
    .Y(_232_)
);

NAND2X1 _816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mie),
    .B(_232_),
    .Y(_233_)
);

OAI21X1 _817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_191_),
    .B(_232_),
    .C(_233_),
    .Y(_14_)
);

NAND2X1 _818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf2),
    .B(CSR_mepc[2]),
    .Y(_234_)
);

AND2X2 _819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_31__bF$buf4),
    .B(_113_),
    .Y(_235_)
);

NOR2X1 _820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[0]),
    .B(_235__bF$buf4),
    .Y(_236_)
);

NAND2X1 _821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_113_),
    .B(_31__bF$buf3),
    .Y(_237_)
);

OAI21X1 _822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf4),
    .B(CSR_Wdata[2]),
    .C(_112__bF$buf1),
    .Y(_238_)
);

OAI21X1 _823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_236_),
    .B(_238_),
    .C(_234_),
    .Y(_21_[0])
);

NAND2X1 _824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf1),
    .B(CSR_mepc[3]),
    .Y(_239_)
);

NOR2X1 _825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[1]),
    .B(_235__bF$buf3),
    .Y(_240_)
);

OAI21X1 _826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf3),
    .B(CSR_Wdata[3]),
    .C(_112__bF$buf0),
    .Y(_241_)
);

OAI21X1 _827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_240_),
    .B(_241_),
    .C(_239_),
    .Y(_21_[1])
);

NAND2X1 _828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf0),
    .B(CSR_mepc[4]),
    .Y(_242_)
);

NOR2X1 _829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[2]),
    .B(_235__bF$buf2),
    .Y(_243_)
);

OAI21X1 _830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf2),
    .B(CSR_Wdata[4]),
    .C(_112__bF$buf6),
    .Y(_244_)
);

OAI21X1 _831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_243_),
    .B(_244_),
    .C(_242_),
    .Y(_21_[2])
);

NAND2X1 _832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf5),
    .B(CSR_mepc[5]),
    .Y(_245_)
);

NOR2X1 _833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[3]),
    .B(_235__bF$buf1),
    .Y(_246_)
);

OAI21X1 _834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf1),
    .B(CSR_Wdata[5]),
    .C(_112__bF$buf5),
    .Y(_247_)
);

OAI21X1 _835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_246_),
    .B(_247_),
    .C(_245_),
    .Y(_21_[3])
);

NAND2X1 _836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf4),
    .B(CSR_mepc[6]),
    .Y(_248_)
);

NOR2X1 _837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[4]),
    .B(_235__bF$buf0),
    .Y(_249_)
);

OAI21X1 _838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf0),
    .B(CSR_Wdata[6]),
    .C(_112__bF$buf4),
    .Y(_250_)
);

OAI21X1 _839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_249_),
    .B(_250_),
    .C(_248_),
    .Y(_21_[4])
);

NAND2X1 _840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf3),
    .B(CSR_mepc[7]),
    .Y(_251_)
);

NOR2X1 _841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[5]),
    .B(_235__bF$buf4),
    .Y(_252_)
);

OAI21X1 _842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf4),
    .B(CSR_Wdata[7]),
    .C(_112__bF$buf3),
    .Y(_253_)
);

OAI21X1 _843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_252_),
    .B(_253_),
    .C(_251_),
    .Y(_21_[5])
);

NAND2X1 _844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf2),
    .B(CSR_mepc[8]),
    .Y(_254_)
);

NOR2X1 _845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[6]),
    .B(_235__bF$buf3),
    .Y(_255_)
);

OAI21X1 _846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf3),
    .B(CSR_Wdata[8]),
    .C(_112__bF$buf2),
    .Y(_256_)
);

OAI21X1 _847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(_256_),
    .C(_254_),
    .Y(_21_[6])
);

NAND2X1 _848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf1),
    .B(CSR_mepc[9]),
    .Y(_257_)
);

NOR2X1 _849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[7]),
    .B(_235__bF$buf2),
    .Y(_258_)
);

OAI21X1 _850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf2),
    .B(CSR_Wdata[9]),
    .C(_112__bF$buf1),
    .Y(_259_)
);

OAI21X1 _851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_258_),
    .B(_259_),
    .C(_257_),
    .Y(_21_[7])
);

NAND2X1 _852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf0),
    .B(CSR_mepc[10]),
    .Y(_260_)
);

NOR2X1 _853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[8]),
    .B(_235__bF$buf1),
    .Y(_261_)
);

OAI21X1 _854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf1),
    .B(CSR_Wdata[10]),
    .C(_112__bF$buf0),
    .Y(_262_)
);

OAI21X1 _855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_261_),
    .B(_262_),
    .C(_260_),
    .Y(_21_[8])
);

NAND2X1 _856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf5),
    .B(CSR_mepc[11]),
    .Y(_263_)
);

NOR2X1 _857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[9]),
    .B(_235__bF$buf0),
    .Y(_264_)
);

OAI21X1 _858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf0),
    .B(CSR_Wdata[11]),
    .C(_112__bF$buf6),
    .Y(_265_)
);

OAI21X1 _859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_264_),
    .B(_265_),
    .C(_263_),
    .Y(_21_[9])
);

NAND2X1 _860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf4),
    .B(CSR_mepc[12]),
    .Y(_266_)
);

NOR2X1 _861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[10]),
    .B(_235__bF$buf4),
    .Y(_267_)
);

OAI21X1 _862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf4),
    .B(CSR_Wdata[12]),
    .C(_112__bF$buf5),
    .Y(_268_)
);

OAI21X1 _863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_267_),
    .B(_268_),
    .C(_266_),
    .Y(_21_[10])
);

NAND2X1 _864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf3),
    .B(CSR_mepc[13]),
    .Y(_269_)
);

NOR2X1 _865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[11]),
    .B(_235__bF$buf3),
    .Y(_270_)
);

OAI21X1 _866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf3),
    .B(CSR_Wdata[13]),
    .C(_112__bF$buf4),
    .Y(_271_)
);

OAI21X1 _867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_270_),
    .B(_271_),
    .C(_269_),
    .Y(_21_[11])
);

NAND2X1 _868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf2),
    .B(CSR_mepc[14]),
    .Y(_272_)
);

NOR2X1 _869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[12]),
    .B(_235__bF$buf2),
    .Y(_273_)
);

OAI21X1 _870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf2),
    .B(CSR_Wdata[14]),
    .C(_112__bF$buf3),
    .Y(_274_)
);

OAI21X1 _871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_273_),
    .B(_274_),
    .C(_272_),
    .Y(_21_[12])
);

NAND2X1 _872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf1),
    .B(CSR_mepc[15]),
    .Y(_275_)
);

NOR2X1 _873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[13]),
    .B(_235__bF$buf1),
    .Y(_276_)
);

OAI21X1 _874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf1),
    .B(CSR_Wdata[15]),
    .C(_112__bF$buf2),
    .Y(_277_)
);

OAI21X1 _875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_276_),
    .B(_277_),
    .C(_275_),
    .Y(_21_[13])
);

NAND2X1 _876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf0),
    .B(CSR_mepc[16]),
    .Y(_278_)
);

NOR2X1 _877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[14]),
    .B(_235__bF$buf0),
    .Y(_279_)
);

OAI21X1 _878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf0),
    .B(CSR_Wdata[16]),
    .C(_112__bF$buf1),
    .Y(_280_)
);

OAI21X1 _879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_279_),
    .B(_280_),
    .C(_278_),
    .Y(_21_[14])
);

NAND2X1 _880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf5),
    .B(CSR_mepc[17]),
    .Y(_281_)
);

NOR2X1 _881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[15]),
    .B(_235__bF$buf4),
    .Y(_282_)
);

OAI21X1 _882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf4),
    .B(CSR_Wdata[17]),
    .C(_112__bF$buf0),
    .Y(_283_)
);

OAI21X1 _883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_282_),
    .B(_283_),
    .C(_281_),
    .Y(_21_[15])
);

NAND2X1 _884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf4),
    .B(CSR_mepc[18]),
    .Y(_284_)
);

NOR2X1 _885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[16]),
    .B(_235__bF$buf3),
    .Y(_285_)
);

OAI21X1 _886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf3),
    .B(CSR_Wdata[18]),
    .C(_112__bF$buf6),
    .Y(_286_)
);

OAI21X1 _887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_285_),
    .B(_286_),
    .C(_284_),
    .Y(_21_[16])
);

NAND2X1 _888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf3),
    .B(CSR_mepc[19]),
    .Y(_287_)
);

NOR2X1 _889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[17]),
    .B(_235__bF$buf2),
    .Y(_288_)
);

OAI21X1 _890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf2),
    .B(CSR_Wdata[19]),
    .C(_112__bF$buf5),
    .Y(_289_)
);

OAI21X1 _891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_288_),
    .B(_289_),
    .C(_287_),
    .Y(_21_[17])
);

NAND2X1 _892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf2),
    .B(CSR_mepc[20]),
    .Y(_290_)
);

NOR2X1 _893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[18]),
    .B(_235__bF$buf1),
    .Y(_291_)
);

OAI21X1 _894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf1),
    .B(CSR_Wdata[20]),
    .C(_112__bF$buf4),
    .Y(_292_)
);

OAI21X1 _895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_291_),
    .B(_292_),
    .C(_290_),
    .Y(_21_[18])
);

NAND2X1 _896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf1),
    .B(CSR_mepc[21]),
    .Y(_293_)
);

NOR2X1 _897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[19]),
    .B(_235__bF$buf0),
    .Y(_294_)
);

OAI21X1 _898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf0),
    .B(CSR_Wdata[21]),
    .C(_112__bF$buf3),
    .Y(_295_)
);

OAI21X1 _899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_294_),
    .B(_295_),
    .C(_293_),
    .Y(_21_[19])
);

NAND2X1 _900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf0),
    .B(CSR_mepc[22]),
    .Y(_296_)
);

NOR2X1 _901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[20]),
    .B(_235__bF$buf4),
    .Y(_297_)
);

OAI21X1 _902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf4),
    .B(CSR_Wdata[22]),
    .C(_112__bF$buf2),
    .Y(_298_)
);

OAI21X1 _903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .B(_298_),
    .C(_296_),
    .Y(_21_[20])
);

NAND2X1 _904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf5),
    .B(CSR_mepc[23]),
    .Y(_299_)
);

NOR2X1 _905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[21]),
    .B(_235__bF$buf3),
    .Y(_300_)
);

OAI21X1 _906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf3),
    .B(CSR_Wdata[23]),
    .C(_112__bF$buf1),
    .Y(_301_)
);

OAI21X1 _907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_300_),
    .B(_301_),
    .C(_299_),
    .Y(_21_[21])
);

NAND2X1 _908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf4),
    .B(CSR_mepc[24]),
    .Y(_302_)
);

NOR2X1 _909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[22]),
    .B(_235__bF$buf2),
    .Y(_303_)
);

OAI21X1 _910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf2),
    .B(CSR_Wdata[24]),
    .C(_112__bF$buf0),
    .Y(_304_)
);

OAI21X1 _911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_303_),
    .B(_304_),
    .C(_302_),
    .Y(_21_[22])
);

NAND2X1 _912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf3),
    .B(CSR_mepc[25]),
    .Y(_305_)
);

NOR2X1 _913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[23]),
    .B(_235__bF$buf1),
    .Y(_306_)
);

OAI21X1 _914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf1),
    .B(CSR_Wdata[25]),
    .C(_112__bF$buf6),
    .Y(_307_)
);

OAI21X1 _915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_306_),
    .B(_307_),
    .C(_305_),
    .Y(_21_[23])
);

NAND2X1 _916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf2),
    .B(CSR_mepc[26]),
    .Y(_308_)
);

NOR2X1 _917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[24]),
    .B(_235__bF$buf0),
    .Y(_309_)
);

OAI21X1 _918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf0),
    .B(CSR_Wdata[26]),
    .C(_112__bF$buf5),
    .Y(_310_)
);

OAI21X1 _919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_309_),
    .B(_310_),
    .C(_308_),
    .Y(_21_[24])
);

NAND2X1 _920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf1),
    .B(CSR_mepc[27]),
    .Y(_311_)
);

NOR2X1 _921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[25]),
    .B(_235__bF$buf4),
    .Y(_312_)
);

OAI21X1 _922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf4),
    .B(CSR_Wdata[27]),
    .C(_112__bF$buf4),
    .Y(_313_)
);

OAI21X1 _923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_312_),
    .B(_313_),
    .C(_311_),
    .Y(_21_[25])
);

NAND2X1 _924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf0),
    .B(CSR_mepc[28]),
    .Y(_314_)
);

NOR2X1 _925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[26]),
    .B(_235__bF$buf3),
    .Y(_315_)
);

OAI21X1 _926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf3),
    .B(CSR_Wdata[28]),
    .C(_112__bF$buf3),
    .Y(_316_)
);

OAI21X1 _927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_315_),
    .B(_316_),
    .C(_314_),
    .Y(_21_[26])
);

NAND2X1 _928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf5),
    .B(CSR_mepc[29]),
    .Y(_317_)
);

NOR2X1 _929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[27]),
    .B(_235__bF$buf2),
    .Y(_318_)
);

OAI21X1 _930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf2),
    .B(CSR_Wdata[29]),
    .C(_112__bF$buf2),
    .Y(_319_)
);

OAI21X1 _931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_318_),
    .B(_319_),
    .C(_317_),
    .Y(_21_[27])
);

NAND2X1 _932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf4),
    .B(CSR_mepc[30]),
    .Y(_320_)
);

NOR2X1 _933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[28]),
    .B(_235__bF$buf1),
    .Y(_321_)
);

OAI21X1 _934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf1),
    .B(CSR_Wdata[30]),
    .C(_112__bF$buf1),
    .Y(_322_)
);

OAI21X1 _935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_321_),
    .B(_322_),
    .C(_320_),
    .Y(_21_[28])
);

NAND2X1 _936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(CSR_Wen_traps_bF$buf3),
    .B(CSR_mepc[31]),
    .Y(_323_)
);

NOR2X1 _937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[29]),
    .B(_235__bF$buf0),
    .Y(_324_)
);

OAI21X1 _938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237__bF$buf0),
    .B(CSR_Wdata[31]),
    .C(_112__bF$buf0),
    .Y(_325_)
);

OAI21X1 _939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_324_),
    .B(_325_),
    .C(_323_),
    .Y(_21_[29])
);

NOR2X1 _940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_),
    .B(_157_),
    .Y(_326_)
);

NAND2X1 _941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_173_),
    .B(_326_),
    .Y(_327_)
);

INVX2 _942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_326_),
    .Y(_328_)
);

AOI21X1 _943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[2]),
    .B(_328_),
    .C(CSR_Ret_bF$buf3),
    .Y(_329_)
);

NOR2X1 _944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[0]),
    .B(_108__bF$buf0),
    .Y(_330_)
);

AOI21X1 _945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_327_),
    .B(_329_),
    .C(_330_),
    .Y(_486_[2])
);

XNOR2X1 _946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_327_),
    .B(_175_),
    .Y(_331_)
);

NAND2X1 _947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[1]),
    .B(CSR_Ret_bF$buf2),
    .Y(_332_)
);

OAI21X1 _948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_331_),
    .B(CSR_Ret_bF$buf1),
    .C(_332_),
    .Y(_486_[3])
);

NOR2X1 _949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[2]),
    .B(mvect[3]),
    .Y(_333_)
);

OAI21X1 _950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_328_),
    .B(_333_),
    .C(_176_),
    .Y(_334_)
);

OAI21X1 _951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[2]),
    .B(mvect[3]),
    .C(mvect[4]),
    .Y(_335_)
);

OAI21X1 _952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_328_),
    .B(_335_),
    .C(_334_),
    .Y(_336_)
);

NAND2X1 _953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[2]),
    .B(CSR_Ret_bF$buf0),
    .Y(_337_)
);

OAI21X1 _954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_336_),
    .B(CSR_Ret_bF$buf5),
    .C(_337_),
    .Y(_486_[4])
);

OAI21X1 _955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_176_),
    .B(_333_),
    .C(_326_),
    .Y(_338_)
);

XNOR2X1 _956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_338_),
    .B(_178_),
    .Y(_339_)
);

NAND2X1 _957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[3]),
    .B(CSR_Ret_bF$buf4),
    .Y(_340_)
);

OAI21X1 _958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_339_),
    .B(CSR_Ret_bF$buf3),
    .C(_340_),
    .Y(_486_[5])
);

OAI21X1 _959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_333_),
    .B(_176_),
    .C(_178_),
    .Y(_341_)
);

AOI21X1 _960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_326_),
    .B(_341_),
    .C(mvect[6]),
    .Y(_342_)
);

NAND2X1 _961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_326_),
    .B(_341_),
    .Y(_343_)
);

OAI21X1 _962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_343_),
    .B(_180_),
    .C(_108__bF$buf4),
    .Y(_344_)
);

NAND2X1 _963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[4]),
    .B(CSR_Ret_bF$buf2),
    .Y(_345_)
);

OAI21X1 _964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_344_),
    .B(_342_),
    .C(_345_),
    .Y(_486_[6])
);

OAI21X1 _965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_343_),
    .B(_180_),
    .C(_182_),
    .Y(_346_)
);

NAND2X1 _966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[6]),
    .B(mvect[7]),
    .Y(_347_)
);

OAI21X1 _967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_343_),
    .B(_347_),
    .C(_346_),
    .Y(_348_)
);

NAND2X1 _968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[5]),
    .B(CSR_Ret_bF$buf1),
    .Y(_349_)
);

OAI21X1 _969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_348_),
    .B(CSR_Ret_bF$buf0),
    .C(_349_),
    .Y(_486_[7])
);

AOI21X1 _970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_178_),
    .B(_335_),
    .C(_347_),
    .Y(_350_)
);

AND2X2 _971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_350_),
    .B(_326_),
    .Y(_351_)
);

NAND2X1 _972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[8]),
    .B(_351_),
    .Y(_352_)
);

INVX1 _973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_352_),
    .Y(_353_)
);

OAI21X1 _974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_351_),
    .B(mvect[8]),
    .C(_108__bF$buf3),
    .Y(_354_)
);

NAND2X1 _975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[6]),
    .B(CSR_Ret_bF$buf5),
    .Y(_355_)
);

OAI21X1 _976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_353_),
    .B(_354_),
    .C(_355_),
    .Y(_486_[8])
);

NAND2X1 _977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_326_),
    .B(_350_),
    .Y(_356_)
);

OAI21X1 _978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_356_),
    .B(_184_),
    .C(_186_),
    .Y(_357_)
);

NAND2X1 _979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[8]),
    .B(mvect[9]),
    .Y(_358_)
);

OAI21X1 _980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_356_),
    .B(_358_),
    .C(_357_),
    .Y(_359_)
);

NAND2X1 _981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[7]),
    .B(CSR_Ret_bF$buf4),
    .Y(_360_)
);

OAI21X1 _982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_359_),
    .B(CSR_Ret_bF$buf3),
    .C(_360_),
    .Y(_486_[9])
);

INVX1 _983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_358_),
    .Y(_361_)
);

NAND2X1 _984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_361_),
    .B(_351_),
    .Y(_362_)
);

XNOR2X1 _985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_362_),
    .B(_188_),
    .Y(_363_)
);

NAND2X1 _986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[8]),
    .B(CSR_Ret_bF$buf2),
    .Y(_364_)
);

OAI21X1 _987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_363_),
    .B(CSR_Ret_bF$buf1),
    .C(_364_),
    .Y(_486_[10])
);

NAND2X1 _988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[10]),
    .B(_361_),
    .Y(_365_)
);

OAI21X1 _989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_356_),
    .B(_365_),
    .C(_190_),
    .Y(_366_)
);

NAND2X1 _990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mvect[10]),
    .B(mvect[11]),
    .Y(_367_)
);

OR2X2 _991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_358_),
    .B(_367_),
    .Y(_368_)
);

OAI21X1 _992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_356_),
    .B(_368_),
    .C(_366_),
    .Y(_369_)
);

NAND2X1 _993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[9]),
    .B(CSR_Ret_bF$buf0),
    .Y(_370_)
);

OAI21X1 _994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_369_),
    .B(CSR_Ret_bF$buf5),
    .C(_370_),
    .Y(_486_[11])
);

NOR2X1 _995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_358_),
    .B(_367_),
    .Y(_371_)
);

NAND3X1 _996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_326_),
    .B(_371_),
    .C(_350_),
    .Y(_372_)
);

XNOR2X1 _997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_372_),
    .B(_192_),
    .Y(_373_)
);

NAND2X1 _998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(mepc[10]),
    .B(CSR_Ret_bF$buf4),
    .Y(_374_)
);

OAI21X1 _999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_373_),
    .B(CSR_Ret_bF$buf3),
    .C(_374_),
    .Y(_486_[12])
);

endmodule
